`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
V9fjqhLmJ82PDFazD0ucMWcFBY9BITDqvsp3Ku7A0AVrAxczp/IiUYOLLNgAtH/tpyNRkdzuwoAP
EJv5zrsbJw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
AjkdpdDjqsDrpBtI8KrRd4EBKsFJPg56xmPmrzKbEagUb81sKZHNAiT6rzNgZkJJM0cgNTD8y52h
z4sSsZYmZLpRBhZYxchS0ZC8WuZiCQYMi8lZz04lgDU/xJkXvNWOIuJfcuN2JV4I71n6snByvfbc
rH1j6MkywWjxa1DnBNM=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2rpPC0jQWYFFbxUR7SjYwZCotNh7v8TZDXBF8QAbPwFIKMlpf1mt6QarI+woa5SeI4MaRzYl0/V1
QxWEN9GTn2YX1lwIpSZO/dgdFgfB6+CfYD2936vFi9B537eUUf4IoCOvCVLqlH02QUncN0JQq4MI
ilm/UHplvZlJfB/NWzY=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IK1IVhBG0OBjzZJ+lbZ9m6ad61iN/w7PK02g5mI+n/vZFub6hGZHtA4TfZDy8/Azd/20BJHFkQ2y
vLaMSqDYdKiviwYRuLBlsFIjA1JPBe7I5qNwzSWowBWY+Tz6p3GF1dhNI6Eu4udDS6R9SjvjDfRX
KfPfZykRmxhmPakpFfHP17r8QKsBQmc7IBzjdfwJCqifh3Vezh4zVSGZ2npz33m/MqJqCNMcZD9N
KMfFAhEG6nenq99DwFpEPHiKuZwF9F2thTm1MZx0beFzMQ7vGjGeI6GlskLsznrY83gjzt/aYHsR
rb6T3P3OcuTGXIb+mvUzPgMV2xLFwnwAqMnGYA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HDX5a3xzdZbgrKLFF0sB8hU8xh5y5RVU1qs90ujzF7Lpw2gh7FqRNaYMfnauQQVWZbIME9ImheHq
DrEGGcM/12GCLJtzt4MSE2AldJSQoGHikzYITF92vmW4SXwZgv8LjTjh0iPTmJccFrtIGzs9AmFu
kzu7h3vEeHESMY5Rztw8EHOX6A0/d7tk6HnBW5mB8i0SSm98PKrqJg9exPrwm7Zbbtr/BYVArS0m
ECyg121HBfLon/KTNeg21klZi/cEiihwYs/J48o5RxLYO5/R8SVTu2hYmJbWekMe8IAqJsJZ2T0q
QTrO4NUmLB4Yzn5aRro69gKXXmxekJvzjmS1Aw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
O18o+ZXV9y8FX22WmYGVCqemJA1CaC4IS7h7WpPatSfHkpOEpdGxXoyXcYl7vvrUnBD2G3xMVtBY
Ho6YzCoQxNWpSpMg71NYr7CG7copGhp78kWQaeA6Lgtf72q/l6KWxdm3/qhctzKn78S9+3PBCVs5
fPsp7Nt1UQKtt5jCpJtSf29Ey1KE4ySkoPWRV4H+ZDu0Cy0V8EJd91mIj6Y6bVON7c1hMH3vi6tn
E+ZSPpvXrIxKktpz0MfHda/gNjkWWHRDpCuT57G3x2SW9+ngKSs+iqFqhMdWOpqv8N7iNjxQEIEz
VjVWPUK4owPn3/P6WXnVkZWx0Wo8grGwoyho9w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 779472)
`protect data_block
mIstQombYn4BQocLjDAJHm9fwZN2RSGWGkbueKDwpCCvk4j56Jmp0dlSwRsp1JQoZF1/j9latsrx
8MMn/6Z49wRp/WuQ9xb8sNesz+ezvWFIbk6dl0/BrcuEqUo9iK2fpxzwrzSEy6zG+laKAC5UP8ff
NvosG9Nel5ZmMbxFdcuRual58kzzDPg9wX1IT7ve6ODsc3kKKbMgpshxYjMhYTQlLEdKCZRIuI4k
8cax1PLQANQyB0zeKjuC5TuQpXB8+EghZYknDCxVSSldT5AYCZxu740jJKcJy9pdd2yF5DXqKZFP
S+XSdiiNAwXnNkMZ0uzepkwViKdUbUwYWxRZiLU/i99f80HaKd3YJytgF4aWXLVGi8mLdIfPpuux
WW960oX4kYEZM88tUC9rqCl3KUMiE7flEsG/I7OAepinjFaI0Ihcx92nm8D/KPkQtQ0x1wD+d/mC
6j16j21eSy8869QGQpMJ1ED9XMi61sBHG0WoeVe+MdI3JzC23RtSRe0fySHvfJJw6qfEUxu73wAl
zuVieyUW1c4XtgMnh7SM7CMmTKINLlNxcDKGdk7b0N4cjSQeD1DlAkgsHnjO4D4PWVEpaQNPRvOR
RZ9FWKuP2a9IRYpLhAfEXGnq7vJJxx3zwhfy66C+/56uQot4Sc8cONGbdFqPxWQ4a2Z6vsdghm9b
r8wmP2D5z7o4sBgKGwkIPXWeV1ZT861CRkGI+hfm0kB2we4UvQlwbygz3qPTucyxGg0272WLamNb
6zxN2KrD2YzBmg7FGt5FegMJzr0bC05aUDrdG2eYoE+G8w3bB9iDPGUs6SCBlL9cKjXPrsCb8YFh
3YZSP5/K95X2xKB6Mvc9FBG6WPCeq6NfAM8WomxQmhlbJm/8qyQtJceNBNqxpxOdd8u6OckIJNUI
LU1ONAKYS+Vj5dFylITlM8XR8DX0u12ZTIsO2ziM3jWFnvNRHpad8CCVLA20MuhNipuK+modwUs3
ZHnpUGRiDG95O+OlXef/E+M3rdTDY3GVVN5DutvJcL2AmH0uWEdNnJqD9wIX/uyM95UyZU3Z+MVU
y/mjwEPVNjMRKGz61gAmfcRYQjq2EzpX2oqfgZ58vSeuOtR8CrJ5kUERq276y1YqCI/65a+DUYgz
Ig8XDnN+mAZmnDXnk1zVXdx1EymtwQoZeyjMkldQUObAda1zTRDc1XPP6YGecaflO6UQ85x5XI/1
z6PupNu6TDyCI8qicKgJy4TmX/wf5LNjem8gJANWWmI18psfgUUCdul75LlB3mZU3DhTU6gpARtG
dVUu0s14lAoy2aFa/eCSqS47X/PvRSfzFeLbQtzmB5RtWyw+sVzLfn7HYOfj+eCWGwnAyEnNyRDb
mxvL8vV3jIjQ2fi3KT4LG4vUNpjHYYQoNGPk/T3GHlhrGPR54hKiYVDbs8wLiDn3rrhVRWgJioZY
RHKOaXAcn35zX6UYhxkr3Vu5r0NCO8VSw+yky8POxZwOowThtnADblbVph2ufstmrWHnr2MfbcSr
yi65ptAL5W4BucUCfEjWIuzVWTpD8vvmO0mXcOcoQZ4qC3GXTrihCtYpypgQWcxvHYQUML6anXVb
gUZe2xJGZOO87UjbTrAIuYWFhuSJs/ed+P6nYGiToNWEUmBgjdZ059RLI3+oigYP4pmZvIjrMNzg
QuP8KLOyPyxF/2A8RirckzvWcEZffHlLLzQxVPPOV29RKeRkgjNh1G+wxDY/ZknroB2tqNQYu80N
gahD5t1XJUklRTYm5ZTvpwaawjGhGi5M9HdA9uOdUdY0C8uAIt++wR5amLz7Yf0BYO+eaA8a1IhY
Rr1VBMwbPtgldso3zH8o7N+cz9hjXjUs9E9y+rwlF9Z4ABp4kyWjO+opB7qtEZj4aKWs71nOF2EO
uGjPUFKorLhf7/+la1KLBtRaN8AxdBgpnBopdzYttDTqO+G1IuUl3dqmpK2jRszih91UOwY9ejhm
Fle9jmNNKSmWqnN2jqOquuObbnIBxLREikmWoHKkZeBZC2GM+y5pABfdXaYonIBd8Azyushemivr
qa0ogUkK7MnOcbjnjLa9exiVT1zX0B0OlzMrf0zyxtjtDjEaLF9SOgTP74ldg54Mul/pyG6GiQFj
t1cDqvcsFz6JEPokJ4/3+Yu8/atB8bY1wZG1Dfpir0PX11mG0+LIgyMZwDFEN3HTOlWNRpbJUmx+
ngEdbwbq4ZqTUKAXRr5q8WiPyqTOtWvJ/2SfKzTehQTIs2wNddT7nefFyBMEnPDl8kXULrVt57Xn
jMpbVLplN1NOwC22mpk6DAznIvD6Q3FF/3UH++7KI0NVY93s85vCIn2/ZvaOXWRbrRvk96Z9f4fa
Ulo2VhmJbjUn2EX4LzknEHvFAxL30BZ3u5MUw/BrkNsQ2+5QwvWbiAPC33/J3irFjkYyNndfB4M5
qnmMUw/TotfcqoByW4iffJEzs/+1WU3RxqbRH7Z0BA4vipONCwO7wUVcjtXKWqSJYWlBmcjuoTuM
ifcd5SL4czbB+51Z5gPMqGD5cZT58Tjyb0AyUdbAnNsM7otxN7s1wHApQAIntTwo9cRLtapZDBVw
IFI3LjZqX7y7UdJd/fyPBHYGl5wgITJOEnWTl0UMJzI0IiPg62dZIaRToik/12uofKwbtIRrpC6A
8fw5sYs4DKCSUo/4c5y1WTH9hBJdjOIiPkUexY7POpmLu/WZtnVrcw3e4u8fDkuSIuuJkyylK2M/
y2Ek4y0PBGgwqkJASPz1mLlbQJnFnpU/Jukz4leQZUsO+LtJE0QqkbdJJabZt+1UZ+r6dDi4IPh3
17gZhz8hd1q6YeN/yfLbKSwHIJhxCrAqT6UdIAN+qZQ2yfiv6JeApVRN+tJdT008ElU6WY9LwknO
oyHNPN/B/TViG15pESbMYxzoGuLtrd5LWF+T1UuD6Ev7pz7aPbzP2um/Ffkh1GZiiEEkDKD5Kt92
VR4xOIYRuWrcp18WRMto1RXdIRRBzHmiQy1lxkyIHFoA1YYS/pvxylGtIrjEEdJx6X2BaZFfgsZT
PvhKTZK/1NFXLgpbue0NknIWCmcaIqrWq9MCwKvlkkmlfLo3ryySRKjhYvO+xoPrZ7Aei6ntZtdJ
vUYZQYdeu2nzniAH7OfvmJQsT9lO+ayglLjNGl8oS9Atip8RrH81kS4gByVL9T0/xNuSNDqkKsEg
NyDyTBDvXFX1w0yZNZxPO2Qb2O01xx/cHshvjwrXhevAKNX3gEU43LaNRqJJCVajSgxbW01/aypa
AG/As7meXKam1JbKRDHt5PJegK5UI/xBAtCThoEHQAsvy+9OmtxKaqc4/w1JnCadkJYjxOPXI4v9
cO8RTW8XnFAu7HEz6Plau2BAOyI8nzrTlaOvvyg33uED+ECNxvACwWg8OhNEDTv0TwxA85UkH4uX
OoPHWOZjtuRRcYokiAfQtc9W4GTi2MUu5swjrzB4t8xh8KdwNN/ZqsMmiD3jr4okf3qdYstluTPc
Wpb/t3BjEpqJ2Uy8og5d9cNzaGm8efrkD4ao9ozOY4jOU2nNK+SWqrIqDTnHeIQccMwRmeQTUJoY
nsA2HgxivLZfGSCfYXlsKbH7/M3Nyf+pcn5yLLdBLgCqMmfzryBofAlRl4xtdZrtQuZssMuM69qP
fIPt/nu+AiLqQ52vbF57J4gW99IMDS4sXlAk8Ja1yZzaUnp8HFzpA9rY8LiD+8BPyPqg8+GYHOT0
HCPRdEFPx4zjRB24ugg8Xs8Z9oUxeXGjd7/lNa9rEsG50LSSGHdtQNNsOOASYUOjz5ROiOsihl7L
XUnwgyz8Y9sjUZ7YEs/gleBxrzw5dX0XgM16BH8FIzoS8bhCSLn8EfwesrLl8vySaq5UZmLlkDMn
E3huZKamLinIeyrEodJW8G1eRiyBnN+Dq4T+PclEP8zVaM6HJvtU8Ye2aoLDjMc3agwOh/0Dpv5z
Z5edr8dK0/YI054VW2F/r/rX1GTHu5Q/60JnhjD2DBLQHrnmWF9fZUOYj1t3Wi8TYGhEDo7KbVs9
OcBXgbrv7ur1PTy87qLjY71awnOpqAOsovgfP7vxvghQ3fvbUUgd31nBIzlvA0Uu2RlR7u8Afmvv
n2Ec/SYn2dNCp4WhkK/Ov9lOWgcDi99kn6i/uBjTf10CbQ/vZ8KDjh5/7vXOOkSQEINAZ8FznOTM
PhgDfwQQVtOmF4dbTgtkkuV1mkrRc8MWLMvsjlCn4LMrBvGe2mvb/2fC/5Jl1XJRMy8nUPpJcEZ9
fg0BGJ0Zo920xWddasqnwCznK3FCcw8eT2Ebhb3MP8drQumF3rR4vtOlbQ98WBxrqbZlaE30cqi5
Yv9T/4m1n2tmfs1Vqs9ZcV+fvRQVLqS89X/X6CycBaApfNGgBWFoz1WBbVUPSJSNZVAIW36ALMj4
u3gDrBCxBYuy2OnUmS+SooQZ56j/dTR3eBpruNdzrS+zuYq7CdJKOzdQWOPUTTeMt/Ku67c/pEhm
y9FInI5D9BtEfc1q13lpXsekMRjiZPD01tR9vTa/70KBT6xYOne6u0/k1tgk4qHPQS59BqT6VsQ/
NLUhMQryzuviv6Sbjg2L28EyrE0wGW0MhctpUNgXaGv7szchMbcwtsIkmMFoIPD3TFiFb9lyDL/C
FVik+dGsm5ScSvUAY71MIyDsIELj4aomBUBW5UtAdWV7BKNdfl73/82ey7sCY9EDjR4y3xI5kF0t
V7tRuQ3pfenmeWnqvQeQRK/AQPXfM8FZzb5UuYMPwnQ2EjUKkArwNNisBYypikSPwLbQZ4TUitK+
2Llbt1Pi8NLY1DiYpV8+SzM2TgGNhmgEo1l6HdV8HPib8dHg1OYhQJBStQXFUxfZXrzHcsyrQB9q
xV4GdLqe6HtX9VAMyLj/F+kFYzAmqlLD4wIXgJh9qHQs2IcuPu24K3LjOhdLjJHfKQ6a8UqwBGmS
TYiLDrnCwnVHgR0TnZ4H9EJCt0vbybKFCTilVfCH9XQtvrhATjMKDAuYmfalGF2o+LnRGbyQAf2S
o7XsTVhRcTsvXZPmNDtsMRZUWRbTAhngmrRa4KVebktbvH76PHZfrViOAPFYvHPIyicXN74yyE/z
zjkzOqsTmyZpWy8k42hvhpUDr+X3UhpiVwIwZXvWhBKhMw1KoiE7vp0rd4FlOICs5EjH0xle/Dd+
4faicGf3yIpMNHx4kS3HCDdsW1L4dh666wfbDOT4pjYv3m7gUguztAM5qNLOfCsHAzJVUvTl288w
GQYmoeeUmPb576vn8QoBpzIlN6BkKaySr6aNZB0TPDCyXGYkogJcqTgVnp9sOSrBqwYD04RiqxZN
Oyxs/WOG3mvgv+o/yLdNfpQoZp/4XOcUxcmdS5jXzIe/GH5zHAuNHXApfYk9GOqtHMQU0jdF1IUH
CN6NmD4TLRi6GPgUstwodjKejopSSIn3qg/dCDjq96OKl1xhOjWSZA3FFbJ9mYRd4rEgmtsqMkfD
BqAfH67I7pO1HXlygNJkvcI4TyDVyibr6FcAkNWrT7vbZSeto+3prqjesHnsgb2gy4StlCxcyqRu
TIPSRKzD77XHAxQBC3WRrhio617Hbx0wmM19AHvC9b8jOVzsLOYWOXU7TTjbzmSk2Ir/uWJv8uTb
7VbVWUSQo4GEzAntRD9RQNnihGLIM1M3scSOYfD+dM1kIL4nErJEWA2ub6zFFqocJdTmOqGHTkz8
4Ro61US7ZFhrUhiuilG1dBQA7ZoV6qbgim4GJ3FVhp9D2C06zM6tJVz+1b+XHpCBqQth83EhKXkK
fLNEZR+JQ5NaElbOn+HYSnFbDS+EjX6jUYB+8t+qVN8ru/Sq0pXwB8KP+3aoJ94Ejibw4N4loFVp
pEZg27in+vKRH80tbY0fGvY3SfxUa8FqHz1vNla0Iv4VfcSyPnRnmEvshgqJMK1LlIG4abQONRTu
L0FdYb2eeae5luXn1ov10/5IwpJvnQz0aD8VaYS0A6eL6R+ABh5Q4tW6Nnwn3vy7sS0E9kwODcqw
B0095Vl0714QxCYUp1Qz6fkMbDePHxKeLPRPqULZFMwfEygOBcfsMC4s/0Q1PV0W+teogA8vfajv
vd+pSeqw+EunjAaQ2uHMl4Y1xUSTvdwuTqtLgEko4wcnkoYnt9kxgL2XYWspShSbcFcJ6rnZ3pJF
JBWORVlCVCANr8MNco0/smdQcLO+Pn3Z9/4N8cu73j8AHO7M5g7p8ftui3ew6VW+wn4NBz4UZbJw
J8OM1q39PXzPbkYYiT6nf0BlYGgiuANpvNnJVxU2J3qZSVKge5sx3LWBmaT4w6MDDtccgruO996t
BdIsXQyaT68cafE5pLbtWtPfIwpr+8xCwF/B7HzcOewi4cbknhGl4wAnQaYO91gzaW0sS2be7hQF
HuPTIBPmu8TEnmz9jkyn1VfxDptVFZ032PUcS3FekG4G1ysfk9h4DFeDt79AxY7NHtQ66MMkbulD
Z4hyzya2mhJ7m8ptZrEipywEYNQIPug4OkxoBt6jEaInlLsPp6Hq0mKHt1mHcHpuLmgqT+i6gOSL
uingPzMGnqPOjVNxsfk5+oBOCRMsVi43WCdxN+0qeF5YO6Vd2SZ8WSFSGfwjaMCM7/oZ3sjMj5cw
cjMvjVk+oJ4FglLYuH4eG5rAdeVoWa/O5hmcCJkAAlvvbo8N4smyeYRXXGWOAFmjWLLFi1gTM2yX
kvPeg1ozPfO9jtshZwSDTxYdx1No1L/X2SVVy0nxWRZS2NPPsMhsLjH8EAVkeQw5IykU3RZuWNAB
CuvORxxU8GoEwoVk5W2xg/8yvPsDr8MJj836+abfL7G61UwjaW5EzRL16FVGmgoXctX4ZRzmmLDe
4UIyAfkpd4B9XUnKRu6T3vPeLAdrzaOoxj/wFqCZQtBPblxiujw3D27HOv7qqNFYGCMtjX5jVuNq
l3S+z96aSUs2HbbHWso5iBMFz8D/8ScgOZlq1hApQXKCj3G/dtpm0zxU2L8udWKd4mhUGxnc7Poa
zI3NAfOz2JIwl3XrYuCQVvq4ZkolUdsj6G+M8w93s92QUbLHaqQ2fZej6orMnSWdP/uP0Gx+Q5iu
Y0wLwH2bSO5eSBPKmMhkVbZ9H6zzO5FfzPEf0FxZCW918PBfDn8ixGb/qjVJ1tzn9ZDo0KIaFhMf
l/2WIwG62hwGKLJk6GrPNUqwwHWYtaBaWTJqay+Y+TrfgzTf8qFxXQbbIpYOy2qUZSY50cIxNVfF
obIHKUXmItaNo2pAChq2qHS9ziqKuvgP7fy0/22wlbXQ3DlatdjDIGx+QsPm95exVYFNdUXpfAGa
/t0FiCdT/3XytglGPe7MfoFDmadY4Xc2CoVaLoxxtZStHKdhr2H2crj9OB1fifm0SHNqdHZxC2h7
EXjrwYDN0YwPrTB6/NAGqUdJy5aHFscE8+gk5QVTEaPPmnyTmPWHlajsCVp/PJ15A1e8ppzmFoK5
0PN9Tt+BFncYmTFyYlpFhR8kri2bB6TUz5oPW6dknp5nOiOmfDsWF+57s2V8NSXCJmlhgs3geuu/
8WQGFOri9CPtVIfc04+AYVcmSwYpu7vQ8mrGyGJpAhmMlf18RqguGqPfKPCQuSR6r5j6tRptFZ7F
pNsapC1CaJEFTTvEV0jHNg48YJMdPa0v0lxDy+Ip7OgZjUku8FWI1Ubtk45EBjVXNvx72+ppofTx
YrLAPqZYKLD4ngJe53MMu/8mt+7og1BxV4/7QPeodKZaxlmryr3Nj/3JY63mUOMMRuo6QniBtxPY
i8KGVtEJEBn7XR7Zb7it1l3QV3Su/k7sJ6+Kp1e6ORrl5u71job0N/757gJXsBs8udzqp1ieLXsp
vTdJ+GIOFtUq3OkSQtkIVAGTR4QKgSY9karUO3uN2ZkOVplegkOPcRWQlQa2e0tMMQ8xR+e/S2mK
YiG/I1/TIRX+pePtYR2IdgfvaQCrY4nF+tj/8O+xNgLNT153Hdb1mY3E3Xkq27/KGQZRs0T4iBiF
pybBboBs2uM3dlNpDDoxbYypACX4flM5Cw3+zOMtKkh/lNlonVbBQIFnAQDlSgHwQ2aAw/ZujaNp
+PpHNZbGEm+yUlSVdfONJM5vFebWybR/AGPqU0xObwNoEprnhQ8RIeSUwLReGU3CJ07vLaigFZ8Q
d+QaiJftQ8GPIvXlnyY6n5Usw5XyyD5oqAK8EpwgcRR99mjMi/msojAPJ8VIHBf3yYirkRokRsuV
r2xcWpM9yw8eDGr5nrT8dxNd3z2a6YGpe9jShgJZ4MRZ1plJF3frfuqlY7d4KudGUpf3LITLCHDQ
zAc/v/tR5vxVaOPQ8qMagI1Y85HKnJurxHvsK8coy1AmyZpbLroCbBJRLZJomNoB+0WjT8vQD2Ph
Z3lC6GC1Lj/5M6EXxgSwk5qOacsj0z5WKJ0sz8+4gP71/pT/kcQyRFhkjkhL/7vAAldDuysDKnLD
bbrtUFr6Ywt/rxOBJF0CktRboNoeqcRRWUs18mHHUIR2GLBw2EVMfb3X0bBTs22/9dfhp/Df/FMR
dWvFCgpAj/JAHEq6XPQl5rKlSeo5j7MHyt1Y51kNTFm9RSN1oo5FWEXLBtDBoszsGop3W5grIWs4
up78+m4ZmWCgTnrE0asPNV/yPlVgHrXTade6vT6ubl4yvecIF9p3o9DGRbvZfFjSegymSU9RfVPG
lLdj5vsvj/3qFT2WecaZjPt4iZ0jHDLyQfEIP5e/R2VlBkk/Y96mB8h1gEiz2LMqnBDZGoAUbNp6
Igqhz7OSDWwkDMiYr+JgyvT1fO5G8yPGF9It7EKSd5VSOJDujVvCP4Qyu425ZnyTUYzdTbFMib3T
r5sL0U2nLOCQK00BUHTNBhbxKkWXEQmtRpu0dOmHOhninhzBBsKRImPMSEmM6HVuqZToOMqJFvH3
qgtBSUDPR86ITHt5ZxDhWL28oN/81HmeTqeiCQNs/tf15igG+ZB3oOK5rdX0Pt/c+JeEWisqzCsv
rdEU8ZLrgqUA+3aViCAi3PYRSvecPFz4UjtTuYKC/XKIRTsft6p9NO5sRyxD61n0mMBSkWDTa4aw
QwC4Bgq5ZHDlLPQC3hnfNGHHfpMMDxDXTZ2k0EiX1j3Whkjpf/rpfMAQVtsuWqE5Gep1dJqTYEDi
8w1k78wJnH/MiMdzMmYpYGidtG4cCQIjq00WdyXvS5iUdc2ZoeUPZfGfY3R139T/ODluOs7mG6gY
JIZLcWKx6ue+YVH1OAOqchI+gokN1fdFjbtfsYbXxw/ifcyF5CqrHbS6u/yZLS5HqDCTjYFJn/5M
E3oqy0UCUDvqNB0xaAJ+taMVrEJsd5CTwS7ufWzrAyRUOLj0poa8e/Ls2bNMdN6lw+12rjTv8uf9
HSy3C1pHkEvlQjKkxNrPwAanP+jkLit05Xm2FDHyB4klCSVb/kDeELldBQqgo4ZJQXDkLRwH85RK
O3LO2mARget3cB24UbAJo+QKvObJeDCaVWeXO5aAeO7llBPhfFlk2aD9qdaEq8jvD0+gIqDvC7OF
MgLs17kYpn8DOWv7UyRmz2wEr9IHRi4KjVdPNmXoe2/kR9CqE+1qD6YpXFPMw0wejhy7i/zD0clf
v9k94hkdUVi5L6Rn7IfIMgQxdu4yeQfzxNmSBM0yGUVHG1i4dOIRz9tE52QlKG0twzihDHiUkqGH
eTd0Li8iXWeUWNAVlK6arP74XkgjcEnW3VfVwW7bg+tqthxFfu0ez7zc9lfkCEx+YIUNsQauBWXh
59cmOTykpdA2o9PIQpH53GKZoyG9sCd9qG7oBw/qO93J0XgFp8HuShflSZUl1gjdxglIdkxU2VtM
r+83Y9Eq73epykTMpbpbl1/47zKQVjkzmsQDi3gLRV4Vu5p+tozV9XldRyZ5M9v1tnkAGDOVJ6vW
yk1fwzFMVmKRn3Tojcg3630PzX3wNc7Ta8J3WBsP7twkVzsb813IbHUF97THfo+JhL9jclTsadWF
6dwAYtWPvkNddsJKCB76ZIEEdSaDVnvF3SM6safwaXrNkaV0I151vtFxf1XYhzUoK9Vi5OW16Wa4
efExlv7PSHsQ3zEQ9/lLtEjOsnSjQuTiKX83s7y7uKd9GUp0DHS9kdNPYiyMkNC27F0JVALnhiXb
Xw2XP1DycLFQU8B9NxGhkyobJU0+wf0MuU6uwl5O2tjEcLXTVqKwPBI9WyTayORvKi6id+7levs7
O1M4VmbFta6dRHH0wRcrSVFg68suS9ThipK8CeiQ16JXJa5GbM7Ig5hpX4hFdtvoWQxSp7crZObh
QoOmkOWKpHgTp7x3wIZnmG4iH7CPhf52t/6BXC3IpOMAaK400sZjC1IPEvGqtrFQLi1anUF5A4VU
f467sp9Nb75VWc0kEIhZJZbLRWIDcO6SRGKPI7X58FRu8W8qPP9m62oX+iHr9Ca0sNiOOqpRQ3gV
uDo5QMSzWNR9JL6UO2gfaAZyxvncKte9BdAqCMULA4Em/nwbeaeArW5CSCf/HQb0qiuQ4A2IFV9O
pvxbsseqtlSU9SIfBAMHvhEYLp1bJmCb/WhaRcKFiH2tJCT7a1cQP4E9tRO6jVzEAYcrmXvpLAWa
Ub4CbUAbCU6JTCjt12zYp51vih7TwkSVdNI6GoheNb8ISh9TSo8e24P9kjhIvYKpVvl7xs4W46lP
lyp/6hrlCL6N/xHITrm7S5N/hhwRlqjclhs4aVjzpDCeZBGP21yzDA8U9xWAOKBfZHamhIZPuXrN
nqS+CWqKs8sAR99e8234e6MKQ7I9t9kEmbuewUmKfFYb0yeNbzKc0guMtaumYQZvwEyz0TFgo819
s0w1DiNxpeThun7FTipXUxky5T92eP7PEUGHqs+k8kvcYrsxmnjTBq/fjVhhfk4SzQ+vIxzkY0P+
Ndy/MrSh9Iflk9ssGlF/3g4Z7MIzkiNOpqE6A3b+fxwB0l/Oh0VymTZSRyqqR4P6tRabye6oUvVo
8Af2VRULj1KOAzJ4NhuqudNr/W8u+QHUA1ILyQM54zYCPxEziixFIpVhGKR2j2JFlOGkBrhQhIDS
JANkUr+OEZuIw/5XmPYeR5DZfMV8towosLJOH9vOZfxgq+207s8r9BNqK36DkQd7k3hvFtGMr3yn
W0b8sC2I1a7Av39v9j5ZHCCCXCRHV0NLAO5H+X2GnPsWzidOMutMTDwakJYvQm+yTcGFlMWjIW5v
Qtzxh2CwJT7qDcDlB/MmWFmh+hO4pNf42DybrBgotTHHsfteoA0U05VodgkXHotkXZ36WpFUEfOe
OQEeiluJlEARWmCFYkCijZLBO/tj+hMHakiA1uCt411SoN0Sh1n1HdcwwexRiNrSXJPULH4sH7Cd
uhD8guBOo2yGIahRRqpmo/yrGlxz1RQJFCwHNQS6lfLPenS4tWI0dH0v9WyEwS/9mxK5Ca1pB9Qp
/vSdqoYPVF5LqBvDvxD6N/50O9VLgfrnYpikKyhd4/UBvm0x14GpSRmaSpcN1dR5V7PADz2/WR6u
qEchWUAuBe9W66i3xQnumJA1V4LHOgXzdDrpReq9eJtgfA4+B8hQgOI39HDkZrwe7EuDL4oxBBCX
SbyMwEfqstzVvXoOorDtR6DNNTVdLWwaJRRxJxZ1rHXUgM0DaSDDk5yc8+BX6joW5/zAn/7EZqdK
q2MeUuIuss8sK2+z78I/1pFdKDLCN9dqaw1CqqtgV0lOcdnvQ429cg8CwPbDttr5knuJe50M/cIR
RJKt9751vicepqnNnw0APPzKZxomH3tgK1kqs8ohm7YaYxE+Ad/o0H+lVyZivocVlqWMnePs+x/w
/4xy86o7vvO+nmWtyaXsWr2wuT4L3NGFcj2N19tbo/JRmt3Xn2OHYOAzevXnG0uTNqllYZf8T0GM
26iUSGK1gEeu1vGysboZ+csEBlpIUaoNGK6y9Vcy5krD4zCotkTniMdSlidrUVzxRISNkLFhtHk2
WsEh7Fieh8Q+aKW2GE4k5kUe9VMuM4gFgL/kjKgWPb4A+SB11jo40nbQOGbT3E0hF3MCC2tU8qN4
ox1LVGvEFQ+WrsSPOmkcTk/8S8r2uEvTSDhslW8+j6J6IpMZcHI0Blk+CgKG1cn13I/uB3JDjRFC
thufQUuWAXj9OhpFjDCGef2+LEpn8o1EScZKWt91J7rfSXzdymNlA2aNiFTdhGjWxlBKS16tvZ12
+g0Etpocu6S9moui9appJpr8OjziTz2FP5of9zaRSoDlbP2SBE6fB0UrT9jrbEgbNG80m9alZb6D
azeDaZPEjJB5jU3oSQiKo3rkKEZ6Zu9rAr9ek3TWNSOusnROMOHY/B1ZR7KcerafjNmsjx6+z0Q6
z3Yy2zgIxdNaR5TJMEWGaQ0Lg6ziAtTizn28n24OeznLRcvyD0LmFQlBUG/ES00SikZiWMHLO8Nv
p/F6qGLQGlJ7vI1Ko5KrHGV49F9W32uzGda3dl4sPxh7oBDim/yBYccMMdeQfU2BHICXVi9q5M3R
3RUhTmdyy+wuvfWg4thOP8yLoqQlR6NPf39sZSiLn531AHcPLAlM8+FkGrcH5UXObGFhgUqG1NG+
NsF8GheLXFS8HiTAp5AfM1oAWMAkxOpgOmfYosBnI+0ar67wNIgYgD2pSPXIIIf+tC8shA7d+sHc
d5oaunxHJdDDUGnG0QxJrhZZs1dvprYnJShNxLHsQzZW/QY8p5yVf6HnmT4AzlX59p6TxkWVPhh2
nkZmqgdADpv/Vl48y7E0vepT356OPmmz0MO0Lve00MRD+6LrbUy9AUYfWka6H/6ZUAP+D5pnqiTl
+zthBcFZt4jt9BGy4Jmh3vRg3KuTsQbuHhvzFWdbZ0ssSuxSWqOfeQ97GXAU8fdZNwwTrg7Sfl5S
8jsZvZyy6I7kAmNZUCAVPLOUP8K0D4hM7vY3L4VAERXg1Yo5jUwVjiKDkDJyXylZx9G9O/ugID8x
tvmmrK2201iQnpsy5WQ6Xf9piCK2pGttea484JFe7csc1mrFccorVGB58Nsgpw1nrnIebGiboD+v
ruvoiI2M5Yav3r6dpvK4ZZGgVtiG136wjtryyY5LObO9MzeSc+GOe7s/qB4hUy1vdfHwdp18QKbE
zdmffjYJKq4VMi+VWGN9Whjw8q6b8KweMShB4+Ya0WCuuvG/6q44/Nzphc2VuBcEN0F1zsWTgLcX
HNffoJYHWL6JeZhbNudVo37ZFoxp72+qc+7yU8r238m4/gdlBNeJtUIRYBW5wkwwO/pFOmD5g/5s
hDIIdw+B+1lflPFHFwYtoSnDi8cFIA7o64GiH3F+fEq9kz32uIPe2jEx/qatD2L4K/w5eqwyQ7ni
StiYgr77QYOgjaF9PpGKYJpr91IsIDZZnMDAD3vfCEluihrdSvCdodexs4S5Eb4kTG/XoMLXIYBI
ac8dSxNW1H/z89MMuOdxlP75IvZmHB52q7fpWxAycdqv+Zm7kNlKBFqc5HZq17Ua+tLV0VUuzdk+
GFU+XeeKIh7EpLWjYpMV9CqOO6hTwg3DHhaMF5YBMIjwdVAKMwWCLbQ9Kiv5EJy/t2onmHVTEHtU
RTBv17LgxakZAxwLvnv19LjBM3rfAjWFTa8/eNKisu5Eehh7cN7dZa0g/MHCakJOmMw/1YKOyIi2
GVLnstXFM8fJDcLnE88EZ4+HOQnEasHxf4Y7U3KscdFhPzPXGXYwTYEOqy/4VLtHLCpxadRjmjP6
deFU3uzYemuzovKoEUc+OWFazPa9o9AmoZ9da+9JumkqiolpSrtJ+cuc6XGf/UEPmJepFx56Xt55
FJms+zHfN+EJjc4FmblYHlqNfxhRv+nX2rLTROlMgn4eMopjjTRRm/GapQlhhM+Ak6Eh9xjZZpTG
hlyZ324VCevG3WRDaPjscDBa9K5wYNXvTg7fYKLcPHIZN/5V9QGr7W25Kf6xFc2FLhG8XI+R0EE4
5bL3F6VhbIPUR5HsBG4Rj1h5imI5E/evABhpJIQvs95ZM7D8KsuCnR4lHVn5vhSXDH2vgKmgf+x9
joaMp2dyHQi4egzoLwPNk1DMIJbzkWv0FKXOx/LtbsJX8qRoGFP5K6Iquch0ap4s8NHzXLI9zEmI
iHhvy/36a/HGP/HPGqCoFqy8G8BZqjIPuKtnwOQH8nv1nxPur0LAYoHF4wM5oE0Db9ebohClTZ7D
NjSd5/wMTXpsHckNAh/ztRFzZqjpvNCjPdUOaI+a5Ec8C7pjFbHELL1E6txqnKShYP2o1hnJve8N
RH9yMcrmsf3uZSC6Sb85j2nqRF/iL93elEA5qVqs8VXERuabVs3w5NFjlVixm6vtZ4ZExRLK/1Jk
g9O9uGpZu6r3f7vrum3xYXzbs06rtwI247fORG9i1Sv0yxr2YoepG5ozzmV3z3exaojgAyojhdxQ
lfniQNWWQ2D01n4F/kyIn3qQ9VVA0cJkfu1aAxjONOn9CTJkkGT9qU+x6KC87MxZFVh8Ru7tEvJW
G093vtUzWFF66a/M4YT5RWZN5dWPatcU4iKhS4On+nj309fIzmosvfWs2udwQ0Jyq3mMnNhsaBpy
gReaCWFfTB0/cGEe/4ylKR40jUGoHOlW6WhkN8P9gEKHiH7vdAJI1e0WS0Hwu9DMlIZFcK6kvxnz
+GBbK+3RyzdDtvt7jnJBvdVQn97fs5x4yLZNqBtP0larORmtIAg4L9144HOH/x21j9yaECdVNB1R
j9Zitru2mcHMDVT2BPJudIkRjikAx+UPgM2V/z/XiRZEfi9ousQfIbWmHaGWwQL0L032ww0x9qsh
C2760kA/uqF/lxMCJ5iKwrtDu78H/rpwFljttp3AsG2SqDeILUS5XnndKOoxK553WJ10oPw2WA9B
gULpCOKlEsbiNG50m0IhO3cwbGtx4j+2xFLtc8imt3fmQUupwDAQ4SU4sUDZYZwGGeXxJbstvCeJ
Hy3GgTZJmRgLdvDJHS9L7sMwZ9zLA+vj8doSoRbkGnpV2HpCa3IePzexGyC1pzrzYlI1swgdH1Ka
3g0QceankvxDDrwAwCSy0r/528jybnL3U5CeUSHDFSxwuo73zi/GJcNDSYg8HVhWvoOpHEZ9UM6u
aBoIp7IIygPj8QEBygYJx+puZsoQb9zz+m8jFYftL4D3ODDPXgKSXM6HCmVYMLscoYRUcAxg5tJK
xJ92OzNThfiorl+LNAf4ujTf3asWnIAOqLkwTgzgG6wF8K4VDNANTWgvRNmAAUk5oByEZE3gSl09
YmC3D0niYbx++cP2nQqkV6V7Gt1IalOka0rsdLXPrmm1jO0OR5UtoeN6n/fw7IfE9eQ1Izq12tZF
z2lIyOhN42H7OWcOA4+uS9izwKLAok03n62ePD2y8ypdwmwSrnJ5pyjyiuiiCKZqGjcKtLXS+6Xj
O3L01mV3ri4bU7+n6+V4K+0T13QjhVA8kbEdHRjIc5OgQBGlBZi+8nQ9Y0J0a8WqeCCVkKJ8ovpk
IjwixJ0d5oWsk/cP4IHs5sPivANXfQZky8KRaXdEo2bc9sHX1gUVbfrNIlk6OtRUqvHc9eIHrcjJ
0+e0RfuHZ+sxC8KcwHjtBY/CupyukhLc8knH9EGXO1RKUcCv0j2xknbWmVtW8+xr0E/5RDH4/F6n
qgk//3zLsOEQsIKFPHVZ05X+63PP3B43O8VP171COS4ulYr/dq+tujHuggOhvE+GuJrV/gf2PFE3
NlinMHyjPlfBDSr92OgUfZPRsxML6EF3NmTKXTMRiCkmm+X5PqM/Gy0p+CzdrkC5+xet7f06kvOj
ubCguLZG5m0iKv8hXad/8FiYHq3J/YsL+bc0E2yiSSeeRSvk2w3zhEmw/jGQOvR6kasWrExXx8HO
WfNLMCxCE+O1XCY18X3Irmy9jgXKIfmd6raVdobVdm/EuLgOKU8wvNCz6fPGf+JIleTi2LLhVT9w
fL67gFCQiCXXjv8ZSB0AlybxGrriuVB9ljxqU41wSzBZP72Wxr7LCdvdM40EuGDDK/8NyCfGVVGh
Zdcs84QnoPW7kRtIYPyXJmpg/CCBD1qvcqwf0J9p9233guU0q/RRbEOxEG47BJj6PwVcZrIRXZa9
pNQ3jEbet4bFCqBLmU2j+u2iLL1IPrbN3hHigWt82N7lcM/eZXagqgGTVrw+z3ghlQH78oX5y2ZS
9gPkQlG0ItF02urDfaP5askNBo5f6wwGAhe78KQ2u6r9Yp5jDpgDKbEcui97bIpDuvUTv4vraa8M
QPC0+C4bJkjk0ZBK0GVj/IsbqHP2JAOiT0xFvhQglolk8G55OHoy06LcTXzottMvDKG+Y2r52VAf
UW1jRPANb9u8E+q/Ry+4cF5Yd61nu1v9Tcudmfc6v4Sqfb9G4tVAeU32QNQejYnHDdxl7rFUy94C
8LljqZSCOdooPbnFpXoLNyvU/nrjTBskrKfsC1qJixH6hxOcY6411opcNe3KMZz7bma4znL2UuNj
SaAEpDDiZ2LExWYBntl1J4TkBS5EmEinK8fzxq1Z3Q12R4CejDfhfZmAR2QPLRHY69hexodNHOJe
ZDKTLxSlsQSrn0rbQXCv6kOJtMA/HyUOJNjfulyiWk1KlERmXOmUjfd/vZWEiHY1xXZro7aaxsrM
aige3t2xP3GERIfCpU3ygLpnCuXrolQxCPDrHUkxxXmGoCYoTb+Tbi1Dv4cjXuJKzEjo9NEHtSLA
xCjRIsyOtF30gqUKvKPcJjQ3BKrZjJT0j4je0XLmisLBbKpCzzQ+ajm7BX23jAq5HOdUx768tpTL
N1uYWE5wclr3r70xEIbZ/EQ6wgSjPS/XnDK9zCDCjgR8MtE9jUfncbMCVvrxfIQ5K/lkPtyZwoME
KypcQFOCX1pwsJvJZGLkB18jVEdk8n99WskPxFW65Qsy1YPIH0KlY43epi2aUUaWFqLbvvln3mMq
rmd4KehUvoCmgNpL9Cboai5Fz1a//ekaX/8x1KVEQ0Oz0CWviJkhG1GdxBwt6wo6eI8C2gcFoRQL
B2u2CC8X92AfVDci29QeIqajoNEG84Cs0qCFauX9X+UViIpq/8tpk2z7NvC6dUgQsE0KT7gN3Mmv
ePRhYaOOleiyKtvWcDF++ALvLNgO7jjGYXn8CPzEAqnMlGTg/DDS1T24eTnLuW81Whnm25xzFZKj
HX6kfSbFAkrbmUN+DDjjprZMVDnCVSLBhP48+9OEjRPmNO8RYzjYvT+cDhG0ZEaxx0iW0hdzv8Hz
gyGYL/hvpeTANonQUcOGW4vUmDa09qwrZN6hJiHbt1SaCPdd8lQowmP0xetIt+Asw00SsYM0mn7A
VwW0MQ2hBfi1ZQ2cCWlpwJFXupOxa27IJe83ppTaauOjZhlXX2zz9gBPYDmBtQXimvP7h/SNawog
WWgiqOz0+NcsZMxt+Mvq5gY8FjM6ZGR11sgXl3Jc9u5xSL+WxQD8e4rbeu94fs2y88rZPV/aOpQ2
RcnbjU05kpv8hPSFXqKpCazopqxynjWRDBSK5tCC6AXkx/slO34U0JQJMrdJmYvOPkCz3K7KqNYU
ShfPlB57BcQBZQ1J63JgQYq3buc0KY10yjujP2TEuZnilQHKIEatdufqm9JmzpjffEETGfNd2irH
2S4SUXAMXbON8QTGDA2PsI5SW/5lrPl8JXo7VaVft7SuBf40BSuwV1kqGrq8LQdr+HwV8dxPGhUH
P0/v44IfqIXfWqcBZo5ScpZYVY1hNBQSYt8sit2cRcUjECM6HHdJdWD0p5rl8gL+1P+HAj9RuVPS
GURrOY3peJbVabe5hVzSSk/HlYoGMSAfNbdlkfpkyZy6nOz5kemz6fBS9NreFotVDGwoLMg93Fnj
gPSiyHRx7SO4WnnoVZr5uaymzQQS9pi8R3A8VOo9THx+yvQH9eVD/1rD0HkfVog+7NYTvmJEc7X9
uPzNjOBglIgCpkTzNYFK1bkejX86A27QYqMFAprYPqd0aNLl9gkQtAfcfzGJva0oMzpf8bRAXWnQ
tP8Rqbv9m1qz3T7wQTTxfRctZPJvO9BaqU5BBjk15PKs0LRo/Alclll4ruXTIk8PxXHZTY3s17xE
s/FfZmlPN8VQGf/UfTED6iqEXm5reGcykBNGj1uNr5tIf2mfZqfYM8mbM/xipHW0zD5ykxF/oAjn
rIJj2MfRcqgMkWfIHpW6z8iKFJlL5aSvK2DCEJhgPJ/YFxhUxtIb+lh4PYnwAHcFQBQ6dhHMHiu+
al1QnQK62TJjmhdBKHp0rmGFvNgirDPf9JSCP/SX05D2k7w2cp8Uy0PdW1p3FBflH1ssTqj8RVTl
qd6BB9HCEQOLJwDNaDZQsH/fz5Wfg+2Wwp0RzI0tJOT8qNHMIqHOSmJ8xHbs4VrGXAAn1Q5VC+8p
DGZnV7f/lyomXg8MYSqvFvaQ2/BTd1L+q9Hf8FDqsdZZlkbvB2/0n6k9suwvToW6b7e+D9xew+DL
B71mGawvpKPX7AiTUHcpxsKMWqmBCb24/899xKL53C4p8McqPYVvbzEjzAGp17L4z0uHkkST1ACI
xBsCUGO5aNhoPZDheHrx1ubCbKiFRv3UcPlGWZXkW+Vq/GZoFrhTrXGfKHa2ZJaeTFg/y483DqnI
SideMCAUtp0hppjbRCik45w0VATT28M46qvuPVA8bTTuO4z1JawYvHag0cfe8gfFEom5uOkgTEpX
1GNfx+L4lTjMReNZLBWS6rV5XcMMwFw0YAe5qSKnT3RQS/SDEdPg0g+F4PBcJQGU4LwPUTRo88fB
aL9oRzbJumwr2b1Zeb9ZH8OkepdLQqOk5TtxqetAK5LLwpLj7UGzPEbDxV0wHccoJC5TnX0nGwRm
dHlqsUbzF7jLEhwZMjCDgigHZ/+RApuZGLzQX7tVOi5bsF9vPRVPuQg3NtBs821AcNlRprFjnfPb
DeVfR2ucufIS0OIWiXNCzGQUCXdU0D4JSORjQe3kFjcOBUrFoDZ0xvoFdCTrYYlevlpFJaVbH9dg
sLNxtgmKyvwtWsS4+E2Cexn58dHWtsbo/Z97z12gc2mtEbg7WdoMOAeTJjm2Jcn2Ootbm6E5errq
sPwOSy7BhyInfly83HBomhmcNxJBzXG57nfwZI2aObYQwGZqlddNyJP/qgktMUwY5PlDySDM+o/d
dg2rB8tp732pjoRwhvobGUR1yGSVuEDIjHfEttPXEul03GXOXgqfosC/xFxuJC5iD8XjfIkytElM
PSiIWpapCOqsCq6QjsVe7lUUYwFwAl1BT/TjhD1p559Te/EQZDFQvYVjcHUvAyDwLA9Kpxpu1yE5
SS3sfPOsE1IFNTf7VEnNIit4LvC9JKCGV94FiKfN6WLnkViOxDDKptIiIO2BAoSZbn1IhRKOXGLj
qUhLUX2n+v+1YirXbKMiYmwkQ/HUofvKjYWv4wzF5P7W6ail9sPKO+C2SCpjV1f6jSLdf2QuO1KN
+mDD1T7nDsRms2sRtpT74FUWFpMNYz+PWBwTSNWJedG/kzku6Fkb3g96CpFrDJrR4VeLmryRPd5X
Nj6dAtsoR/uzW52op2UC42Cv94Frj3r1Rxh5QIUeKQkIVTTjsyHo6isKJm6TLGnaFaICrE4Uvec/
f0czyzXxKxC7+HNLYsFfK8P6NXhqKxjW2xX8LTmJnjQK7P+sjZGg6QmovCu4rzqf2trj3MdIjXkx
jsQRNLhMJ9RifG7/Mv0V+fveA6Nm1ejnpJBmGECr+LaYdUchhDiC98c+rReu0V0ksFmhpg2r3urL
gVH/MCyWZoZFcI2MKHBs+7RkGsJU9TqwWmZNP7TbRjkHTV5Lz3iMtwiKBvf6S/C3tFZu8Z3kvaUv
mO24azZTAcm//NFYD1210AXX9xXcSJwR2Hc0aQZIMycZccGE4syPmdLhWKAZMea8UhgQ8bdfcX11
k51CnV0unlTb2oaYTfdU0osdt9YWWrk4VmAPPnH1ZXnIDFdzFD2EgDB0csRmlAjtt3JPQ0WgmzNs
n0nFi8S+dzSKtROstddvAzO6v2M2a8m3KXrOjc3Pp2e/34aXi30D5OSMZ80fZY9g/Qpx39q9h8K8
7nR0KtubVagmEhEIV4gqT7y3xgySaA3EN1MNKKNyrPK9oAK3pZoT2EfHmoOiC+5ZNtZTQE6L/URL
ID4TouEBMVwRWjfAOT1VdjtG73am/0SxRnedeJ6TLCeSsqpw4Wi/QEo2dcHumhwR/KNKUmA4n0AM
GIFwZdYoLPcmRSTfG4stWRsEX7jSIagQ9eavpHW0MDN2juudLnQIYZL8WrTEsrvIHIg1TsQkRCT0
Bc4lLPBv6lf0trbZzLYGDI2swOddERf6yZNYaKenslATp0MHCDDHhsePqHiX8lh1lBd+DgstSWet
RPK72aB0kVA7gMOL43A51/IhvcC1yWoH3qMc5FIPCHbOGDEu4lLrck8lMA/VLCR0iPlsAHP5djGy
dMk1PvIh0n1SyxxG06ROlYkTGCkeAgxgXs0AAR1q75y6KLaSX75xQKPfKeNJK018C+uhG9tvaqOS
u7FRDaa1eBBrtL4Z2HAAFwBXal4loj+v81PPVby7ZI1kiD3ERazzjafDNdFOjdNy5Xd4StfF1AM2
gLwKSrFrjWLOiRgbleYh4uKlKMhi31AS/Q72GYls5vH5nQyKbt9KewKqvJOtmF6fpA2QfDl2oX0s
qo4k4NlYlLpArDxxlPxefDcKjA+US7gEN/1OAD5UTP80805tu1oAZRH7718gQb0IJKHdnQxjrELa
Zk9za9rCcVqYX+czLoXRWTzWSPfjxpaNbjVxY4dxt+toyPkGy2FNIbEUPHcoxXcFeoRSC/uiWxbM
7wAZ3IPxt8esOSlVllEhKyMaNbXNWOHwkAUhsl91FITdOvIqI+ksmAkzfXX0CB6sFp/jJP1OmysF
f+1uK3xbNY8Hg4cdyhavSMVpEzvblHSw9SPyd9lbrZjnPdRqyJ0GyvvjtsgRtxAtRhZ4dNT5L6Pc
hRMtB/nUXJzz3OHMXCSAzsFlJaXxJqFjsfTZR7hTcVGJCyuftkT0qkW5mci2TqbcD6B1YWu7PIJ3
7mCrLQ7Ar51QL2av5GaIUpqaR+jmU/qPwzdFEh1Fyh3OnhUIQtjHs4FBTmKp5nb6Ig7K8DclLWql
3fmhxrrSnkcNfma0opRezjKgYCDTUFkYZZDBP6WthPV/Vay/3/EN4P+nPQljc56mt5upZmsGvMXS
N7LmAbsXv3ayEzPPLokidWnxZXeqAdxDFUEPJSosm3MCr7tP+kcG3kv7JXoVClG48B5Q+5Ypv980
fhYdF52EB2N2cLK1xdTDqgO/rpg4Jfz4Pu+ltBjEGEzauTp3Y4A+1M6ww+nVbgC69Kid71YZPFKo
60kDi2VwTLp9n/f8S0eD04ITICbn+vPVXB+kEvL48Gt12lf6U16AW+TMl40vsStOGg/hyIA3EvfR
fues6h/nRPB/WPUuPxON0uN2T4AywxJ+NYlMXZAbvFbiNpW3Og9JOFsT+n0oxcjeKKRV8SBu3YN4
+vh72m8bLr2i8BajWzndIErVE9dARFNdj9KN/BwZNXIA6qgAXlLhy5Q3nHA8WnIm0IrE37kqlSmq
Z98IdlDoyXltjq5vcwstmQ8CcSFmhm9kHWqplDBLY3WrSozkKCd2eRh5WYDTgpTIWNiEuJxVMLP4
A0MgYfV//FU3Ru0155x99lfMeaEfWek/i9+UCr+4Y97GdaoEsIzyk9HAMoeVgodwuafFmXxmHxhb
lRJvsKStn14Z7QHwT7SLeWaFWEjINEg+g6+hmljWQlwJDDVEx0wUcNc8wc/LpVZBwmQo6W/27Z4W
VfScDSKSIz5ZRW5ZMmdv2tTpnuA4qeDEBRlSKSckTS5CjNpFZ9VjFyYktiZCjeJX9dTsIGFgldx9
hpVB3ShdSu+1YbkCw3Tupb9JJm3t9eIDN/a6Cu9pMz8YrTR3athSHos2jqU3TlsafD8vWvLk907B
VWTDGPIDgd0hBb3HkGd9s3ZxFWWJY2w42uRj6LorPOtrK62jUdR6CVS6+8asAvT0r4laFdHQCLpm
wx0q+0dodznWcEmOJZy4kzQ2KM31sEqGSPLfrHVBiap1taCdFtfjHQgjQxipElKxxK+NRsbVrJJA
yKcgb2Q5EtX2IEJou9hfGYG8BA9aBiRbhB7blFzx6Xs7iYn5QMKVq/PYAcSFJ07sLFv2W9dMuPn2
3hsMdbfnvyMz89SAi0tbRJBeVfMJiwOI1UnECL3++EWbA0vlPQbwRJ2Ty5G5DSVlGOm/8kbvDiu4
YxC47lDWflAUz//Gff0Med+qqh6+we72v44kJS05Ug3S9DOWMnGXHf1P/OvsX2GnoiTcsprslKue
Hc7rENWHmFTWNMrQ6DWfh4LKMy6wD+yz9n6uncFUOrArFGF4ahcPln6GCHN4iDZUCiypusGuBteA
CSJu7Nd+mpymOnfi/Q6SJHm/ipewWl6NGlBhL56OYaqu+9wS5fp8IUXcp05woUF4iSA5gPMFeJs1
ekPa2+snq6F/cEJ1pfBQZqMXEopjuvARVfQB205C0PmAN9ZFBMaLfjgtGJ9fZHoMN9Nl/IuIewY4
xe0tF5XXwYXobqziDalEJgb6ax8QIM/KToM+9qdu363gQ1cJeg/NGeIGSRLDiSkS1yXoXUzYBWWJ
u4Y14QjBkYyZcmlGvXreLkba4iQjtuzbq9ulBZLHq0F1v+2jBh9RmpKz6YzdGML4e/W+bubvGkg5
f/lNe2xhhUJA5Q3cCt1azXmhPiWhCXUvr6ltRHgsFyU9+Pv8yolvwb0m4qSeb/h1/BusC+wfIDjC
Ko+sQxZLpx10MqMmd8TeI+mxYZza98NXN2EfNJwstmHPg6YXaEFF0xJzBVKV87bZqLqvAETbmsGM
mFwdRZci7GcnbyeGR4+losDM9QC5fcEsevskbyVI0MfmPxdPKhg2fNJGo5e6UctWNhSdcwbafY2r
q0rojympzZcYm8lUjkLdbXi++592Onnx6DQ0yn/oS8fZllxZ5hfdAxRT1P5FvYW6+YL9EeVfuzN+
cifAokZ0SQW++ecfIxsNWJ5ciO237QCMVxrxabqlcMgVDRDwXcCnmqlo26dGqP0QH0LGyeFD5FmZ
Sdgb5w2wZ9vVT1wjTx6lPbo6eVFdflsfSssi6kzsVw5MrLS9HAk1n9cTX9l3tsEqIsEyaFd/8u88
m7l+XIzfUBg+XfDHRXeg5u1jZtcQqQUnrLoObyC71Hmo2OXH8iqf2jY9FkQE4yAodYUIk/USOC/t
XPg9ne92BqzQQmJLYJ3F/z0hPk6QbLAC0w4HC5S8w+nW+nVpNNU9/XbKSO9Cyny34DFc785iC0XL
wXXt754hlhmT7CzLt8DIhKTO7h1ptaotelopf+Ndc2Cod7EUWMGgZeeO3F46z4VrR1XpG2dp8oPZ
ZgWl3syN95YJf/5H+kBBeNcYxGuPfZ5trkheMLm3kBjEQwy/1i6OQpbyDg6IgSCPGs52lOI82GEL
P7RJlFOiEvb5AX9cTKH1BSBCy1ASfaW8FN22IyYqvWTsox//95kndhU0FNxXOY9O5+Oz2RI46fvg
BgbOLkPPABlISbmjxzoHYWYH8wrLqrzep8KxUxWGyJ7tLhI2FaIMdbBDOTSMZ1FH9roWux1iFL//
Df6PpYT8OJAIcXxHkNdVdl65cbjn2kNfWhLL5epJcKwalRoWUI11A60/Qw14LO8wslxp5hxn6jX3
LQ2I1Y/mMywDPih5thSCC4obRdSKK97z9Q1eqAM7uKkGV4hSuEMuihTs8Jd7QY26NKKQXP3l/jip
RlwlIXl7JVLOFNHMsp2n+skRapQee30822khVTmqHstxw+A/DJTx9kgkHexGBVMfgqARfoapEe7t
Ra/tDUX7AIECf3ikZyUuDIQ4yi0bPiOsulR2IEccf03NV7NXOr8RMyo7eYt1SmRiys0fJI3wytuR
TA3mJz+Huw6fmzW2mGTOuImsiE7bV2IOtqVhQ4ggq2BqIQEy508tRLp3vxmn24BvXIaY4IybSz5J
KSf2bXZE3vvuXiVUNbeOu0EGOaag0o5cIqr4u35iMZfH6Q3L7XJHRZWJnmq4MddqpB08V4zxJse6
TLAOvC1DGkvy5CM2GDeBQqyspiCVvSh1N5rLqCxlssngft0DKqdMAY3zYk5nq2+TXWZSc1IuFB01
M66uF/+3e5FhO7a8hKXeGzONSCBDYfMwLZtqkfASDPMs4EZIzW6ZcsGJ7ITIsI/YdVecCPQ9NF0g
gSTMUJvajSeTZ3dACn6zsPh0J5yPi2OD9sCjnqGUYDJ3/TGOoSmarHUyM5YK+W2n3bA8uABFJ6AS
GEqRMSxTlZtS4/bwMosFalP/qwLtzhVhigQVaX05zg0e0yyXQDQHAL0HtQ2sJ4LZH6SnCoNEW4y/
H87MupfE0VJ7mv6JaccPB0pEduWkZ67nX/vQU0DomZAMrn1E8VMza9ozdk55+IMH510edOuydeFL
wFL9fX6gOqjgZkcvgLBnIcDw8H9gUra2HK1XZ6rgUJmq2s9wKooVoODq05W/5Rw+FRx63jLhJEyE
nEV9U7TCM9tJ0iFGqqtTp9Q0CXy+NWdrFKOaUKBiazMVZMcca/IgAfqjlT3tZHbvIPL1yPiu3Uom
8hYxOtU74I1CkZWnDHhMskV/FLBHFjGaFFRrrth1Kut+LQnN7iU3gR5P2ZI/7Itiq46NKPeSk8uY
pGD9b3dvAWBqkiB0asdUvE/+DHKyB7XAxmkbTlJxPiRw7qwhKoywSyvDTFgTs09tgy1EOb/5wQnJ
543DAiTup/7mS0QmFH2UoxmJxvIlnRs7yXaR/F1uia69TVOogKpQg2NOLyf8KVTE20hM1b2IZ5Qs
t5S/Y2d3zwjjsnLv8HB1TKdBBGqdTkG4yFJQLjoeVBpEFcrHIFA6tkR7SIngGOJxvEo0gr79zMiO
KSDULXx+lx7Q+P2AzUdVb0g4jG1lcr8Jvut+nAbGr00Fvbd20JEkMBWFHYhIXcZfHFa4jtEF6YpY
p0KHMh6bqJKHCpclGMMmmNU3PPVFKi4geQRZlfXYD7FA4F+4oxef5laJhRL8hcohGlDXn2UVFGYk
148m/UxHffYlYd9e6aIIVpapRmf/sdfKSzOYzqggfJGGJ2ZQm24Yem7ZUSLuvDqSVQvEODtAYSlA
T1XkewEHuhVNJqHLF31qVoCLvyZVPke245vkqGtzf80TtgHRl+PqpyExpfnpVxOuRoOid3i181gG
1L/opfsS56Bhpf3dKinfWEny751POFlpJlnJyx/Rhxe1M9x8+D9wsiixsmrmoYV6U/kZSCCndwQB
cksyIjNXpyRZtX0PZpJpwYnZjK0Xji78vbuNiXXdWZECNOsT2/EV1UpScXwPPukl8ozCOQHFtGQm
D+jnq/neo9lAiuVMhwix/ZmVstfmp+e+PIw2egoD+26Dl4+xz2dc2R1grE36+A0fkL7Wm6SbM2Dj
PjdtcrAeH46Ebg9P5n60/tunBnfb8LJdVj1AnyVtPb+gRgNAVL7nTOU+H+8oJl+bTXwnC95ZRnb7
V2FdWSGEJ0vIFIQuEXG29r/l68K++3CjObSro2xlAQVxgyGAR/ucMXEwsCvX/Ss9XqKz5yaeAG/f
iqRQe4ZSR5Swi7vmWYbfCoZGAp+syB3QpVJXGC+307b9izElMTUM3tUptThury/LiBIAReMUU7RM
AzH25yzeg5tWh4FXRkdygF5gJmH1GvnwwkoL/t1QGP91fcxMAegCIp8wJDs+7IKjjet0mkcNBbzK
NNKbWHUYTasew489+SHutPPYCjU4jQfic3Dg/PTrdIPK38OiNYoD2+qtnqX3BXoOnyNjEccW0pq+
5+wxzlSe/gbk0gEcyqLl0Un+TDX+afK9uk4zMPHF/csnctYHq7FEXa/fZB6XP65ZLWASmktcL2yp
y91WFiBAi/g4JOzh3nq5RSk4V39czXduelQCNA43XIMoAn2ViFaDjaKh7zR6p8qIb60Fdkvz7ypH
tSmZfnHJekVC8NhYcXiG1DDKxxPWJJPYhKKYFl6ecR71ghliL6YsSZCfwnvcqP/FUTYFou0wKOKX
aBsuV0Cre57c8sfamxTrjCZDaw6p/Z5e6V/LSDMmdF2/6vRFARrzMOS+RhFmOc1rZk1up8iMDoNi
p8mpgG2/702DFWocEldIHauY9XdoABBqgbKtJy9wtS7/LEWSYggdrHMWRjqi5xZBDXcTWJONz5Nv
VwLds0NjX+q9r5+AQMiZHiZ0Rzsxg9TvW680uJeEBgaKd7cw7LDzRRINFmO9gxakLXJPxXjhfW70
wgxvqOsTueYcFTNrfT60NY8LQxEOrJ5utRftcB6h6fHOl4IGBPM5VJivYjmA2XxRtP7wvlU7s1dN
8zc4+Gy8/2yf1qNoAHB6uN3+aDqBR1YzVAPizgKbh3cXgLE/OFAvdVNbvODDzxsAbKVA7E9UwLrq
+l+tPg1rfL6Vo894PetoM7GPp17KUpqP1PfXZuW9K0iDNf9+Viu15vcfe4lRm5FF0joBkl52edZm
TG4O7u+9uxAoo+x1YrHGeuOrzBXkVvWASmi8mYmdOfKlJznb+xZ6psHVuD0Ts3iys3YVw5LSSaEx
gJFExAYDI1QlDT5U/f52mhHB6mJCFF828JlGQjkr1TWeZ224Syoa5xySn4I7d9nkvXKPXA127aEC
ISnzhXczjWxtVS8xmdtm0qBy9yLH23BTCqfDm/+0aLV6XLv84O+8h6kZHksEHCBGWdVMypRAktrS
T2Jr6eGrJiLb1s94nk3xL7E+vs073Id7/KblynQOWEHR9ueVWxpE6TINVi21VzFbh47R8+cKKHnw
ApqNocgGcJIjHuaeZmkaacfMdDSRPSI6sfvI4z5ReebeR6YZNjUD7lXN1920EEpwOHCspi0K0PZQ
rVN6hodNCguXvsmLiw9jn1eHqNBa4S+m/kj0zmYKiUhXlSPz2+145d4n/JV50W4LUgLC+wgroz8Z
JSfJfv9deb1cPGmZOztga7qjqxgb/BTj/FWCYwBfMluHh5Ztt6FWItxg19O5X+tqE0BulBPDqyMg
rjXzaiLVbR39oE9PQjDvRgb0kZrWXkyjf9iwvi67RFnUrxJpN+vmOgbaMTZcJ9+Se+Hk/NVOwDPN
RC4Le5oZTAU3YUkXU8unIzDqVxxDeL4AHA+PHvmRb8yiMJFY6vdFW6sur9iJ6QXilf3ZdePdfODl
Kr+mu4Dgz0KD9tHRwoXIiElEpEi4ZlUQEcqEIyOlcf2ATIAwItVz6cxt3c/ddTlVcIfoX/4so8f2
CLngLqo8Kt30SBFOluhI6jNkA+hPdK2Q0eePT1RfwKFPe2v7g7mBPKweUF80weITysA0Z7StBqNi
hGuQNYFTCV4slEuhF2yfSZPx/WYH5hJl8kqIdTTO0qTSRU8/7O2gLMxkexo5OdVcm5SIbnJj2Sfh
1l5ahzI4erZ4VhLZ3ta5zk/I6GOVwFsFRYXZiSVxeOdUvgiQjhNUg3rgyLzwYZ2Krktj6St9CjI6
QNQOBGQIaLPU6ehqCbNtnuKtwtgrdMsDCKXrYjtB2xxLx31NtNT7MzhPyjiKhR05FNzxQkDrYNm5
aqP1deh5x/sXCIQaiS/ei2eFXGCCwNvjwJP1JsMq+H0SoyQeqzuXQiawcoXAmMc26bwdaKwd7/mc
SM+d2BR8hLUIh1PwvUBAB1CCl1sVGK44nWpQp6cQedfx4IKUbVCqn9L+aJL6v9PC5xTMPFe8RXI6
tGoykU+rcODRUocXJNtJAcVNxAaKGh+0u2X8dIOLTrr1QkMC6mc86bA2izbK5KEQ4EU67VlqkB6V
6GyrWZhIgdui1wiXkxJtvlRF8MX16sU2K23Goef0EPPqSXYkCn2JeVkLnylNoebIA+uSpRUQLwXm
2PT7abAr5Iga1++vB9YXhWs0zdqTTnCkkvVA75zQbzl/3t0HVz8sp+Ganrd+x19xuTJ5Jtb0CMCJ
sOBfy739RP+MPRaIBVR+NB48B8gGPyWQtKB4qLZjj6QxSobtnBIeEOs8ZVyhoUU717eFHBxwnJrw
MNAsnc1RQLT/yVOHpn1ILmDr2KMnYOdt40KPDoHZ1gQmLWLXaNDarTU6bU637NX3RQOgN17Qr18z
gIdpMvaVuZSBLtFOuvsCWa6LlWE8lA4HZ9XpIW+I5UrAWVpaF71tRlJEnDFW3+Cx65bIC/vsctNT
U8+E0xs3wCfNpqVT9e4xTUg+eKCP82A24kKAMxnF2O/i+YYCSp15qNdy+1j5/wjJDf0e3VsA1A2G
e9a4pRbdlVaAcEGRf7jID4D2SaAfDr9sf+dn4jlknszrFxI79ro7SZq0HnrjxzS4effoRLNqrTdN
Zg3IsNllllCHtrWzs5msDHE86KeLjtTNUWKiBvoTUVfmCNx8StmYuG/Q/Ba4c5QhEJxqVKMQfXDA
eVKpEdpEPJb8byVHm/1IrIOIXPL/2rDTn2GhriaReFbWEqFpOtHTJjffzXZJ1V6cmFYN33mmCUjP
aF1KNYDoN5VsX+aGk+SZPzijwg3yAr3TIF8owUd0aoKuR2uhSOFqKNsVjx3HvSlbZQVkMmXVrTrF
Nkyj6FrwEp3kya1KelXioPQxo928aqim3E0nj3+levqPuFeKBfP2g9Y3bMBNbxqx90UnsPREG575
nWflpTLO5avb8mlvigNSJjZO1PcvttzyCv/i4p56CZbzFz1DFf+5W56JkYF51QE2k9RY1OJ8Rckg
QK4TMrFRYh0aV36IdiApovy+HHurupvjzafVKAeawHwFOxt5YUONLMAs0rVrXNU7Ue8VxS63ETZ2
7Pq3O0aqsDE5LxTRF9qEGeCpraau4bWw2oHrL8LQJyU1UXczE7Hd2EAynjwRZ2nQJbNjyA3v9NN0
240lDJFuiyRYph/lej0sZdYwJvM0L0aKbzr7/rjvx5xuIYIhQvdPYirA8zJqcZkMKnSPu2OUQojF
P87Y9iTVwGUbHKMQcvknKwCnXfVle7JMJEH1V1RdZbsob5jkIDnH7yp4qn9PqOs8kgNJYbeP+oBt
Y3Gjo0slnciJiwJJuYFvWa1YE/HSQca9ihVS3FWAp+YRGd3y71/tI0FOEJu35lo+Wb5cUt9xBQcp
F7vOrJrgTYbz/Nd2NHDO9UFEj7LigyLWpP6eYiGiklclhfLSTA4WqevaiNWKcLe+nm6rgd7PM+pT
id+8K0JvBIBPRu60tkPg37Y07knjFpPSVhEa5Df3dBS7Zv+ix1W6L11QyEzkLKrdDns9DXqp6baL
fNLD6lnL8c8OK92RLKSOT+FaBwL1hL8+t2JoPEii8LsUc9zAZjtch8XXcZCLwYXnKb0lxeEqJOnn
JsEe+fuBrpel2qWyeVrSF78ibgDHpnzH39K63AFZYgAGpubi3y8Kx95yNkBWu47KWxOvtjxSaCnM
OVxp3Ajvy7J9Te0uAdcNAwWHH6zP8kVrQNcHsMYsvcHUMYUErMihVrYFawq9rm0GgTEr4ABPivZK
Sq4Hs5MIjgBoFVXNuiHib4PNX0dN9cDr3b0MDtnrg4szCKQ6gWdqTBKkHrgx92frXzyWSG1+dg6b
3JX2LfhoUYwQ+nE0o+TVlTMoSypenZr6IzuHQdqOYGDf2SlpD9fiXtMJxpQhhDAFI6GR3zou545D
mzrTLoVZKRZ9WbLQK8GDU+FHbyEYBYk1PRyZptAJNdlTcxA1dVDL5DyWEQJCm9UFfHgvQoYAPdv7
oCYTfF/TvVQBi+JsOj/+N3Tl5DTuf1oUhpBUZ3T5IyJP6HTMxkJGaTuadtjrWZaphAvKRMzGUyiJ
O/LyUsBbp0soUoWgRb/h9+No+ZVvDdIiR20cV8XzaQeiZUmHOgrT4FY+ERhr9o6MdzijL6W55hmg
MWLfGOtKImrmrG8u2KvHfKzBYJ47kY5aTSMrPfUWdS6qNvTkyg7LpwEw4EELk63oYo7ngBtFKdQ/
lSGuFpWZL7EoyBIOPbcx2vEKeHsafojlHZTKXvmzLBVHb7aDw3BpPRRM+gTGTpvi8gtr1tNIS68y
JdJbxsfsJyxInpejAd6GboDMB1LGNYAlxTpFrpffwKU9k99BEqE4Acan19XoNqkbZKZJt4lP8G49
Pr15WVQBy6wpqSUinD5ET5DxRZaDp2rY4jvg9wRRnjd7PUFT5CWpMYnTNrta9Wt+Ha6qeGt9G4tL
y73XHUNTWPKEiMAaMiIT99Y7Tei9RH+UKYazBikH3yw5KtqQs46U5XIx87thFVmyPx65EDT/oyeK
53nTXf1l7UaZDwxQtGJ/O4w6S9x5hi71rPZMJTXFykaQ+ag5JY57avF/h67VfQid1mhZUJMPIKRY
0tQEgUlWKmKTqiVeiPdkUxOxlsLOj714ENKkYq7MuS6Q043bP8+SRLPHaLGzZoRtRo5iWtRSsbin
k7h31JFH/wR2OhkcbUzF66ZxfuH5IDFn55gBRbjOO6ybTakxCtVFPUUdNt9cibFF4QCrMujot7Rm
CoHOf1pL58a4zDyq/6oJ2A1pJKSBKMkh6XvwGjj7nIw0XRFlBN2TrLeNrXRS87Rg0/CXZ0P7ASmR
AzHCVzUarCiPP1hc8DFiy2Wuegnqu2fYFmaKQoBHzvfpd6L7ENe4p6Ca90KkOuEpJU1qgaWdDuAu
5ugiRuephovWNuJLzHageH1yeCrszTdcx0x/n3/0fQ1UznpJ6BP4sq1Jw9v14nF+nQ2waGdmBeAp
adrHQNd/FGyx8cBaWLSFJ5ODiF7Cf+2m3hXQ3fURfAov65YS7XUF89MBM1ElOZViAGNSuWgqZftP
wnVYi7uKgT84i4gPmSyWJYXnWft1YrwcsXBjZ+HblrIik0Y21fK+aJxT8eTPhwLNX9Ij1G8VqS0+
18SmxiasQrVI759b+iI3cxRUVdXXsld6PoU8ds2pGs0cYtY+PjPqGfuFWxXBfhwSkwNZtT2kbDUW
RzMu586IKD9fZ2HfUtIHh5MsF0X/W6TmbVZc34f1g7FzX44ilNiTqfFULvM5R2w63IJG2jm8KVRc
ELKseb4ov1777TwFBD3j7OFH1v/GoqeZ8cC3scQUOYup1xw+ePZVYmYk0K8DorF9ujUKzsv8BNoo
bT57QierAB5fQ9S9fXQvrtDaGLSGbaFs5TdKSaGUxbN5KHJBMrATC+9jPVT6ggkG9qTgRQzfvh/j
MHMoZ/ZPMT0Onmcb17ra+VhVYR6C2xF6GzewFXl/6UtI9xZOwfju4fRN0dY543nVKAyLwwQhAmA3
BIqKUSL18eIXvD1wFAX1bTfVWNmRaFUFuXrcUX2aHSlFEi4RSgF0pR8m6i/x2OA3Ca6uX82BwNv5
YYqQiL93ILFs2BF+Z18YGfXAVsVEdMbLtPJ8lTieL1dgmqMuFEyXkf3f97N+F4BPf75FyB6ht0TW
aSe5XUyMT/1+lFZSvQiq+cH7u7rqIYJ/+MlwzD0k0gqWMezxfw164321ilZhqW4tExuR55WZMPlv
jVyXqQjTz9gVjXijVPI3nNB3ewtvGmNo/ElBMBpjxZU1YJFg9l1mBUX06QZKdX/hFvIaN/Awtf9h
N46gWzPAcw5kyIEA1ZkA0CR6VOzbgo/4Txg8uPcJCKy5qynzYE1o80/B3nyAhSaNtF6LJWF/JWUS
vE0iM+kUGHtdPYppXz+wRCXPEFE2FZku6q36QJn8dqn3b/xVN4m5RW60u9bcV65Fk4pR0uc5CDrF
dnTi+B1g7xMq+cPsb7/sycIK+l9j0DfgFjt2U4S5JRrF8GlYTgUti7agk7sVlq2y/rJh5pgAIieF
DBm/MaE7SlBheW17DseBY7ArgnZ/+N+OvFtZshjVmWlPyhRYFr68m6+PAO8pCbobICOR+3H9QmfY
unNweKR4x5kKmdEAbQWO2RJWdNkTaDIpuYjLnI2vt6IqOgjoX7WmVCu27/XZDHJzN1oE5l405rzJ
xehwZPIFmALRv74D6/6jXqfhAjXAfcN7o89pGN2Gh2ta/Ces1/E7CsQJOk6wXO+fZh9c8e4ZYZ9H
WCWMVvNTLCIiyVqm24SOsQyeXX0H3aOUhcQoFn1MgYT79pLl0ru74CmK8f6vxngzMa1xQt6fzCuC
ShOOS+EAIPB1UZYer873Y1JEyGSi/KZXzwQTy1MFwVHME5qxO3k9u2Thulm0ep5TDPk2V2H8LRmx
fuF9QWdmUcy992b6naefukKzKO6gDIXf7L/oUrKb4ccTemI+7ynEukc0TSEjUGCpjkRWn5fA9BSE
GjoFFb3gw+kPVxJkxOwYs5Ws21gNXlLHGuNGqKxlgq2AW1Y4WjSCj2A61Dak0P8P21dUo1mb3Pu+
/6WLtZwJV2VGMRqmqkergW5+CgkMW1rHs+83MHr5/V5aEtKWaZ7fOVLkPbGNIyjFfFwQIBBFqkla
vDqBIOEF3L7ypZn0oL80cjdw+Cw+nYBEooW/y3pX4M/MY+DXgSZeBhdhaswKi++o8Me++tSZ/jfO
1QM2KXY/Jzn36FV7AtBtTApZctcN2VMGiuFTdFTdBzTdxwrc49zhaEsFNZp10g/s7Tg2nuS94X6s
veXJaaqd6RaIoKHdt5WLvUFy1e8m2pFa2wxjbG76Xchlfe8g2HGm+u8Mk4w4SNTCkp9Mo2ppaTo8
nZowg1srqQ0Ig2KhEuT9OAYQIoPfdJ40ruWdiYqU039yMrMyBIewgoaLmSvgxB3NK/dAnxly+4vn
1wkw7BVZdvc3vbYgM+kM34FL8P7JrJA1nXx6nX17F6i0QfmYqe/nzHWMmk9+iVOdjzXh8vEMgVd8
vtS63JMHzjv9ALYQ/5J9GMiR1UfKhhgSC7kmyqbeU3Mgi/FeQmKOTGCHlRh4Hf6NObE826OvUmIH
cSjb27xC5xKXHBciX1/jB/5lsr4UL8m0Z4AGFR9gFgDM5cUHlQLToPWG449sfHJDa0INEJ1n/0X3
C0yPpMMxKJD6MjICjmBF0bvzd3Bd09AFz/5WyjgW7HeZALvvJ2dXulIbgenUlIzWXLCwaqSf2I8g
AHUtJ8kQqBQIu+Ph2u3pTF/CoEQ2d/MscHRlohAwrUYeQO8+WH3CrxpXdyfV1c9nbi6/WpPykVaD
mm6e8rrrIHc/jT4jaQtJtU/1QcvRexVXN7yAzaYWIrBGfnvzz+lrBpAdoKOdIPPh5fbse8DYHQd6
CzSeQZVKV8MqTN0nIW0gjfggnOg8WGOvDrrZLEIoRqg6wFJUmPZYjsZvAdF8GubQrlbQy6ubDm4y
k2iJnCKGYUQI7gQVCtNwvsiAWTzFLB0+Hl4LNZn/A1mVZuygrj7puDX2kkZcMZDdkQz1HMr3EozN
GzFHrUdkrH9zR9ivnWWDW1bYumps10/651UESU0+kULyfExU3215VZ+u17bKYDWk8tLU2PIjgltx
3qe1P7/SNLgFAfsV7OppYyZtmAuEdWxlW4Yq+ltiw5sgmmAu94rQIoxSBeCqRfNze4SKfwz5gDpx
qQ/1OhDHqswaVVGS60gdGk4+s3pWUCKi5wMG8ewfOt0/CXlJOSCfQwGtCWm1JCie0ltpagiTmoHI
C+57INJZiGw8MSbhbtd4So1vVxOBSK6oewVVLKQViuxWC1YK9BwI1rjpLOFjau8+Sg8pv4ptOZEq
OYn/KSueFwSKgoOm7lNpNwsr13xlVw3XpgD6fuPeuu5cDfnzQNiiHtj86y+NG5aRPnaI1eDBEOya
wldTRnENknwKoOD9bJFpGbv2osZDW2rsem692aDGxesE0I13r4LsaAgx19YbZl6MWvbH2lWtBn2F
FFyBpRaKziuFXn15leQ0MqyDeaHzN+YNDHQP0QBmaTS95WxdbkZB5QSz3VHI5QuRBtg0sOKYEv51
5B+mTYdhvKUSbUhZ1OEy6EnHdt3oGCk/8Jv+F9T8i9SidapckWKJxMAvMF7JuLHk1X8ktxCR2pej
kJ6o2Gv3sZOiNrDi68siANaCQ74wW6HyXdMv9fQf2RzJSEsFNCNns2sFepsHpSCTpexfGI/uXf3p
kUVLTnQg/LTyqaAajDgmTgq7wKEfRyQVwhVxMPtdzGBbqCGQiKylBecS167evBsPRYf7jOb0IoYL
L2ZUli7Sbo9g54be9fi5Ml45PtE/V1HcvGorc1OfJcZF25/RHO3TazzbF8lLusolsyzWpzOCCKfY
7jI3Boj8MZ5j8V3n8AH1VPtpPXw4OnQJSeOLvllwo2YWR6oQMUWDzNIKk4SGHrdAP0dsYZfHnluK
R7YGVY2uUm8rNLMZJHJi8cbRZ2IKc1dSAQKzJr05pJ8+nvR6jUTFjC9kXCpLHK0Eynsj1DysWXng
JlF2RdnbqDbkIKeTVWsKyKQqze2r7+HUfH47Je29t+CaRrRC6nzYBIKGt6rtdtsgTOwWpaZFMe+/
+NsWpPpielvGLJ9u/DhR8ZwZj8YjNUzbl6rXGAP4s4G5fqk/9EayNeTmG08YBJzywA1+ZKyjs+U8
A7Mfp2PZunqaMm4hzZMCVTtHPX7X0N+HK9SvtpDmMyt0CR7KnHLNUwmobrlCm8X82O2YRspO9ab3
BQ6QOelumij0/ClVjASBvFB/jZTDWiRtLnoVM9ZVJViJd+PyptV4bxM9QcJ0Mh7XFUb31UnTZK9a
i5livc3QvPteqKL1CzJXwyItoFWmeBS7TQwUGic6e0waKxB/ZNeM/MFjHNp0Nhkbij/Gh9VoKMbh
OeV0GYgICGqXXANo22CKlBcJKeWLCO6AWq42P/SUATUuhZzJND8p6ggqhqcOiJqsCzMifoUqEdPC
5Is1HxqSQ1LxkpKYcr1lpd2YWikfS+t7yA/xmYXv7IbO2C9/AzsgwVSSSbKsBwOft3Sen+6CDLsP
ZfiVtGSVx66PZc3oJUZDUMvWuw+k7ANBFgfT1RrNfFEqTSlchkn4C7L8800gDTbkz+lPrIZGXSIl
gdmO+Azdx27OBCISQFTa/5TfFRzDwCgZMAgDogYPZCbR3RkcPWRV6cdeV+H+w24EZUxAmZ3r2tmq
DKK7F6U6qFutFSbzbSkKaSmb1jAc4djBIgfmVzRMHneuak2Me977i6tt4G8Av5U6acUOEtHWCm0e
/94DtFmeC1qy484Bf3c8lDna9OtZWh+Gm6s9IvIBV84rpAjKQMFzcP2EcAJ5Z/pxh8iRXhhrzenG
EjSXvion+3knPbmk0fyiA1WLuUuQybqXXv+vIThKNXKikXmtflgw7C35l2fEuNhteWzf3TXRLxun
6M4Vpv4jTB+hTEK+3OjeAFyPBwKDp4WDMDJASlL9kMDT1CIclCpgqHi3dkxV46gncASAAyfn4fz9
O40pNNoz7hARg0jlLYxkMtp+C+l3rebCXRN9KBukPnYqdbG/CNBQsj/6zHD55iJwavdNgK2av0Qr
uuiP3tcjX2jqTci54QaK/ybFGsBcV2GgAOqkP6werq7lC4XE8RcAc0iqb0srYKFGPtEW65tDd8YR
vlStf9lm8ZVwbqtaDny2iX+t5zYIt3T2gaRPsiQebrf2ZdftKQHUAFa08RTkRSAym9qvUvmwNaKV
Ynu9hj6BQnYiDRVZWR5bClKy1jCB080NkNhNqNhP6mNItDamk9utQLe0ehjj+XB4psIfNxiIJVjB
2JYln84go5io5EUG1wkPKJDs7uh+1CCpx5UTkXdxWbTgBp6DNCC32KxfB/LIjg3mK0Y2Ferl9OFJ
KHZsogT7Np6nqodYVMApg6sNYcga0cJzpzpqNbjZ7H/MTPFhDV1b7H3briXNIubhY0uqDngVD7jT
+wEzIs4uAVlXZfYi4bu2k47hDfLxI3rKcUO1ARxuBSjjpc26r9Fq6z2phgS/wL2jySpCk+Kcj/zv
YdoFM4FjJp6vajHGzCIp96ddKmqzxryddnC1rDUxo4SKgYLwLq5clDpJLsWBvEyHlfyD8sU5syPA
aHLO/KDeycWE6cyb/r5pU9J4N7HVFdoWKXmVFuPLFX3iAoDc5bu+kiQ23XOPBJR8kLFGuXvuKfNb
oEBggb80IYA8LuJEJVvpabC066EKVjVTaQ+sccSjVx+Pvanvfu0ALIMJ1XchHvMnOpEisljRr2EL
5euquoGFRLfFTCjCxDES/DPZdplfsgUvZD9D4cKhSQEPZaF5B1Wobf8vriIGVYH4e0OdyfubmiNe
Z9NCMzDmfdPa5l3hWVq3p4T2rLDQG8S5Q+ttcBYh0+vPTHVffD+84ppM+tN9+KLegwl6mDtQjQlT
RWJcmEw5mX4U4d0sKNN33cyT+ou+sGuaORSk4YZJQJkteWHZPTJI/EoUCnMgemmA5QdgSN1trZ+d
ed2SdWvSd0S/B5X3u3TEEnKELRI8rkacU4Y7oUn+zvdc3xeXuz78dCI2yqs7CIiKrE8xtslzGM8V
pbFRdfuj2FGO3EQlticCPhq0QGfhH6FfgTrcwTTDPv2lqbPRWMhbstYOYt1oakTZ56gk5m+gWWAv
C+QoSW7YFinz1KRQLdCS3X1pfjiwFfIRrzM11ts8wCSlJIpe3Auk0D0YiCyCgfs0CdRsoG2xYCzl
sSaXrlV6boioneoAuM/1NJBXGorEZGn+XOFUaeJETeYRyvegHyd9QV8ZyrEo+Vbqu2DDQwwCOzWJ
JZbmy1dY5vVg3G4F3U339Rx0fnImdBKP4swEDQjAsolPch0zBPyPHdW9fVWZZaGKWY/sMbgX5L7y
VqvYo05OQw92F9Hgm00tiYpHtMfuWW5StFY4feJbByRH2BOjsMaMZJj75+O0K5XrsxR1Nip2dWLc
BWK0IEDz2eizNeVVYPswys2W4Uj5mSxB758usXMsERR1c2zCmn0SaREEfxm+NYYobV0u9+OOiZoV
c0TFvh8uPxwrje7mO+z4dniUj41GggckP9E9sP2BKs03iTE064ZoAAna/oHhc0bjM51z2gS3lbeW
oohaEXmN0gDOCydSHbyWPcINyirmjAxCojxMMzUriIevhsQQ+UoYQzY+YEhztmhhxWsrTAH/xHst
FGmUOVfkuUqxAkILKIvzQIlBt40vNafkZXdUAH2362LAALyDfVLkPA3OFLxOAyHMxfDxZ7iNEgYT
CFohR2obnXTb6L2mvivk1lnwfjsHWO/sWgu9QzNCwQAD4cG65pc9YaujAG4t3SL3fUL3M57fiYRF
3ZAwRhouW2jwM2i2Pta7Wyy0Y6YzG+GaAYSSnHfe9Z2fhrsnynNxyGKJX4NzSeThHtpPRDFXm5/Y
5H771iT5fXmBjqX3y/OYIBIRDZ1yDmQWwPyMKOix3q4h1kaV33TEsVj6qS31M1uO+O1GDnoy4v9O
oXftWDpQOkDxAGUXI7zo/W3O2xJ6JqryaCf/Xj+rxybr4ZHf92xXkhA7Ivgl9l4umkNXYQYvTf7u
oMtcBk3wWae/el5dciZ1kbqMQwQ+yjDkwKJmGz7vI9tRtU7TgX4sbsA1vlIhYdT0zGzQLpG6ZPPG
R98EUGuqp/DInBCqPtPKKb4y+GhgvEvrzvIMa6j993lkZDUHBm2Mej8QfwWBXaq9bcsYy2cP65UP
p+QvwkPaGoVgxtZVI7q6QQbpwlX4n/cSsVL3aUr/k9uyWKVWKsSJgbuy6CrF/zJeOKMEw+oyc2Vt
TrqA/u+PmInWJkLtuVwJE5mpLO9BcJQzbCMNUZ1QdDuJ0c65LwUfYyGJn4hBMMKHsnM5rAI4PVPx
LLxvdJhnCOUOGlCNPsAWcODcMjjfGfnu2pahUGz4M3lbKe0RC5iar/fYm3FYNOd0OMg7YDKUII2q
er2FhsUDsH4sAnM+/R3iiukdbACglCKIWt7T4/uXV9qDM8JqnGotMnigkH3deZCzVvQT7TfVuOzP
ocSqUNTzedMcXabaqT6IPE4v5F66v+e8DYbtMoiJH1HEmKcGt7vKMgMIBKq/M0/YS1CL+/hOnzkn
UOqhGwJos0sr74QpbB+jasuWd6SIFetrSXDdkZQQ3XpVHl2f3dukPnooHWB5MV0DHsKsKToFTnvA
iyxbsNNb7GH4wVgRtKo+DPMJHk7wUW2SDYVy1eW+KIB8J+IH93YxNXq/Xrq1+TXSyAvCUjF0r9Qt
oEq+KfmLm8+1Hrqere7MZWxubAMVNF/2/bw5oDpI0nyCS/QmxUi44GQO75XHVd4vwXXJl1GlUd4n
3sMGYVWtFcuuAuS5a+ClzWs49URbWpCuM5/nRqilZjQ2iz/iSlvkSpQ1y50TsBURYNpTBfWLFJDh
dDB9pQWvxuxRfMAKmahGU4Z96igm9rQPB8bmSRMBvKeFEAP/VV6lGOhYJmOdzWZtRozfda/ya6zi
am2nqJ24TOe2MPsFRUdIXafz9X/jDQbDV6qiHVEuJ2OLbK18ibHGM2j4Bll3qVX1XBlLo0VoB8q0
FoEUafyH04/QXsIJOOzUUWPcuVyx4s4cBZy1Uan6wzohKT/vJASr80tGcb5YkfePszMohBthS6Zn
Z43DMLM7ABDJDx/ydBkZoYrgp8L8/MLsGbpLY6yVDowJdr7UilcGrxj/AO+ai+pLHfXhWyTSO3Tv
xJp8UioxRtwP8swcuHjvpBq15lKSDQolzK0/0f7RnkIGfC0kMhL8E2uGijwoVGhHLJkxY4NF4zuT
OTZeECsWQGAr5f2Ine+8ZSWmvxt+tW38omCZOE2QBm8HtXZau2SUB/ITKqN68jBkFmPZx1KUSPzN
ty/JbWQ9YaU+l9V/qyRv8pv19IyTX6gfiYsBwW29iI257ZS8DNfSsL5KFShtvT9UnNbXluVswjjI
AcxzL1LSf0r7nAnsd/IdXse0xVAR8740QtzcmL3QLputNCGxJRb9SCpYvkqI53+J8Wruktz4IHHA
q+5faUzxO+V7+2HBmF4Y0CYP58SHEYM00G0rpl8PC5fJsqyWVTZrWj1CVkuby572qFjLB/bg3FrJ
HQuCBaDC5gNcXYpnKRv+cQMsrZKInlxlGZlhV2CFqFvj0MJjJdpp3HDQmGiW7Xs283mDzx9EBa/O
rtMom/3gm9NsSHfYbFKekRPVm2JIFhCS8iTAkLB7dPV/IeqWl7zKnSFlm708wpCqwYjKReuEaNVX
bX16OSxW4FVHWNIwhxI3FAn7jaSTDuCANhbIerBzJMbMBzbA16QDqmJcU3ovIbTCicU2PvJugnKG
3jkB1RGQ2cX95OfnrlT5f05o9G0nEaRmiBgkJgxdmCj+02SLSK7HrEJI4UVtJTko7laffx3k+BKu
DsdAvzvkz+IYHreAtERLbkFaPTu6AkXoachFKFDSlzWvWBr+zzonJcBLJjvMd4MsV+XTDndkWR/n
PdJriVtHgfSADSDpRPYEn5baRwQJLyNPvNTBiHoSOw4qsSF+8cgrxCuhGjHBe64WyMEQRzyJ+a25
9FM6n7utnvZtsEKVwTJ0+1aXk/5Exq76PRmqKh7pUo2lBwtZLWPJH385VYUz4T5UJ8IQPLHG7p30
otWVjNJkt9pg8Htx5BMbrjRHf3tuF0YW0d5aIGQYd2Z+hBS9mHemgaDIvZOh/+pwUA/O9eqZCiGP
KqW7UN+BSEG101YwOKt0dayFmxb921Da7anuQCrCpmNJ5Az2kQHk1GWNyWqwigx0SUyHtC+Fn9FN
fxdT4FH6z8Epx+o+p00o2l+Rlc058cMplac+lt7WpzfMjnP2/oVbBb6yvpAMUWU3RtTYWl1vjKof
jptKF3O6E0dIcyNlMuRlnqnhuz8f75gDktDdUAd/B1M8r5uw0EJucu2GXETAmQhkkp/GyIt63U5E
OjTzCQzuGnfihh97tDiAQ5XJJa2NFBtdGpmj5ZmzUBeDxui6OlEegTFnH3UC39X4JQiN6kFTFyKe
QN5K07vdPjnFgECkjN2n11WE8GMhYgV72eRm44tiz5y4lzrpUm33AkZOhYBwzRVfgnOlphvszMUY
GVXBNvrIr2e+pfGzCgDHY01GUkoUjMzCJEHCyxoDM1MS+UDmVGBGxkHvZ4XoZW+S8N5Aga2YuaR6
CPOrybcwz/VZ5WX7v4DtSU6MF92Edz1iVtEhfZh1XOOUqGoeRxgpGVQsF5y9iDtx3p8880kCwY31
NhSmQB4gDy7ijsMLe289PNloh+g8zeXrckmdCVRC0xeWM70CnluTLcZjVtGRD8ovLxONzM+R7do4
ETSG+1G4kWkTyNPptM2xmqxI6ubYnEIcM6PaR6pvuvqkpn0aqCEvr3JS0vmJk3rGbc7J01ui7gpV
aIytL5gWqiLLR/+RIEdKY9bkamNJrZEBNKMjvnwZ40/yvIUSaTU0PpufpnJOdREw3EADJjv3u34p
t/GxkTjZN0rcpmFjgtxTh8kThs+nH2bPJ4gJSq6OgwxdqJ7Z0RP6FHTcmJBHomrS/vtv1Fjt7vuG
T275HZXz94ruoBEFNd56oSNMfQgcLHd53cDzSxbGyBfS7v7h0U5qEmIJxec+jBckbxmPUmmWbv3g
XS8uArUkCOVPxLpPT3u+aFG7cBfIWchn/OgnEmysTzNNWPD49S+5GYWiS7E2qaWfT60bRQ4oD3Wi
F/A3dj+JuRRe9DP7ivVW9zMQod00eL1CfPt8blI4xN21TJKSfy74cOXLa3LcnqfV3P4/0JXLXpVE
KSb2wswE84sbvlKjCZouiVWEXGfebrDVguyNg7vT7e1XukUoRfE6rrd9RyG0KHo3V06mIZrPQq8q
knZgQ0kBm+5/6bcZwcS4R5cphxciIQ4JYzohSXs52Z0ZVaq3mVgSdelM3LvfSmUMKDES57fyKCnb
scJ62RriwxeWt+b9HSYr9WU7Eae6c3lAd2kYpyDrusdsFGH69EZVAdcnGnoxLb/8D0BHTaDKsvwx
AGlfxsyq9AW5fjqbC5Ku5zWzoxyRzMbfz3BtXDkqa52U0sGnBlVoumZ/Qr7DPxSJ7npamvDGIPol
Lor+rbvlkb5Xqa4LAIuCiFkaD4EZcTuoquAtF2SbV3vNku5Br9z0m0kNujiJeT5AIg2BQV83T3SI
fESWo8G3or4sKl8t91pOq5G/suxOo8LkZKYITyxNqcKpeLN1RE9eECAC1x4SYGLeba1N6kh3VXSx
ZWUdxj1NMI+BNcaBT2Cr5UeYHFccsvArU5H47qig4BPI8mPQwtw8cJm30/hxz2oS0onzEsBE8msu
fPFjZ6aNLgAlcGJ4hRsMZj6h+TTsF90haVckue+afWCCkamHqYVh+9jCG73/4eh/MeQvT1gjrU/M
TRFBfyXz/s4xt7+JJNcpP8RnvOvUSI2IIadVtlwTQlHJL117g2t0hXTZfjP0H3I99h5kr7YZTMa3
+XGyC84Qgjh/X6oYw0e4NzWd/8eObQgPfPDoTjy3fQN56hETkikUW+FWAy8EVT4nYlxOgLWM3sB7
6i+csTljpAotOhuPmGP9YKuS+2Q/kS/NM6oTsQLCAxl4WsseufWmZNorw4AvDSw5g7Rs4KKTRMuA
vaB0N3kHBGtBqsGdpb703386i9HGe9SKv+bnqTpdBKkj9WqLw3jIjdClgokRj1+lTK3PkUWp8oV2
K99BO58jwcPf0WcRZ/RjdCxg1ottolFlFEO8vtwdlDVZTS7+fqOlr6bderbN1FpD0fVGkUh6JMAx
MpFmrdsEm7qr0cTLDg+ev3O3Iu/tlesQVTQurDTOQGlT+ItTaLw+YT0nvpBfvfbvlD8fQ+SzJm8J
IwQymbRcONanYhh22kQqEQDuXMv3ul+LUWQ590sixnBgAlKjx2agqdKpKhx/a8moEFPhUrJdmlj9
C/y4yhKpH3lkLIVZQlh18WzSCgHDtI7OWbD+Xu0ZgefsO5WAqa5GH88TEySkoYgeDvRD7c1QHYyT
NH5HBT+nelLVCDgBrebof4Jw4wFb1jP3jF6iXVnehZZBcJITpdhbPphiHP5IJBzYjf0TKzBSDMxQ
Fdut+i5DxcbkeC/iTTkZHNLJ/nLdSpNijouLVK1erSRgUylVVSvWI4IrFrPIy6xuVV3v803RXU29
4KABxcKQ61vWKZXg0h1P1/cVsMlJwI77epayqi84fXOLZVYPk1lcuU5H2DKr5XpOL2t5S2Luzpqc
x/PhqmWgCLwz+iYsmcfAKhPT1VM+ZXjvWMhh05vfFg78j2d1BT1+HYIFCnvh6Bl6yVGSmSHS78zO
rZaxCA75JhuTqVENANMx4Mq4KCwkbkQSBpjKsT+xTU8Vam7VIwE1woiN0zsdZDKpJp7GYCdv3jbi
O3MLyCk+l1y9LEpxEOl34BlPG+EzNRsA73yOMXcH2DXsgP6tR0BXIpORnhutshQWn5Y/T/bgMC//
MER4Q003Kn2BGr0lAQI1MShdILHwxWbA93v9Sw1Xlq3rjD2niSk+6rg73x/fPkNCKLvlf/r+0yKi
6byQHwWMwVBzx7VaETc++vch3YWk4A3AA9RvTzJ6YVc8dfidEvmW30P4B5xguw0PZymqy1Hj0GZr
KxTAeiHISYxqX/7QIsvRnZpyl7rbbRTVbJJEk6YBsAPZ5pkwLtcyCf2BnuaV7qzXFUsQSf6Iz4gH
nKMSUDr6o3AbWzRMMZyWorUurtu/WG8z486/FmnBD7qR2XBxbmE+YYAvTATDo1gylmijKnqNZXOD
ehxn7W9YcfqNYq6dWL6XW1KkAb6Pv/BWwqnFNP4Y3xNujB4RkFF4lGjhaJ5/J2YMBxzTLaO9WYcC
YCG7AZeBl+n4C4vDbFpgK8kFa+wCwHq3a7wJ7VRKkeFS3X3G0PQ1EvOpd21JPGL5X3OyOpLQspBR
t+1E0eGrHc6hXiQ8/w5RktPZPJg9JY+ZxBGM385lkkgpumVqDuznZmmAyGn4kNxXwZZ/+NvyIejx
K7LpxnCfWn/ebrrDGP89Nv8ef1gX7SQ+LbJRUnimK0InsZUlQ+lFLE7GKSiSd7FNafb1AFu97ceO
3WV4k8Fev2YUBPqdYQyesQPih7lJd7xZc+wx4i6AbzYhE4l9YveGo/Q4Vh+/TTgJTvNdioXD3KdY
B13vrFRo7uKv/EfkGn1c/PMqCqFmY+HVK0ODcRIs77LyMUJXfIrrIS4Xx3G2kwgO9D22Yg8w64AP
n+2uecEah3qzv+9OQ05kjtJ9JHnHUBbv8ANIoKWQXGhaLJYFSLzMtflpqLv6OzELG7HkKsDvvZvQ
CDWNif/Zx6vguEXLXMSbPZRXbvDthais1zuzAlK6VH3OtV8qPX03tQ56KA7Tw/BaBvNPp5921Lr2
QaLpVdNh39Mqo5TuikkRNtFaJ3RtoQvFcwkCBHDOTyA4XaxvAHT+ceEnHwwjs5CQM52N2zU+uTPw
sXbASju7EF9rXyjrFikOJdq72F+eZ/LojJ/um3n0y3r8l/nExwY8wJGJUFMN/k5g6R6iidLTPcua
zYElNFr7Ux/zuosgMpzq7imGlTjnZVZgwrDkmyhOuSW8TwUI/RP+qlx6VH4UbYx0EHJYrQ/Ma08D
0nGMHJNtvD+G8kp88Wz2wIo7jYUtOPFs229fOi2t+05vbSwmTm6jOVqBY3C8Lq6Dlqas4c0vjamh
nhdsdJYUenr9bt8IMNyR9Gvh42PxHhIFDN7Rbw11udZpaj16B6HAnhn7nNLl+zhFYJDfLZQlezSY
Am7TzzIhUe0KXPfSIVhcvSYgD82NR/R9GK6rD26tNbGxW75HwcMaLjtuO/YwYf3vxWq46wuz8rkU
H3P3aZmiU3dLePlQXdy0MEjEn9ML2VUniwKsl8gqFN3vvAfZ+bYAUx0JNSWfBS6NlDTBICx1b2qs
/8dxMkS6YUpsy928RTde5SUOlz73yF/UwZLbe3VDHeVIMMEf6D1X35AIejASjvMEJMtBgfaVm55T
oWR3C6R51BMFDEY4R51lHLcunsImC8+JKwdNYdyB9sObTgVQ06CCfrXD93aHgO4Le0/d54glLCdp
oz6g+/uq3yUvPvlJTHdfegmFHZJeE9uk3G+soB6iREBiq52jarKEVWfxKuB0Ld3gZsU/2BQgXxYB
UdHOR7SYuU6ZbMJmnazLaDOVP9l/Fyiqp0mmf9brKHXSTDmDqvmtgSf/uffWi2zRj4VNZqMhGOPb
DUzLEBwNXh+UaKL7EQNnpPfbkV4Z3FjUlqdq0q/YtyEVFq8RoQN9rMlTewdKF2L9xPSm7ZbZ1xqN
R4EV48e6ViHbB+Q/PJgcmqzf1ixRi1l5R2EbNT8xgtJBw/Bb45clIk99/GVP9g5M2ZO9EhGyDF7Q
ozhCL3SoIF4bn9jmuZuRYQOoIWfYmdIMsaZx+r1IlvV4QZAVnfDzO/AOFbjWO7e98VAOEnuDb4MN
AEHmR846c3ifH5rFBnfynDNV97OkRVkA0kp9SVTocZgJ6aY53c+hVtIsmk3p3oT4GfvK0thyjtvg
T4QW3RqNl15dT214eFxxPlhZUWQcHAobfZQDIp8C6xTrkHYcvYJZHd8B/UWYe4wVBsNgrPl6UzFw
DAxudb/ZJSrvlq6+YtZqD0xQAzwcjJe5YeSL3AfmOVvv1dXGoTh5AMcXxx7Qv5kotNQ1N3g2HcVR
u73V+u2kC2FOAAVtcLDnvKdm2+vZtTF8EZZzfhByccVwM0iHtdAaKsnuo68eAor742J5Ozt4ZUmK
wKPxaIsWq99RHBd9R7x9Eax5l3+EBrTNMULiJVgsS0rjaCOytSa54L2VlTTr64VSuS4lINjQaBni
emi4anE0IYqCwaRMdRSK53kDp6MTwLPr5O9I8dMQYx1xnjvVqSshMeJ2ku7iSWhwueK4gBmHfGaL
rZDMmPye59nTOLyWlwPGeIrINNC9KV8+S+VERdzzGuHDaEI6i5rzwVWmJ3FK0RGfC7nuV/qs9cEZ
vaZxxxrXYRu90+cGcTwfOR1EbfpTbtTLwgsgLmJ4YQbRbnrvWzdefQud4XXp4Hc1njkMJUc0HBvI
kB0cg2rufQDuUWnz9Nxr5jUz5s3VBrr9uF2AbXVruVXS/cEd9mLcA6e2+uW4r+21eRmEuc/gyCr1
crthpDrZvJdkGIWQDcqjc40AG6IQ33OEJg/DgALmFvGTyfSGN7K66Fen72B7ntFnK7tT9f/Z25Oa
/ofeT4Z4weOtLuxx+vClE0tPSOfPr2yV4OH1HY8jvkDYLnoa64c/iVON4/AoAwYhSq/WRNJm0DUd
F+UBRZHhPl8aD7zAGJaMIkP/04Qax1WcKStZ2IWQk56lu8eLC2hCO81pEvGdt6h9hxwYGyOIf4J9
X4X0f6b4BlkbWptcqAGTSNqLkHT6c6Nl4fy9FaZ5juA1/4p020jn4GxbksNVp4IqEwRTOMmQx2J+
9SQ6lxBy4N7bDqAwiXHKMgHPG2OZp3Ez9YcWxOiA4wywnw51oQ0q1wFI2b8T7wzIcvz/xqO0p1Qu
8rgshZelpIdbS0L4jiw3FWEbevUACSmSKWO1TVyqnOXQhvdW1jgZU/ipSGzb0qqNmriBlNWjhaUG
KF+en25ft/Mwipl0LtzN3mFrHZ8Y2Iwz5uxMUXK/rdwYfrZP1unJBfVc9giIpguppaQF/Yp1ApXc
2Jb161nJkCgKENlfEFerusmAq6mzulo310v37duS0j6Bms9pUr/qRhgflUlG9rfSH7Q6FmYyVKRW
sw/ySrljoD1+jkRxwGb7+OOCQY55d0OWPEoCwGnrNE6X9y9arpbrqKlHfwmzmuG1+WW9Nmerl4/1
rp1ZvJ1Fep8D4u57UNwB73jDrSRxYy37AQwiUv8+J6Y2DQoWqx12mXscoif/C+JNem7RKMsBBAQR
mPVNdKB2IWx5o4niSlM31E8j31wRbgcPRsZyc/u7FBzA0WVM30FIEEssPW2MZ9hspmiFCjWLzI9s
h0t9kGuGI+wLk+Sjf665UIZRK6mknZUvgU3fzWT1NkptSpnAZ0UEYEAQH5uKjPa+6yGgXXHpwjT1
ytK+DYYK1F4M8J7mw67LrwVyiNvD+Y+xmRS5UOqW2RC9UiVwBNB2S73RV4RoQJ3U/J3PhAWa8BBl
0pk/IkkpzU8d0WSuo4nGOliVc79jAx0yKds5gt9KdVX89DUMwjq/7UNCE0DLXFXVlfnHAXg6m773
VO/nZngIGZ0jsIIxHBXc9Aq5wQMa9FFYPUFFjKxxhXi3LXsuw+DJqDmqHiozLAVwwEC21NxU9qGl
27tvU5RzbGqCaUomjeRPzL+aS+x0rSvJjFA9GvItkZsHPwFuMju8sBIO0nLrf/yYfCM1xocA+L8e
B6qT85wEE7hJetOxCnIywL4ygWrwzg1JxDXPYEybHpACZMrxPRcC6GT0fWmLGR4+0/ojMapP9QYf
QgLQYRrb4IlvIZzcxDj/Pu79vZnvlM7eeW4WE58OdLmd7a6k9VbMBbhpRdj9LL+Pl/fvqJqzhE8d
N1A0re2G9r8RbES1d3e8Zuj/e7JeCu/L1JE8xrUOcoZGfcQygqPq9OCMxRimSigLux4xwJFVDyGO
wYf9m2ogWXEdNbPzobEdNKn+XWeZVq51LeELPSiPjhOptIpUMI+nYOtLMw6jP2OBcjQXTzONjZJf
mBji/51Hd0b5y4hhGGHi68uPktcILd/jhpF4FmI0qsjtbYTGgL/OWXI7sp8QNH14lD2JvRtxMbR7
rDn1wZOb8hvq0XVOh3KFMwTSLpkt5j7rQpXsAlELzZWCy+MjFHd7cm+XpfC952YN68V32zHvsvY7
tr5UosWsvpZZGXv4durhYMuPc3pmOcChLyPMPppaw5LUPxhKes5iyi+DL7FtSUvHqECoG5VN53f2
/8WFTu2Ejh9detzEKqn0rHQUU6sQjv/QprW7LE1oT+WU6IoGH9BeD9xiOZNuYomSpQYNkvMN8gyG
z8sx+vGiXgCr19pDluOW5SZSyteQuZEREsPU2fuvoDtpMej4at6f6V7WQqyD5/qSBRJdVUEKV3HK
kScYIxsVvAFfH47y/Il8+DVYil1roIovZo7LujFaqq76qQ7pYFCKcPgCiHH+NRfkRlZoKcd2ZfVj
ObutQmtAD1pxbrU9dV2Y0R+WralNC36ilnbjzgn52229XJ4Yz5S+HgouyYdwngoQi03UKy143ygm
4pcfgpWaXC6WuLn2jzYFDa7Nz+5IBUNoh00EmFMTY+i7PR7H99C1AIx3nb4DAY2s6muwvDbeEY/g
LTDPleU/tAQfErgwzOwgZmOobYnrUPUBqZJ0RdkEQknk3uH72Q57lJGfMq63f1fb3TMJoQ+/h7f6
fb4bf7as4T6QLMx3YgICTQ3dXj3BaB1ie3DBWgU+sYCndQushVOLIOb9LK64km3MREfon0GU5roc
3d81b1x0ojJZuejHzNSQ6gtdz8pZJrdqS8prhi91k3xmq7ePcZIE1JPY5w7vog/VScCEOs+Ugiwz
K/PlpKgEMion+812ERl/aVTJ2IQ3hQPRSnaX42T3UjOZL65eS34s5Ohl6nD80YTf0EawPN6JUbjm
UyKndIL2WvHNSrrqgIg77ubgzf1yA6g5WF6oApCQTd2SUz7zTV3L0poGd9f2G04vtFWJOdbA0OWw
uvOkvVOKtNZ7n/Iifz4ebBBK9XBEWeufHamoKS9EJkNbxl66EDXewwbp72NW1Ce82k0Rw5ZdeLS9
BnLVMH0RvOgpcRsYk2PCVAW3OzPhKVYrcUdBszGiMC8AbWKwKQpEA2I7pasyHd6oIAdgHyoY6yQy
SfP4efoXVPmJR9smO5g+9o8cVklBahn+ps8QgFXRjVfIJZvs1arJ5PbA5GblLSL4c6h0BROMRDDK
zksL1apnvaid8JubTfYRgcsFysZkHCPpk1kuhTm+1y9tkhXKVhuTs85e8ha8o5fKMDggl95acWKX
lMiRrFrZfv+o0zX09YigEXX4cxGavw0x4Gp1fMFvboVN/TPdb1mmnvwZascmMf/2SRVWwvREuoZg
wc7adIiWZ8Tasf2osqAWCbBYV88pyt1f/9VW6N9z0evul1d4iwUcuPn/cyVNMAMmfsiihmn5dZUm
IVi4mxK3dY6CWaxX0Kra+dvnPHPJgAgKrTvw4fXbaCeXnrQ8vnG5p6v6D3mloMWT+7wXE44m53wB
vMvgRCG4oWfnxGtS6nPNHkN4xZ18f8DrTw6SmfrkmH6g15cIz7ZE9p5G8Buj+mm0X2I9VVELAbfc
FarWW+UvqhQYtqapaJyDagMf7xTHKBAxcyxXK3EgqWPytv57utQDwv4NoN1xGt7qFOBxRU8cJzu+
NCuDJ+dehd6/8y8YyRdRozUcQKhZzMVU/DP5eZ1PS2quR+7tvPu7glJKEsCQvedEkEGWNPI/p23z
XVWhg0mMt68QXBMYj9K2aDGjNafbxe+VFUCRprv03wO4CeJHc+YpXLrGa8qNprqnlsvkEfxYNfn/
odT7cGMwqlSmV/WM69ZcxqmGh0G4tyk+xjkm5IjzsM5VAHwsq+pIJNdYWuLG4skRUEA6pSwizlJc
WnNxw/uAOCUGi3+/27ua0nE8Xi6cwpBCvOSHLzrz4zgN3St/M0czK5ZQJ3Z1ubsZjq5myC3R066S
uQ/rqda/q/RuhpK8g80pYe6xF/KXM7VEp7WslcxpMSGj9kJmfUpFPXbZF1RjQr/FBnHj1DFBLyuR
vWhi2/flCJLE2b+3nL2xEoY9WNK31YDa7hLXVrTqGUeF4bEVigqFvrDZhTkrxKNOqBdXn4eTPTUv
RIhLNUWuWLJSVEGcT1LTkxn04vnza1ACXHr9SwuPLb66VuSN4KHBngZ2zl+5sERNAnNBtaWBK0Tx
Ua/Yd96PFrcPdxqzUVnfq8STLKhwVc7JKy8IdACLgxXDYE98R5cgKuCX1GY+4KoeuH8Znjz107l5
zAZdBw88LYkY9xwG21KhPsscLSoIjSbwsSI+lkQtRe9DRPKIxH1xI0DmiaiS2JqvEL9BdeuwbdEZ
UgbSr6gpFlRCjUZq1Nj/1ZB8Hs6P8xmst0DQDux1DNG++olVDenJux0wo083tZh5H3iU/tjwqqJJ
11RMN8wcm7ns20uvJ9gIRjKvjO99gnIoo1IpOAcOcCd6lor9Oxln12B91rlfNzTVj2mS0BAr1l8k
sdGqGNOxuZhB0tv7dntGD684EOiuDwPuOqaH1u5zxhppRuTOBnoRYQJSsE2haIhSvODK8oc15N4v
Am/uVdu/Nx4QH+hE2PAMp1g5lhPZXzC4fA2+5vQysmRiSKlVGaOm93bgzAmrnUsWP+AQdzm6K8RF
gMUNGkx2ICbTSoLh70KrYvRJgz3joEdOLoFExyp33Zht5SFQvrAR9m34KzxMhBbMv6M6L6rxWV8O
l/LtJIy/4K+6+bJfg8qPgqe64k3UcudUneGHfSY6vHKfvWGGa7ipjThy7mNytQkrCIlTFnRQxq7t
Vv1AowEeU0DZfcX9TCZAF2IVfCy76DBvUV5uvapUbNVoDyf9BtVLI/diGnWgSg5TLXJhfw4Ud+fG
EGNda4aCBuYdK0ftn6iZwoywh8MfZbpIrIJV3XpHPnxLBUPVvWTpciDljjGAGRqfskqvRotwQabg
TI9X5qOywEPDCo68EiKMyX7nw3ZcNmtju3lbZaJ1HOCCCIRq7LTp3lYqcCS4eYV/FShRJhue7jdU
EwERC7Z4YeFiFKWFwS1uAuBdN4Pqst/Joe4t5oc4lVKkDw8xubFPwqfk++M8uOK+RvtbSCNJAnez
HGZJBxGCqFLjuSMQLbBlJsapAnLSdPK81djZjCrUijYa4dnkEsydsUAqHiazvYaDRacNe9Huophu
J05mgNN7TLU7uczvJyHkxRgZxTuEfRSV+o82KSs4c+mhp0ZZ73WC2TNOyebBW9dZO6sMuKEu55th
O91BOb2RKOAhZaoA+JgG1t48hPeRiqsM0LmxH5bMxwRy0zubmYjdvbe8JDWB0LcudAg8cECLGh5x
fKd6RhRpfWjOacrtdcGCoaIn2a8pdtvmlAKRzzoMeXBsx3RXpVlBwebgSyPd1/HLhlNjBsBNCohE
9o86DBNYk6ixcXGT8mfoGMhvMA/Ke6U52PE3zHynO5jPvlIg1zlv7QHqpWK//wy8qAtr8+PuZgSY
uNApiL2nblfA+Mg9+72XzP2gjt4KJj50rD6aI7dpgOa20IFCSU7VF8lcHUyvqw6TCuPDfk6I/jpT
tGn6MiSLvSvuIJ2cnjS3nOtW1mhH1quKLlv8vQcGW6EUY1w23q/KF0M8axYJu663GcMtNvd9Xber
RhrFLZlhYXFwnEXk9YIydvcC61H8nJpCHXrhUjEUx99Rw5YEXS9QZ4psNmYrno0MkS5tHiqVSuSH
IAGdhXC3oRU6IFmNAURR4AVbx0vNpVBTnIHN/KQv1IWunHNh/YEk4EIDuvUYqPqsSDxMI2LTRQaq
o0b+x9EITMhml1q8JWxOstIqtFSSRFPk424yA5Mi/2HXG0tjQKytFi0eNDEGIIePH2hnZO+DX4Ml
QpRSzZURnNh2sOvllKf9sWXqaONjVncmpMTrHLDMOWzvqaqQ5jWrhLHbUo5jAjg2pxwUhoMmu+P/
9p7Kwm4D03X66IIfrG12i0U5iahGFdJ3/EQt8h2C5mBPAwUDscD5kuPwxilwxSgd6j1NOf+Px9y7
z91GjiooFthj8gFPEue0hALeO3BeZwyfRUhyZKtzVVMO/2n1PZJXqFS9McJu6bamdKi5XFrJOQhf
36ce2WT6oOTDAt/zIz4pZwgiiuh3ZgEwnCRouGNfYtijJez+hjHoqgDOHs0UYey5fuewP0gJUdYm
4GW/KQZQaXOB8Ba+WdgrHDPEqwg4ntTEyOl+SLR6fJsvAXHChaac2d+Fb3uZ62MqvrvPkjy2ldyo
QItQupb38soWg/LCpMGd5DmujHmtXUXU963YQiQ97xLSdw8+jZB9f6AExkjy5l/iB00RcYyINU24
C1L96g1yvN6FbGkuJwF/D16RnZOjgErw2gyBCDLdiTZkHFu3PYEYiLKQD2BcJ0lQ/vAKAf08jDBB
PpKzlbJVprPWp8tiri96JB9Hx/qTx67lWlDKF6c55dLcuEayF3IDt9u/hfWB00h7JgiG6JymG07q
cDAy19TocQSyfwt+HL49HeNMscN8XlvWPOkdv3iAz+THkAUwe+/DkaCk1vAHwRUqhj0fjrKPZvTF
MMsMh28VTuJ7z8UJL8ni5U7LqFNChWqLzAVZo3kk/YAzxqJhoAYi9gqkHrFuhtuwR/S42LLH/ja0
rPrXCSsNABOwF57Sxvg0ttmrZmI6iZEVze8vmJVEjQfhdBRpgOtrL1c6R6xiLEM616ivPL6UL699
T4G4ZpFu94jbUxAeK2p6Jgw/2FQXzg/QU5wFhNjrQjKE19nokOp6Fb0z6nZr4MKhCNQvnDal7jaP
WwhsLU+puckiJDHR11Q2xABD+SPuhz9N4saqEac+WkXlUv0uVATadhYqotvxpjCImzjM/Yq2qyIT
z9RuSsEg8ItpH7XCt/V/feH1sfGPK69qPTGvbN1T4GcSlzj5hzeDrZuu4T5FFd5aM+MsZtq1mgHX
kzKGWhXDI3SlBJlQIzqX6Ac8K/K98l3ZW5rdxzk6hZG0gPjHcQUB68W3qypdk24D67M0Tkphdm3Z
8QGWHV9dDYrv51Np0oax/TCtu4yUsTjNDwJm3AUW7twaFqfGfuLTYqEM02OIJ8jlFQfZI+1UBLRS
8umvRn39NyT8kDwleDxDBjZrn2PL21sALq+f4jxuZFXeCmCj6zln0ykdDkidq313TdU0srtbRQPs
Ka/cstPx5To6i5nXtc7+7+f965Q/oh7W6ZJnWZoeU3auuRH/rzHYpT9S8cK9cjKhEX1RBNj4vXuV
sram5CURfRr6/UWwqQ1jaSFoX1zu7F+l2fYyRre5noa8hC8JP98JejH159j1MiHNVO9IsiBERLTe
leIMGE4DF4paYNXa6/JQmnmJAhkNoec613yMf3zce1t2mnNpZHH1LiQBiwJxo8KXaOGBnPCuL4up
k3RHNiwfc0WF0G5xhLJIRYwexF4tk446fkJPfet2PD02gGq1Fxpgz/MJcXmH3hrEGvExIi04j58z
1ESHDsf2X0gi0gRDUrM/24YAaGinBiWoi0z49qQi32AZ+e6WWMDuuN8ijgUcH7KGGSqrJPgAGhDG
0y23DxXFsb1UMyiuT34x6EBu8rgj1MVxIaXlrOpbV3xrBQC4gVRYjgK36pE0EjexiSlN9OrKM2op
pYOCYXYrClRxmkr9NFJCXOvq+jAQ2ma+S5B5DV8mBQV6H7K5d6vffbHT6ebQ7ptr+WKmWlb+Rp8v
HepbAomAQ2+frTpmejIe1M/jaBYbm/WKDBEgmrNyqZpYAkEh4LRZjCsFb16OjCJjP2t1zAIBb20u
6PFNDfh4bDlovD0lAFzPUmN9j4ADQMYG2WStwk3JnYtlUEIl/tHzNDS/gZ9KhK/AprmCBAlNv/wd
rVNqxnMIwo3ZjpFZZzBudJKQxGagBpU8HxkD1NjudLoi/8AB6CFmL5VV4GPrX2MfyUEoe3bB/1hu
hsu3+Dx01ROV+KR6o/mTOxpTmMBND0nEbW0VZloPk0TSTd9/UvmfnK2bQlgEr1QvuRBgVy5BqNC+
YMwermmbIx+YmhyLhdIuU40Z0LB5t2CtnAhni5W6EXRTULILgey8EXhOv6d4hs+BujyupSwnaNF2
dJNFKvOrfmTymv1UPtjABzpeTsvFjNJErPcRWfjEPnP15MO65hrOr6wr4HjhABqry5oYpD21+pNj
2VGdpqtRmKXt3DIB1ERCkRHR3+WyTMtKNV5yv07562PRVm+R2ChA3JqYi0FPTxLeOd/TSYZelMKb
CxnEsEz4WJHxp5bMqqDA7APkg2GalRLhaoku3gCumMTnu5MmK0HtPE88zAVmmNLq19UzMPyl7QaO
ICJquznylt/rjdmCVFmshRsGhJthkFd+Ay5a85EEsKigM4eJW/4rcfM53r1X4r5aedSMAbtn+L+M
SHP6Zukv3T0U0oHl0nx9cXxrsucvN1T16+/aXa4gl3zZyawLaygP3qJ4luSf7nZxRffHyyJNRwFv
uD4ojjYP4mYswwyX6QBeffK91N36E8D3chzjwFpj01+YHxmhEWiXI+8xnIP5Zeq7O70xA/uk7Sci
wnwT2/vcGQZj/KE5B+o7WO745JlEVJRHuRHobYI5AxAXLGxBS56Kyce/ZbeNGCaw5x3UFGwOg5+w
mMxTcC5TvFYXG+ZZ8gys5XQkfce7ci61yZJw9tjDdadE4KDHPLN7VPHxNZPR0vA2GQEBQ+LjlBmS
j+p5oYlOWvJo3BD+ohwslzRgVoi2gexHn9IDPFnSidt2hFKNrJaP3EvZ+4NW9iqYE3ON3/VRrbAz
T3wLAyHMuysvFkefILh2565zpOhi8266T5rE1oB72rb8s/fo/V9FHR7Vz/i67Cjtb2koLYalknDw
wMW+z3RgLMWLqZc/QCMfFsI/jVP9J7VNpOdNg5GOcHUMQGsqsbymy3pB/38OIR6cDUdLD9FRM+QQ
NGgehi7agZAiqK2VH5oiIV+QxvIE8VkWigoLZ3dJuQL/lKDNGdW+GIBCzNX13AkoBUf7kSAj9/Yn
dZzyQ8XmJ5jDjgsFGvo87K1GYGkpYTbBfcTDf2r/iLMFxYb4cCgWno01IZDPsxFt4zGo/NHUNraC
hBXgxXT61/IUErnI/9QcXwDIz367Af+AIH/paOarT9ZZ9CGyXzgr8pMW43UzOjK6f0LNqH+L8B3U
3igtU47v2WgHc/ztEhhX8AB2EVf/Bou7eOrWMyu2kh/Rgzi0uvzMNHTiXIkgF4ZeddKrJge2LpCC
W5LEqK3BiPaw+nDx+t/Y1BmbJFvSPYJQ9hVl2hMUtVukqMUZ0d2wqMPakB4CH1u8OOsUKhJEDhgg
NL3GMuE2qK+3K56CveFHz7NMNW0kxsyWhSVdJymF+7v3knZbIKQ/dNtQQ8H7JBV1TtSL6oM9WIb8
yOADXTRz+UW+LD5xjkBvqzF8eiyFhR35W3iF7tZTw5843FoZcSubOBJoWhWUNxeZqXhslbFC+us7
5iggthogsBFSzDQ6b/RhZVRVQjUy0VsU5lRnMcawH4Wy39z4ovcIUZIuedTqyLRE5pQwLwD8fa/p
abt3IY+ufAOozpZf/wJNgQj4c4sId6FxJMjL++UeAZiOXKQu65FNEQw5NyeFCp/2tvyPRd9+mbUw
hCyIdALa0xkjMhPddv//GUlXbWr9Is7Ynn+zUvTTtTkGRBs4HIbQmcRpIWm/AJcEt953xhy35cVz
vJcC/05fwHVtWB8XDH+ooZI+Ibn9RPh4QGKbKpL2jy4LhBaL6kbxLbRywqCsriDCz1DYhAxsDeHR
Ua6h8iCD0e3MBfzz1m/o+aYDMP1ZIz/gywPa5SsN48JZIQGZmzwchUufLMZ6GJfZQllt/fYSNq+k
2mmjTL/CxFnv++FKPXkOSwdvqMw8VXUcza1d4jQNymRHp+Gy2hrXXz6xp0o7C0CYiS+SjeAsakAd
A/B/t+gWWs2e0SAz+KU6oXJDK25gslugQPdUQBzDl/btRSMJQHaMztGlxnvbm44qKIzTtGy0zQyD
vpYmKe2rivHDBhVkbWVqW9+tJnb1e9nbIQVO0n+p3Qjtvhau4MdE3rP+jxiee6N216bc1iyeBf2g
jMpR2QHp2RnMgYBxt3d0P2WF1DfLmu41PlZWtjqx7Ri5EXMm8Yv/EdUmO9wxZmnMqOf0rg7rHWbK
xvWnDW0lbkq4YgG5XQnotUTa+zrrZs4Vl8rh2PxSmHhnOEud7ohsxg4Flc7SiNqvh53P4Mu9c5ns
5Fh4ONgMKzVK8TP8YoMbyIjhnAeBQ/stTHhY69c/3vrqv9Hxthytogi94Kfz7HwQXDfCatF20t/X
IeMj//Hw/abAiG6npmTRa5SLrAecE7uvs+NL9V+VI1jtXNm/e616ddDfUkpr0U6B5TaZktFi3Qzs
JhBG0Eip8XBixAPlLH+PE94B+IbE3LTyNo1ghCvmadE6lbGPndvdTZSx0f2GzSR3IoAohGb7qJ7d
erJMGxjMQQ/S+be3tRzkkkOaR0dHRA89LFby3R2+xrh3oj8mNpZlcnjBBIk2VsVbwO3ecKt1zVZK
yaQ6JarKVhxx9Ti1EqSGqLt/TcSBk0w5/ApI3k3h9Vg+U0nXlQ5IkIWaTun75/zqd3DjGaSAOP4e
AgAWk21SI0+eiFgh31bsIO7egiOaZoMR+NhWHc55h0C2me/Gj5LxupD41zHSOK6flKqQD2YcEwiR
dF5+guBMkVZOCqVRvxzXgWiyiQbOb/fREtBdzt59K9J5ZEN/C3fNFCbfisPkd993OeRvF930q1KZ
nUwVT5vff4+QopCp+1rBuB7RHldgL2xqaHuEyxyRsJJC0WuVEV+PoXbrkqzIEEgzWIuRFqEihFi/
6DTfFDw8Avtvytt70Qu2aDz2KuSRwNr8nj0bDApz7hEg7X+gJ2NQoVJtMECDFstrZEJ7vO0CiYWl
Oo3xJ3LcoUBbTML91va6c+/Jk0CbEFq7OAvhoOMiVuRPIpEEZpeJeQdBrugYZtMjR8Ae72kEGMHQ
yarq1I3/z/vg0TteAfSDTcMmqA2CwUNvOBzEW86bDU+zmkk42BLcbu7/3birSSv/hbwk1vMLUBXV
TFLcXUHzrzFmkBBfsel81CwtM9VMUdI3B/3+Oxq52edfMNmluAmdt7UwDjuhokjxjO+b5eRitaQa
xDKd6q0W0CnzclmcPrnLtDbF7ng0uvbYQWwFGfoiNSLBZ4FKFtKPRWfpC5uGwJW1MxpvlHMIG74g
IJ4SLdYl1dQX+EqSFPqRfMojaKxC6+/x0fd6JBZAbiDONhSIpxa3WFqcHp20eAZpo6Myp2k0p6AB
Vcv66m64zrQvc/0ARyTzaNJoTUg+4kVgLdgkFatHsZtcursytytLoXr4g7yW2t8mbSQbvOYxs98g
Dy5mi2UbH9loFNce3SFwyhhwotXSbRG6PnLgGybzztqdLVQ9uGXZy0p4NZVZpnhnbzxXi/QCxqQC
NzmST43L5oa6WK2fDHG6CP3HErZ8fuGlOpBiWhGyREqEbiUUY/C9thFQ2bcsYCEjBqfh1yX0ml1u
T/4p1UjQBiLDHF+gL/+D9KO/RW/KUu5GpAFNuzed2j8nX6xD0rFux/maexnnXp4h6nn/0wT8qu5/
hO16dj/aeuwztVfzQtwhFbGqwGSb+XK8C7TblZBviCAa3XhJJlxHlUt2YfrzpAT2qUp3n/2HlkEo
oKoj9TJb8fSqus8JkjwkC/FzZQle2WntYA2m1SLb+Td11QUxf0zi1JN2OiAnr9q6qVyjoEPkgeGN
k7CvDnTL5kCxKuXR62S2pR7mgRXbk9Z1FdC2GGD8qOz8BrZj7PPeckPHYZUSeROM5gLR65/rvs9K
YJDnLXk6E3V3hLQf/7Af8nB9cTYE8GerxTh/pHjEq4u7pxtK3SQzcXxVxRc33+ljqmuJMDipVBrK
Msa/eZzdxykDg2jUMjfRvpe5i/xkmttGKyru99sXgASSsP7NfaDes5WNx4f5jj78Wn8Dfavg9VxQ
PgnQACbpEu1yzDJ7SG4tsTe4z7zOixTcLmAqPagsF/TIYCv9TLQoBbMbgQ5UMADflgdn/2dIu1Jb
IB8xGgOmaurYRjMrJRIalMSx1gMEvG2TiHDavSf5vvInAf0lFcqKdLX/w/YjyALZGA4kqQBqdgxB
O4bxuKmu42SQf+qwP4PjjLVHKHKI0YPxoqJfEKgukzAkoH2SxfkQTkokLPFsSO+H811NolbUFNpR
MRJMT2wiANxA/ETQxt4aAg5PnYTw0R59E/qeN/WYGJ6/Ie4LOFzGivfhj6TAVssWlDT9644loiDP
1PmTHKqc2ZEY3x1ciceHb44aVzGN+gdmxaw9XZMt/Jq6/DRmV3qHo8cwxm1Zq7A3KGOwhoqDl7wF
eI7h1QMb4XPCE+arYMruDzHg2p7dywmsAFaEQ4Yu3LTqZ9Mtjm17H5hs0/Q9Tdyi4rQEwIIi/tT3
+5v9N0IikKA0e4+WgyJk/YpO8JC2QCB4kipAeDAkt5UusMpC2eDRVJKxyyZNpT2roIZTskLDJki+
z5Mm+NBNE80CbaXYK62R1mKa5lWOaETfahjBf6Sxu5CgZcqHRFmy0IqFKOHni06Wgt8KbZHbxl6U
T5h7gZRZRtUzHLzvJ3sDPAjk/9s+TEh0JGumRzPZihvKXzFeHxs5u2nba+nRBxIyan5PXvxC4w61
l9oO6GQwVn2/3BgIeqsuiZsIkO9+2x04KyrxSLGlAUaAgVx3y3Ka6nHqSwJWa2IaW+nrfs6j4xNq
p6KzxtlbWWCGdHe/duRW23JRCuy41R15avFeZKXCf2dvUct0ZX0v3pUujukLgzb7uMltoZoV58AH
wtDwKS3pu/xlr2NNSzsYKLRDxCmHjnd6XTw/30RcP2Bmw/EpH45kO3P/a4a0GoDRAZr8YMxEzGnt
ayKRMuRb0eHAgqajteRdEaWdWeX61a3s9PzUH1IyOqVdmcP87x3GykXwrsjnMgitB0Xl4LpVeXu7
HLK3tj3q9a26VlERuPv4q48udVaY9udm35TdynXfLk+NDES5PuIEU1MVraHVL5bgSxE9nhI1LASJ
WKfI90TqAYXRR8T9kp6IWmniYncfPg7peTTDlnc83zJyRSWAPRBvxznpeaxpX0VnvbG0DbSwp+ig
he9raS9tMZ/oUa1Ivtv5wC6JV8IWmARHTsLLfAX0b7KSIoMyzMFee/nE42UTAzOOOQ/VreBUkYua
DKXsAJSeqzcUEb81zDDpkdf8l6jfIlM/GEq4XDMhjKWsTZVjpdvynKlmR2txE1yNOMKNsr5Xe0IP
3g4fpmCpP6maoMEBp4tlWgDg7chH8vnFqNGk0PX/6rR0A1XelQqEhHP0wPO/0xDn9RYNp1JqVQix
iGthokBfsqiXiTYF9J6RxgSAEv2ykd4TNTqVosAvwV7VyYiL9bB2lOA6CXDQwop0qqmnAxCIqyQP
hfF83/4q2e44KZBmz5z3xCv+oUOD/C4e0a6U+76TGw9F+vOGFhxjn4z/0ikDIAN7Gqxh0gXc+no1
IU8v4q4RC3IJch/jAxgOCq+2rpMeDnOzh392hVmEGQv7pZmOVTMN3z3XnlQdJuvN5wR2cig2U2lY
uKO9yxKuFcUZ04UZN+NQEN3dbUNQGbEFywkzY2ZfxXBK57slJi6I/1C90enN2gyuVIIlIajMX6gG
sONT6oLxP5mMAfoNgApGcOtOGCqX214dYb0zV3BH404DYRui1Y2WCJa7DkEiRp34uhyoHr/a4E5q
V4GmNycm5ivqEgN3jotc7V/a+7KPbr5L8OoYtATR+9s+J5JZTmGyx912p8aLlXY28BA1uCFb3QwV
UMHWT5Vb70mt+THn1eaeIM5T6ce5kUx3N3uxt6wzh1rGaNSVQ8A9xyLjwz3VAbcyqoPgDHtv311q
hzJqP+56nMQXiUfFvx9LcUVHXBE0ZIfv6hZFrDYxFnscnyJeZpcgqvK7JUnME6P+Gzx5P67iOIj3
3kr8yMI/xnFPcdf10CdcC2fjDrctW4R0oBAqWEYevPC+atCqfAdCsQ33h/gjUhuBEOZeCHV7aXk4
T2Qkz/izqbnaJm67aniRyHSs8ByQRY0Dhkr21kWEgv2s8Wc7kIWAnwFvjP2VM0vp4hQ9gMEpPImP
I37o3tx3HnhNXMfL6Z7tyMvLWl/j0qw6uz64Cl0N2B+gSvOx4kdkUFa8auOfv2A/hk6L17PtQcHL
YlY/eqm6pnyADVTDQx6Lei37SJ+iVQ3XJWqJO9Pw5V49GoOBb0tIczSne4/djDB8Hi4X0a/OQx+b
S6/2qpeTwCvJKoCAQs/8P83wMcgmIUBpN3HakCyGtEfz0u/ozrQAUqfhI5RXlFBtbYrVTp5l56vX
tUdsLzSE6sieKwXjYSfWVgMpsJ8mmgfcQg0K7GWkq6DCQ0XY7dNXlOCCA4DSrySsoDRZzUOwndnC
fwL88Bm4hJt0McCCFpRdYC2iuWfWi44ztS6mAnais3ctUB3tIp3HxjBWA7BWGBn/W1g3qLa9xI4c
9dFpXFT6V9Ru7oNbtZlNNKlfoowJN8CDbzI0H9Vc3++3m25TTIthliCckprQT0iaBIWDaVp6ZUjH
rqNTrrtpTQuETgU2mKlK9hy3SnYf0aLUEe2oTkoym5vqduQ0hat0YJ7rz/bizg07LfouCmmNkLxz
GQK8uCbChJiUZIUpAVl+R0FkB5DxIEKA9BWNNOpc+afpLvqusOPP1WBU86BrSzf0mWVXCUk+alK9
i4c0wT+aMXSyIoHMOaFgFBhU2sWFXYSai3sxnGni8BnIDfZLdiJmBg9FPsibAYUzy5MSzN6Xg312
YeNuGFRq65MbjLGDQKUtOXKfP3XQrZYBGjlfBoa+SPHB8oVK/HDput7hV0Wxj9j/Mzt52+B9n634
TWSNzKkgtexMfpxqrQvWkIJwnPn8BSkXY5pLHxbrDQbKehPudPyCmkpicKGtObMkxb/Xn+FZGXW6
FXddD7bnzslxNBaY2WkBtYqb3v59WiHtaXBaZE47C85mH/Ogjauw1L9VuoLpxG9IYI8g1JS8HfWM
AnX+r4H6MI/dBipE+yEmqSoDhEBfNACOT1S99CEiKt5gMKiWD2m5YkSQKCbFRRjxig/KXIs0onq+
t5po1mvq2soxbBe2mMfIf70t8AiKUWfzAz8f1Ga7Lct6sOnNPrJ83ffyMGWVv4KyhweYwMqHO3vw
AQYvIG8oNxbATXkAK1J0skr4HNY0/MdIB1/vwAWniapKQHJJHNz5TwIqWQyTi4E1h/uKvfVk/OEV
T4nDP/y4zTDQAQR9RmvaS7Zo/x9GA8ox+9Qi4IWz+XqfPjWC5HuRX3TckrjrioArT5NqVJe8xUKS
BrmuALH3WvUqsCXEPzbaltI1MuqAobH3M+wILFsMtWTZHvqipljx/SCCDQa/n+2q4IImqehzj/Kl
uZGxbWjG5cI2ixB0QDIwh9os8uxOKBuG5ByPNOJTgm4ss9ZDqsstnf0Kbvnwgqj8HNSyRnz1/Mn4
3hwQVvO3N64BZRuoRTgq1SBv70rc2sURz8W6Bxq1yzu6AWtPSrPd7RGr8EHz/uVeABS2KBAr0Jl2
0U1RvC001XG1F0B14n+Krmx0YAy0Xusuo+GRFR71JnyUPw+kBsGLg3kWwqOoISZhgKOPXpA/WY0G
JlbEn2o3/IHdTu4FiaNpUOdiLPAmzN7Ou2SL6YJZhcIcpeaDS03bPD6jQ0exscbC+VHqGUw0on9g
iZx1qlu6S1vwtxc2GBCBk3TcXlRtzZia0J6bUiQk7Fk4YKftaQTzs5diL5F5CiwymJttL2n+//P8
8OfkiOuZ+lHuHJIo9S3YEoQHH0HRZ8ZHvWgHNzFYB/49mfgGAkYnOCQXQsxOFh0Zz27sYJeiLvWY
KAs8kpjpOZb647RDUMBTI5I+AIKFkuPHBcGvoeYcibTq9xsfLquig/EI6oCs5XhtBp+jJYJxc28h
Xyfd22z0GkiYKxrMCHrgRteLIKELbimgOmyg8d0kGq2bOJPxrsPN8c6V31OKz0OpPOk5lc+x9xyQ
ZO1cRfrpvfnp4RHWkjnTG83/izpdLdNR6eL4jeokKMAEUlNT9sTUN12rlYvfNBR02yZLJWOko8mn
QD1PrccSmNiGReQFwXOVoAhRRx+saIsAVi45T6/cHH6K7sjk1kCPr3+f2DfO0N/jXQJwSUA1hGHp
Wky0xd7f5+hTTT7UgH/owEOT25zwRTKKnpqmZHKciYq7C0upO7W9XbDbJ9OFaCN+TXUNRxTr2Zpa
0QQgbZTpTdkvGDq1W1fw0U79Ezc837R8YTtLOKiXcyuyJBK6+1rj1fBjKflQODAImyY9oskfPH87
kUC57MB9KWMyuds+3EX6RCphKAWnjj4b3Z87VBLKQjyCtF2/Z1ZD7TbSjwxc3Bhjlb/+ea61lyjn
PjtE3qmbiwkPo1RmsvqPmmgrlXzGYomfQV/DlRtci/op4TkR25qRh8CB7Dlcnjhmw+rWqR3j4dvR
ZMJ5d0I/WxHAipbMD0kjLzf5uxLp2NXcFb97ymQRdJVgl14VmPP4QGI/m8PrSOUmMsF5lXTPLZxf
qtJxTdbRYpszJ9GtzelFGex7nQ8vLpbmXzNmYVO1nca6uiyhTn77rhQ1D0uStDuAuvUx9PLlsFcH
bI4GGJR+G+asVTz0NBNDFijplGXgpY/zIGEuk3VJuNoGCsa/orBwa8OMkHtO6mLW+xUimQ7lrWyv
adHJaZxYAHV3/HRlQhZY8wlJJG/Wt6/kQ+BO4TXx+YqfQ+OetpOLMDYFxeQYdsBW4lXZBHs2kPMu
40HtYojc02xZ5LAtrfSHplydwt/8ZvjaXZkm2Jzzywvj5hbh2MH0hPoJ2wYba5A6jHqFgBt6ez4S
bGXBB+G296f+QaqDiQgqqEkIrfChTezw74svM/BY40HCYLCcdqTGk86HT/Hvlh137A1IEEA0FIjk
N5bpE+uQkmmv9G1sZoXuvaqrhExZpDDPUQYVCMRm9JZqFZ00gdBywVUCRvaQJf2kckcbNCafEIbb
3wzXlUJm4r/z+rbiWucIMx7OF910970nWxNtNpyGga1oQG0p/+AkZY6ZBsXM+xe+MzZcp7mLZpEk
UlbgNh308Ib4vbLW6Jvn8XSKM/hu4vnkY2XBEWUh1PIHzTwWDSEJ2J/Ww0HkIDMCz8uK1ciWjMvX
i1ydwEJ5UzLw7UXgg3aVKzaz1CpCXQvu0b/2BB7WzSD07y6dMNKanMU/rp3Z09IzSEOqJuw94fkt
ITox1jhTKfYb56f4nJSj4nH+ODra8W8y5Uiw4frHJsDE7CEmCa0TPng971Cafr5WENSakKJxXLk3
A8+6hYJJT3cnyKktFBt6CvodeleWxhYenWsBr3Zp9syw9MrxykGMC5/8MZCoaxZbsB9PzZ0XDM6+
UXNty3hhzHPvXxuuuTzkjJTQwGGYkkQqMAZqki/3Hf1dIAXPwqn57IoPuRDFl+s+bxlfcW+OV51x
GUOAOPHwxwmG09c2RlUSTE4iHX3BScguXYLjz6Bbr2dfF01Y8S7HIRkw2k7lKDDqEx7h0+s9trvi
FD9HlA3lpgMrVSpn3S7OWx4mCMh8EsDDW++0Eu59bdQwOWDc3S09EMPf44H2wpZAhJwS6ed28QH7
mkjn+fs4SzDxH88TTs542twjL8CQB0962LawCVD52E0qlaES4AnY39reSkWbohRGPgSxBSyjqB/L
CLHB4kNBAC5DFpXxVo8bW0u2AOSAWORm5t4KuXD4isL511If+Sme2HbbyNfBsIt/jTuoff6LYLpT
pdK83rqu9DFG6OMerk/XKRaHWRcFNuUUJAys5jdcdVTGnOpN727CyGkfWbo3g7tU1D3odhDH1jGN
SzY9umqW7Zl7NhbyZWQDOebzLlLB3xuh6zt90DAbxWpMfvCMMhoXmDnYEvzoYOF+/iXehksS1AmY
o3SVlftTR9dt00lBFGHeS9lxU8wHtZdlGJ4qpWP2Q3Cfni/kb8aJyTRrJQJOaX8FcEL5MioOr7Rj
kVHc0H3tqLDEE+pfPRa+TMLZ+HnStEX1n8gMttNluiSWhKlqRYWJkxs7Dc+DaaCz30mJeWHdr1Jw
HJAhzDaC2dsuEg1yjAUMEelG+OrkJqxnc9Gu5rmI2iCCjjDCj7G5Fzxisu5ZTFRvkzX+XZVaJr6F
3NSv7P8zjCwngjKwsFNHPbBmBTecHuO5dnhLL1NbLVRLZ5i80TGRqHLQImmM008ag6l7TqeJYjdY
mPNJFYB/vRM1No+4UqvLu5Cf41WgX70loYKVBkTsg6fDkIQqUZ09gNDG+mXsga3TIwnYlEdU3Kx+
W8g6umExmysjUl3z6jXK7IJPawqNSkyVr2JlTsgE6uChOD6bm2ravpq0HsR1qmYGmHRAJydx9js/
w1nsUzT8PiMMYyttTkgtmgIniSyfzgbLOCwsm4Xyb3RWRj1uE+qR2JauK+PnOrSDXP56Z4KpGbqM
aqknfVbkWdmcsd70AUylDiYWmRZVUbiQV/5p2BcMUFWwEga93+HjH3n2RlomS1RMVJykdrM2kS2M
7YPjS8GsAG5hYVfh7b2zjdkkpbNe0oGa4Xcj34EbABs2TYEV2eFiPdOVeRZw4NsJVMBLxrOwC/Dr
Z/lYcn61aD9GVImvhRzHpygv4a3zo64ZVCKmh2A17A0VlSq5mpNDqdsXzPsE9+5+hMcG4Ifo0o+2
xF54lku1wOBQDgx07oKY30mjy+Xr0LU76fb+2iScRdIzVRDHowg/h/CHwkgScnkxyEMqXVSRPjXM
STr6eMz7CJszK+CdM+s5pV3mfAljM9HJpYGQ9q1I543VG/ExFr6HESVhBSE1p+MNAFUXIVpUS/rI
AQL38qTWmozklw4yCIVHn//jRH7d1R9crWn5+//bSMcrpcvafYYvg4qtbST/N3ZO0GLglzHFH/RX
QP8V1NgvKv4yE3fLO/QStT9b5EVAb/qS2SddviXmFP/HP0oh2Fxl+THM2E03MrQExds4qAzj39b1
2KQLzRR6CLka/eluERUrqrGZu6xxLm0e59aArifsBQA17vDwVjGaQwRGshDOkVfMTAWYqKvwXCbR
0y4NCRmqqKtanswG6HiQXQOMhd8+ZINOXtPXI9Ov4zVgLZuAU2sOdDGxiw//FE0NoQR5O+QBt9Wz
B4bAvcl41nsRcxg4t/jbmWz3MJo2wXBNadgdevr79TIO6mLOT2P+q3YVHnb26mMkuGSZDvZeaham
zyO/7tCdiyL+yT9G2fqRafUrR56F2Dvdv96RTdq8zgPkS2BMDr0N38qST5U/bP/kPzHGbMKt5kE7
fdZwN/lTlQWT3Qy4y9SKoYxvtqjKoRPC304yLsB7d9oBLSC7gqgL51dwySLBYkgoK3+5DJ7eYI7y
zN1F6xCdigGDF/1uw3bqt4Hv3mYizIlqxOV08A+5R8b1up0AFichA6spKLfyLE6ls16BBczhqJEv
hu6f8a7BGEKtZs/CH0WLw9DGVn6zPWwyB0/Kv1gTP8lR5xXzQlJd+8s5/TRqfHY6oA3LuYT4s26/
dyL9leLZnK6bdSwYz7l5jfQHrxSElOEMBFde4ObEGYnco9mz7PS4vPuFsa6EGPwebvbvQ4VTsIVA
SS+b15tUXwhhACcHYxEW3Im/7g9iYoeIORJ3afZCT1dWHSi5KsN8AI7eSV5DN9+saXOVkKST4G9H
fMdBzSVM5k00cODKML8dNt7CZLZtttomFQFvFA2COa7PwxMR4VwE9lqAO+9DBgeB2ARagHgMsC9U
myYDyKXeVycoKdk8dNkndzNov+9sTt2Xs0gEKjbsV2ORn+uNKWvZl4Jzf+svVoviBnyASvOgOyd1
H3GCTtQ2i2zyanG291m+zM1frK7f7/Pbgr8zACmWAmUUR8fHEAHz1vehMuOmf442YHZoJVdLpb8f
BAzElMG2+CRa5u5i3WQ1MCHcYPZ2T8TBIyVNxQk2Pjc3pa3wvuYMVNlRpwB+CnjSJMAkBpzCq4Tp
kvN8u/Rr7s73d5Syvvztyq6iijhJkhjbF56AtV2Afkld6zXr1F6qPiDdJap1+/UXI+dKIDi9/9OD
bKQTvLJRUy2ahacGY50H/s7yL1b+l7GzhZRvqmhr385cZFIi8koSrkL+Ge25VsYSp10SqPxYrMHw
8kGEImOD2Y2oMJriwNvAnTY5gf0dOEpaS/KRun1bAZ5JJPImM1Zc5TS8ranskVzPonGk5+vFlDPw
f63PBj2kyMko79zgJROcjmEA9fgX101Chz8URGwOvX6vRl2JVNkFblJmIKJPM0UYdsdyS5aHGw68
j0FApq3OuAuc1c3VeD03Ghhvv89cXknNgglKNckTA609yuv9l+HlyCV7QyLCnfdWMCvomzWYmnWB
3lLxBvA81swBVqrJ7CIO4DmCOOdsgkp1XrFaz8N21ElZc4X/p/FlnTlNZJS2FmEVsfu1cQea3DQh
eh5zqLrLATVyU62gBPYHYBQjTi/e+f0qCnPEbOVUyyQPT518Zd2SuyJnWqbVE0Tw5CqMFpXLWHxf
VYasT8HBAiBHKa0uLCRQXIS6+o7qdzmAgSsnaTI8+EaIspJyw9fGSIXC4WeXJBIoVURZ41MkKgLZ
J3y6HGbGCefB//i9bn15BDq9ueFSwhJVWw+rr9Rf2QIR2z3V5ztZ1RN5kvBM6EkeyUjvFhPatTTU
dHh2unjCOR9g0u9wFNsdplT1iWMWbgiJ3Oa7nNBonwKtyxIQ7w7Wyjm2sdAmWrIdwgDhJ+WkdkLa
kuTACjvIpVR3cyrF6xVfw7DSJb+zPyLwT3WZDFzlOI0Ug2c6Eo9FN6gIMZtnQRYFt3J8gn1uqpC7
T+LcsHUD38bI47kNTgDGwZzQRjPxIt6vydNIYhzPjZGdhsExVG3pVQNDHHQInRCQDsg/Y+AwLu7K
eSQ2HCqC0n+b9vp1kVFhfXu/DApVEfDH1dwgua3WGjMFD551hagegetIL0eRt2pBJgkqUGBg6Pfp
sJwROzsZSq8/JlLCq3StW2l3Xa0AJH7IVQEnVnp1WEFbjFJLBRSYPYV2WcdqaJRMqg2+uWztfUft
U7WrSZZ3CFnES8ugC5l0YSid8+BxdTudWxowaxp8upcbzPp3H/0FPNf5WTSgmeJErPfKvpzqeYgV
flVmpmfpeuJcN5thPrCskjhQYCRisRHnk7qs1zj741VHU+85xRXvZnVVCjmwHC3K7Qlw8MAUGMjT
wUTiaBQfOXPJRBYfzJg6egbLSgPvi3O6FiVJoGIrAjWZ76QYWsCp6/xp+mIZEL6zhEi7stM3GndH
NxX32UfhFDFedmNYjZu8jJ15r1pZvSImX3CUkwT6ZFKHkOpu9ygRDGcgq4JusuxkYPWL/gFmB0dP
AgHwqud05tJ5IMIORt4jKRRvDtMhFwvmOUznFwcVOX5GmpRGXzD+luD7jOQztPmK2x3vc+2m4jRP
KP79OsfQ0a3Dn4CCm+88atbKbAbQsxj0qXeswVUoayS08oOYNwHrsTki0lEYjQLan4kYLOTMeBqd
FqoA629JiR1rMc0ua3tWd69/b+gFljJCANVZF7EqPIJqiuWaizBAS2gv/EAimrIAGl4yS2fOC/GN
zSg7VNppmEWLtgl6X93XYaC0xHVcb4l/MqemLm63xY1wLV/APqkQvT+ZOaIFEaQLkPCGbCARnqlN
QqoYuMu14rpFeJxfWNQ+b10U8iRwzn8V7wb0e/GhPxZebmSVWn/AW3/3Se6MUTKY5v5iTKWYSPmY
wm9EwYSLTWkHk/8ut5OsizOlhd3sJaaBDfRsbamoG3OQ5PjYarHE9IN2ZIGDZtMaCJmSryp4EmiT
vBj6X2anZif+Ohpw9aEw6UPjt2BZNcMISA8OPmnd0m2i45+aYD1MmLdBO6l3tSKd7et/kNHvyNLD
No4LfmsOsq6oqfsOyQ+d97kA+MMuhbSP2fRpGsXMwFGIgnrK+tWV3cYVw1a2pLgcBqukWQmxaE8S
7tl9uXq6lh0n7XPX5yF3vZiG+EYGrEcJGvCUb52M6PXgYeiF3pUNS458T0uAOoQNBF+Uo61azSYv
c9QEp9LqjiojtMKD0JT+6zlTzim2IjNNjG7HDc4FYQa49+6eVATJOGtxA+e6KaZsgHbNJBAp4MAc
67yoTlYIQnTua9MILEvhDVBlp4gc3J90I92mSdTnL1YFajy808RD0ZWGwpSv9PBy/gGtFYNksaIi
W9P1ioknTUEfrbqfI64AMsAHBZgLAtc0vvS7RcgPjqLwD64QaNMX/3zFjVGOpB6gXiV+IDeWc+Tz
uWZuKln4e6haUEbNczBjvkQvBhIoAzczyhiFiSa27CZID0nSKLgvMWTdCIi8ozfk9ysqshia1GbX
cCfHTDSrCGV4nOHsWmuuHb9GvGwwYl+0WzNmIgcmOeF2eCugE872+XwXhqNZJ8ibj58tfH7CAwq3
XFahIuI7qG+eFVCGq0DYxVhqtjf/GPMLVmgT4g0poPMun37pTKZ1IiCqcyA4ML+T/5U1MEPNaVOD
1FGMVrlw+4q7HyP+MqNAtonkdSB6y7pRwwNVy9VXQN/Xzvw0+zrQZ1EmWpEztlSWjPBflmo2Z7FW
1QJPaMnm4v2BGzUNch3ADHr9y69gJVf/6ZjCTzNyb/yBU0WBE7+IdXdcnOO6T0C0YLPgWByrR7BG
pYLBQm9CZAp17k1iNGn9QjWRclASOzZ3kgg7e46KDaOlF7d3Att0gpvMTesPP80GWGfyUJBl7mR9
omH/YY7ZYCGoCRhzHv5irXw+dcDviZjR3KtZg8fQFupChdfPmxL69t3XP2n09f762hsUGqXObnln
q+eaLiE+94kJfmkCxu8tzwLHJX2WpOvsjmAJPUWX9Uo/3VF6jBXee2gSXi+LY3XBTscjFDhv5swS
UMefrCzHLt4blBB4uAEIdA6ZeNo70G5KPXoLUYz+vtGZIf64Oq40YP/ZbFvRZoEuoJ2gdZSO2WO3
v2FwwmkEJ//hRellQFrODXv3MjUoE/fz7v9NSTCfQLFigG7ed6nIriKHZaUQUT49A/v/1d17ZYO7
hRtF4jE5nAfm9bU6wg1mgbWl5ga43GGQ/KTV7mE9zCafsRkT38QaRHMBcRZnsg/8+yiCZjinPZJJ
/BrQGhp5UYmqdfItuWAPLbjV+kB33QNkJAbgpB7OWeoMTdo3e1mC9iCU1m17BeUK4mnym5eahdiH
fYpDsL7fYHIQIqWfACDahDxR1JG0I04Yh9r8xqqZp9+9y6leKaquptpb+N6Bf6abvQajElmeQSQO
MM2pEbiNDuCug2xqMWMU0ivrDK8da9HZorx9z7jRHJ5WlHMQMrcTr0wk8HqT/nKD4EZlpHXOBtv9
oFPFmJlKk06OTdInYrPy5K1nb2kzF90RXgxwJsGLDEsPCeewerj/42FsA9BAa92DCOrm/sRQ29Uq
2mqTTI6V2eE8TjjIhyyW5WYKygc36VeTt9ru4k48696aNOix4w3HLNH9KTSaknQhfpHgyg8bnOww
S62y4Hn46pVbkRI9k9aSPhPj4BC6b+SXAAYzT/Y8fTX2M1QN+yJJDie1INJRrYK4XlCb1jTWKMan
s7+CDkW/oPF+MIF5RdJtURoaWXlrjEt8jFRlI848GEhHKUbF2A4J6eTJXoAqkGzLAGE28tOPSqgA
KekP8OIRg4uA5YPA2/RTYmiX4ORHlNqrNL72sja4tDyjh2P8LgugiS8XnwAMxZWOu058H8dt5c1o
+4I41N5ujRxbVIV06DI07Qy86sHsbQvMkTNrZ6KoXAyiTVV6cnFlOHMEaY1MOpNOpE2rLBoXet4D
v55xvtnbeoElLzfHO/34oQokwhGrsO454SLYUrE0X0gSoihLrTf6iqXHOyqMHjhb5Z3f8M8cFgWJ
vEK2lLsG3WZHIpzxuEcSEoLdErDBHHnA9KpYB9+W3e274aFGyao6rGQWiyunhoz1uSYg3w4FB3Al
Wlrw3W/vSWCq+1dpqVCRwMMRg4Hgg3GNW16LTpSSdP0/+ww+PMzelKHU1DWRpsZfDippLxPfUgqD
s+UYzS8NC6gfZsLmTGygcLy1HnYrkrxs8N8/MVvc7aM8Q4PQ7EziRSju4RJ/zopm2y6wmPy1b1mA
ZnF+jp1JM3j/7l99NEmtZDLk0n4tpaayeKqgCSjx3VLto4G0/5AylqEf73Keq6tBgJW4fQfzTIaP
7FtjvOLj/bae+8OC4+5dsGqBxm5LkVMEOthgtHdqqdK3SkOrsrVfaj2cBmUjCei4mgVMlZFpqcG3
g0wrUkAVjn2iDJk+gj5OHl1ue0tdHHsXdrRQortvLeYKyIhctjkJOleHfhMZEx7i8NQ893e5ukSS
mfCf7HeZ2nQYESSLhndjo7UQ5fEuzpBQ7dh1NhPJ9TRuPku2m5OEaeaUZXxtsfHd3gCzpLKQI00I
00pTEJQJF/knVyI2kDSTsgruP4L+TxkKYacgFyqOHTNgxbzJZCEguEb0DGKVxY53epyE0XsePD6s
TDbBexMkBke0NAO150DCKFizmUdvv4VYXOM+7A1zHj4xUmktN8DlZRzb+rNor+MdcOghPMtDTHBp
Xxvtg4UoHRCqA6wUH5LegvTuLKxrFRHgAkSmAk0e1YJeKfVg1W3mCygO4moPIrv6WrcpTUUKV8kX
HEMr5UI384QPPUdvhUHYtKGHiEAWeg7JbKzgSCLlBxSV9PJWI5bdzcz7CSw0hijQsnr5G8stzh5R
zCSr07LMh6+XrVN9tmUJIR2/NWRMQbGzhbPQblnxkKMibBgXLqco6z3PLstEau5CjP8Ab8UufJmp
NZvBz8KxyDkfte8NGX3OlBGhGZs7szpicR9hzyQhpwnuSfCyLAce3ks6wAvPLG/T46EbOsgbkXox
HMLqPGKqysTGf8vQBlPL5L8+MXmFUrQIC8iaDdbOeEp2dSvhlG2PQce2cepi1AOEa8cnaq9XQoKu
PBva30pN0DMqqxgwE8gMThNDHCZnLdqE2llWZL/R+As6fMGq9cHJvjJy9fzyi2v6yKr7bKHv4csr
NUtZGdKoGrj+B4jp9KFjrYf6uM4zv+igNy25TI4OusQybsOvrA5dTzgi7GjjCuY08a8OGr/5st6h
NreSA5oWEOhEO43n3F/4HsiL5f1EtAXbzf5Nju3rMvytJJR0oBHfSu0W1tO649QwZb7FEpLxBoru
k1GZ8h6mij1IcBZW6jXeRCqbNbiQ7lyrqmc7xr69P559Zi9LqJ8xWqfpmFk80tVrpWMaHdcTpeup
oFxLNuBoM+Si4brM6Owxz7hivMtS3luZ2FWXKDSAPiVjxt7tlDq5gOYphd7HuNpaZYw2MhG9uu6R
Hl05RSlPFUYgeHZELcai3tY63EGVwyWl6nSVh9NcVrlztqSbXspzFRn9H0TCZVsbhpEbGOHtmlF/
yH7+t5wd2+ld35pjs+s0p1/qJUs96HsnlAY5zEPUVaH9O8sgCibtCVCfo8XUqIRR/krFCRJt4/Jn
GXwMdNNu0TkLx3rXnMgRCQEMrvgOJpC2sClQvg7gZyqOcU+zhqIheBLgkP5Hx+ZGAfvDx1SgC5CH
d6S5p+42wt8fIDyZGXLzhxOlla1uX+adfEI39xchmhwZtjNXb7IXX2Gsb7/qyUPSYVYwq3MmAt4K
xndH2YT6AO71WzycroN9sOWKhquiHJhvu6rWyNqj5qwGk66Che8ZuA748OuYYUa3o8dlr+vclqjR
6evxtn5cCPvq6dPNBIgGhEoDre+3ZrP4un5F+RDIJ1Mwph/yCX0JJY6aaZDIotQnra+d2SjNboMZ
xMOVrLLuD35oAsSxPVOxpc43CEKCwWbIl/OwJ1D4Oqwxx0PJV/At9Or5hO3GWXw+9TdlN1GzHqBP
mVHDJEl8FLVHKBBFIn6baowbJcA9cCMwtt1HJtL51eHivhy1jVPuFHtu74hOKWNEJIIcx+2Quz/M
zFAnyuQx3A1sMyA6hjt+hQvtacfGN4Yp/Q1t4dODLohXBqKc0rgEtvrJv10RhPWLZcUhwQiut+AF
k0JA/DZW3EhmA/cY4aueJH7G8KJjJGV65mfSw977a7NLU24nv/JQGTidICYz6P+GNZA0PBYlemHO
EnY2QIFb4TOoLY6Fb/YA/LGiuG50pclt3MMNayxATMbpExjmKIc2yaZGNaBWXnlkFrIWww7vyPI5
vFK+QDWGcmWQfkWOzZ1JzkmunKKzi6kE1tYuVSrXJFPkWHQ9Fptx7CRER47BRQWhBKTXhSclr15+
fa5OjpigVu2A2eDE/0yTko9gLX2YU/ts2TtuSz0Q7rvDwUAwcPcs3gMg4BB1finWSheGxOtXaA+w
BNHGc/UJick+QGBw/7oHcoh/WBtGMPuSOoUn6SyRzbMwpQhLEegED8HJjtBOrxS+lE9Onxa0fYZN
QSqzYKqTJeRtF2Q+so1ichy4sv7FYGls2M1aJCIDSZ9b82Jae9GhN9ETlMKnJ52KQhOJyQzhkcd4
8otXclLUSOCclmsum9bDryXs7qqES/pv2VZ2nJ1pKQOzx5A6MPxVBCVbHug24PbhErm+vNoM4Fip
r3b9Udwmcn2dqMJncOXfar+RIrH+KB74uszG+YF4ALwTqkANGTzAMGFD1vS9jVQVHgdv86pZ02ni
iS/10/hoOT35XK2uSI2DEMNdjThBwwC95Ij4lJCsWIH3USDfJqWzDTouXz3wj6XJjs2vu1SRFrsv
9rvZlKqdPzh6cqBe2cqKsOfYjIAYqOwk+RWsxcRrfWRX9Jf96hcFdrmUzwmmZx3B0t1AebwkTffi
b3q3tGP5fxCGR0pQWT4A/9MJCUd7egAY3OyHftfVpPU5lDRsMemOFRAV+HFSeK1KLO+GsKS3Zg/U
ZZb5KQUj6BI2ES1p6RUemuOZg9TfyiafMX4xJ/64Kl70B/Dh+/s0rez9+eObbMwE1ZhjWLPPL59Y
fglxL+knTGmpTOFK8mgJEzRmh0tzkb5Mmw92Tbd2V8p196QArZH15wzAWLS55mjyaRIH+J/eSepN
85WClT0AnL44LIqbmTYG4VZd3LRGhjmGOiw53jAAc41x9P4vvRHdqGjyaO5k/wWtkVFQqGg3fUGQ
y1QW8Qqlpxinzhduwwu0R5bPiGmU7OZJjLWprZI8MnyznWva2FR3pxagSdwFfOgquZpiLsKSPI1N
J4sWFtl95a1NzUCikr/np8cikZS/6w67ZKUD2yqHE7goznq2/xpdK0WIvuGxPW6cXTtXozIhzhry
rN86S1E973gYGyr0cHdzxrM0zXHJfrrCMeACqdSZmsunomfkOT/eAfgwXKoMSpYaRz6G3QorA+BJ
B9gA1EJFJGKCS9as0d6CZo8O7T3NUOPQgykueRx05JSXI0J+cIQs0dmrNwUKfE2QlPj19tj3Svdx
hajjOLtikrZEwww8iZ/tVQuZdpYOIt54DwuWtGfwfnhw1JpN7B+Fz4o+F+g+2BfTqV7gW9GOOnBT
CyA2/9I2ZL0oVcSwpkj7wr5VwbJIkmuBX/QNI/MT4T7CxPJsefiyvxZ09egMJa1in0iB/Syg08Pb
16JqWLHP3YlikgKpkgevttUoiAmLwV5pNWJ2lcDxa3LyuwWhGuROVSnlCJLScyofKGbE8qZwvUWH
vssr2pR8CHeZKek23W/FBPJ4TueyvGlkuKdqtg0XSXDg0vGZXDJl81ZmugUPVibD8p8NWlQ8ni3q
Sz2ULm0Q9NMNCRz0PQBnhxUeLXS3mIbb8mpYaEQ7IokXJMXJ1u3v/mA+7gLrukRX3Q8rXZoHEf9d
nVnUPPEJ5nnx65sMrytZjq2inrDeXx0UoW8mmiUoJ40uoIYZ7DvLkDijKCpwGOHAsQ+UAb/ZVIdJ
UNcx/P3av0cvaNzrRwGJupizdmwErAur5fzS1/97Qol1/7BtxDZg/DBnex1JBtgCfXNNjkhsTxw3
hj1zkt3bFLF5VYO/jMXNDhIqmpmw/YAF620MSTtMoEQIT6VNWpelR88vpGPub3MDVPPFvvcXlKgl
TIzlsMk68vL5f2AHdRoddXQ1a9iKnW+JGxyZ5Q5FJn5N2AP419Gt8386o4ZxiXG1CxS3uiKJdh7y
1aYfgo24oQp1/HGWWIl9ePJeJAetq6JayraJNF6SOhvloLQyr4/co5qwxd27KrdaZV5y+ZLVu/RI
InQRjU9uQeV8grkr3VaDKdibQD+6Pv1P2hMvkvNTCZT5j/gwKpgCvMw1ZXfi2TJsyLYiUQKN75De
SAPn+pZ30ms2gX5PtP4SXu1U3v0lIDGz2nHDrG/UYyXVlx//CWkgbH6u+Q0HQwAl/6tSjfQNBhd2
f9FTFKfOXhVvkzR/aj4F18pkkJXG2WVr01dtb5TBt725RYrL49Ks1oaNezW/lLJ5YVh6qn/P+uHo
2SS6PGpxgS2JeC6p+n080a5h7jmU6F5x5S0PSeTiVc2mpuuvg9yeUJt5nNyKvzgnSXzCfymv8nvP
MCfx9hx0ZdYaL5xt0ntVaCrve/VC/2HMSL1NA/mUyUj4qK42EC7qRrkpMMojVVryWGQk/4/Eob+8
I+2hdh/uiR2kq5DNpvOXw8vNIWPoe2eStJwTsRAZVBur5dm29BET93LuXQM/pQD32nThZWOethZd
DcRMVMa8NagM+lsSyvEohUL3M50Rlp13tzvsWceHJNXcM+KAm3jcnNrj+tPCBCKlrVxi9949eK6m
6Fyi5aXkJQJl0eoKJIKjgso0CeE7os3aDKlbwTgQ8aGduSQJu2ELjBAdZ9jqUPNLC9LZ0i0TfKsy
fd5iG9NArWpfiY2J12EyqSoHAUd0CvsrF2WFIkn7WG7oGjay/wugEX9J/+bR62mzyQEhM2orKiRx
p03qkdGvYFjJ7uy/wUqx+aaOwms3gdkFf41yezyHQO1ElXCMNOFzvA62KYwtOneosygTfl68uU3c
tTF7yBAQWL8mmlUZkMR/QMHJOUv3P4THMWB8zTAz3hkgKMWYFZM4jJyQe9GyvJVyuXS6/sELXr71
YaTiSGO4UQQa3jkie5LxqE87D651lkpix6kJH1v+p092YutHit4tPFImZh0MeAiai61smIu6TBIm
h9CjjLDLMmwri/V1zBhzh9P6rDrMDmvR6ZkA23g/d6YWAOaSW4+sDq2Z1eh6GTQC7SbuTrZ9R0hr
9t3O0qkQzMZjiGKhvkGVfnlydPred7Fl0siTrb0h4x2z/ogRvMbDJezihcpKPPDd9Hu5v867dXr5
l7Vggy1u/XmquAJaF1wmLcid5efOK3MpcQ0KH6oyNajSSYkwFZ4Cy/wV3MMwU6gHC2k4uzJrfRE4
F1KvjibtPfUauaSjotD9BJIkQ2lvLqUh20SYWpOr0R2ck3ixaqP/GjKW1NZmMwAhSso/rKzRO7aq
KtFhni2snAv6vrj22w9+ma8c7SnaVTAKIxQ7OmFfoMNVN4Ycrz0sQirNKvrezrKwVH4qi4KUMFyd
SnS2Z/6VbpN9T6i3wS/0z+zjEAYfuhUSxzs4Tp1D40DSLVV6o8PUC7a/GnlTKWMb31RK2ckhncFJ
2/AtmnH5+Ah//PTiD0Xo8VCxtgOlYCrzyAuzaJtCZjRNieFccVxSig1L+3Udd/j4d/ekkFH7SITp
3Lrr1h2eYKgJYNKMa4mhjrkW2RoG3h+3xzgDFBH2DHzTJblZv7xfwCrYtVaXEQWT9WHUZwSSSR7l
FnJ05KslRrHOwZ4RTkV7KVH59rGerf2q+faA1ItGtK7EDSqW9PREtYzFwh9ZAhuQO1m1tnmbm59U
+FLN+86aLfD/ly9kC0URWA3BkH9qO137mvwEcTsv1zY4IP9A+Sue03BgyeHqYp/e2IsqED+8Tuur
bwLWb1LS2kalg45C4Vtpjuy5ijJ59dM5mloXT4Fir5zefkaPRXQgLKKLpfW8SCK5EYiE7LXhnfRs
oD89RhdAKI0DcfWkTuLLhFXRwJndwOw/8Hlhge77/AA0B8S+PmNkMqi6fELp+zD4Y0u+1g//DGCu
R1sbDb97Ez+TpEyLOfMSk1UltkLhPWePfEU8NdbAnWW1doj+noP9X3/XPV5QD95cUi0Z1/luO46w
LfGH7xmuzvbFaJWAFlm3y2qSg1kgLZnIb9+o6wIPPGIkHW7xdYmqP4d7KpLfQ3wMWfHhpoWx59hP
PCHxF2iqM71IUAbm1dFXRMtyOEwPNXy6554YmLcjqMwrkXFll2zPV4XVK/96Axw56pkD0t27UMbH
I1A04t8zgAQctWwjMdj9KZoqbCxhSwb8xF56lRliU8qTzDTCJrH4+VpMLPTYKispYLRO3Jpm+N/X
qce5iiGdY7khljlgjLv9fmkU5tQ6n+WJbZW5BekUL3viL5KvuQQ4ExWdz3lno4kT8n3sb9NOs/U5
4cJHOlFKokx9aXdo/+cvJDHGZlF3acZOHfg7Iwdr/DVnFg2+inoq7gcUBg57jkVOHFnaPVlSVMq2
9v4W3BAtfBJlWcVwfOOWvlhHdEVMD4CJL/buwvUfLhcA7RfQn9UjAx3mXh2P/wy4ww1aE72bVDaI
5qrZ+hpBVlje8esuEcqW+LHuhCaYaHBbfExeS9+4/n0d1i99rJQ6wC8WRYPAjgzc3w9qszORWb96
N4gHfJhUu+ymDaTtGEZAtl0RgbB2LemWMtNZTKArPq/SfHeWWMZnqdBNH5uW6AIsqeFGzKU92dbj
WLKw/35EM9CuEOtIxk9SdVLMveU6b8a4kl1qv+Ay3ips59URTX7CCT5NqvXk9/FhYpC58Yv8q0PB
0FfgSvFWyYdub/io5SbM1wDC9lRbWcwCzV2ByupXZ6RG+dUj2xike3+R/aJ374tnCZ7G/N+P2nV1
mv4OB5Z2CyhrLEFh9cAAzr4mFAympAkB0CtkgGoGYWvRS5Utwk2H3fWvxS2Xyn7Lz1cFW6vt04Na
01sDbp7X66rnXlsjA+SWPPXx+hB++HVrxuXQd4ZXEjizTsuWpPVDxJU2e8KS5BpT5kNeBDNaJ3cw
zznN8Ovmao3/gv5kVzihIgCWpLeoM2K8FBiUIBdk0ja3mmzL1A7Bd4rqlxTeaZ0zyzoaRE/iUQvq
RSRXXITjXBOTWzZgtAt77sZeVqe6/G8rXxZZik6IUbvWWXiD8cZLhki9NyMml2nt3otDoTfND2yO
QBh2ihNOt4ezz9DK+55Mb3J9lHBBqkw0eTs1Vjg1OdwfxeH7G+OdIfsW3RN/w2R1j9arw799er8c
wB+8RXdK1RMYW2KsOkzSXDBZ+a3nCeWvz0OJXtAUoVnA87zEYOurN2QNfrJ+wGb0iviteBx6jWSw
nZ3dHRleXC9AvGMAioYSF96YZHY82deGtjyHsJcFcCEpb5LP0nAUAVkMDBi4xUljKpArvpfZ3/Sz
X7nF5bLxMDY3sUgEaEgdVmMZ5W7FfKiH6Ny4xr90lyzoMdk4gzEzA2sQUMeIFa0Y4zEk8LIoQkQD
qoJnjIqUKXMe7XGN4P6MCYj5Ycd2zT/wPm0nwc1kYhnPNbybfDMOA+gYBZlV8VxtbqawlbVToJE2
bGnwWzMA3ZIPYZf7xn5NrXyR/eF5aPKMqAlm+BJhncvO5NhhhGp8M3JRGKrqg2HY9/IVI2lMcQIW
sXIx6gzxvypZQBtqAV0hu6HHeH6A+bmunucpRhWYB1zj9maHGkoh+2dkz29aJahrf4NwsF222AH4
ec4EaD5+opyMEqkW5daZa1IMlzz6sQNOC7ecEDQpf5U/isNr0HIz04PttCfJ8kkA1Bx7fXsE8rSM
KbGJtGIONgBKzk666OjK2XyO1g1jVo2QlSGbE4AMV7TGEqFGYQkVoLguW8APZVgQi+N9TLgFSDw7
rTBsG8LvV8LNW7RKj/eK5Phxs2aEEPzKLxrqw53lyQXMHZq7zTJJeQd9gaCzFNfl+IWYKLCAum3a
FNFLaEZ5qKGggRgAHXIMdRWO3rJrC3+Y+Rnzabm9ErjJwAFoUBl64e7NMQxh0F+6c6jrsBXUW1vC
c7OdaNWO/vM05Bs0qDlKXberxjpfjKMDTYOhb9lwpxqxCAUJuNY5Gu4zgQeXyAKtvrrbC/aBkYUs
9JnvTGLzNxvgVxHNU1Qbogoi57/4PwtPE8i8LmhD38DL7HLjfG596+gOAPKRNxNiz29miogWFGAX
Jb/HK06suJHiN/p+gjE44pwN7waA5WGYfAduQ5+lmJqGgPQj6KoBW5IwuQMFn/Z51DCvCr9EwQKj
odimnVjqX+ZHNB9Vv9CfE/AdIqae1bghOJ+SUZEfZesMFseHWmzOUnRqyhyzI9TKg2O3+5d10Vy4
6ifIksbsZu6d4rDco1MRjy/TdbsnS1mgY4GXkKQKoaEvBs5JcOIBq6cJYQL/sh/3eMlFBZULHkeF
/YOevXNBhCGaz4lleo2CRlvLzRnwT7EcIskWfUrcit9gEsaGwknYzCPGiIrjk1Tq9cUdEjYso3TD
C4ohnPBmkY09loslO4Dssojy0VnK2iqSwSthjh9p6uLWFmjkhTFikJ1ICFbXKSM3wtyv4N1ZOU49
bx99WPgOb2rCrWTpATMGVT3rM+v2ihZVZzUjt+vz0beKPD64xixjkB7iVr1Ax6r1wtxg8gDbvikJ
lKlMi9gVVGuvbbUEQP+ajNJTzKUi33RyOh8je8PCbj11/k18dovRfWb3/YbK2wzf4I8cnmXZnGTU
pMQUiFxwF5tPGlwizIjtxJGKyfUDI+TuRhtdSn0Mri4zpbgHSqU10dQxEE4vmKQ1YlShI+MOYlXa
amSDdeEvh1cd7v16Zm6DVIEi11DOTci0WUbjcSG1aDXfXgaZZV2JYiJaDLn4f2ZTYbPtb03Yj/jc
P9HmV+V21Q2iQyiVJXaFmXL55UZz798MdUctNToZ9f5/IsfOngugAs5yrjjq26YyVfiEA2t2roBH
aGKGS7usLH9pTYLXWCMgX3xj/9bSBXkCZwMIsf5FtlDtnm9aCBfZKHbDMU566f+piH4A0u/DTlq1
JDDdGz3pvWYrENirTzFTquEX5uGV7cv/GsNtt6SB1/gJG3ovt+FoeJ4zSxAx8e/k0jcpptLJ7pmX
QkJdFQRMstcxO+Kyg1tUAmglw2GL/dvb1BO+8YXbCYDXyNIjTZ4LdMBzezteBMx2TEoH2gqhujFY
WJLsRfaGx8MVV1ATVr6kw0wxZaExy8sTi00lKjCyizYHAEPWFtS0gw2tLDZouadKn16VKguM17CH
BA+ZWsmQzd73HVeiKJZJKOVB4vNzi/9Y7c8LVsEO0H7uj+QHwkn1KixSYvJ5ARMi799TdYt5oDf3
DIlQR18B7QLkHyn+2nJrqF/Ykk3E6AaJweMteTLYbok8JgICWXGTZglwBr6OqSOwlWbtmlo8+jLd
lpjj6opbtEKMm7jOwkMdZxTQcCPxukMKPlEBA5Dseyz9sI2L5SgJzrhh6Mt17Ck++4WeGLbgG6Vm
1tACod5GET932jZbEu6FwtiQmMj99pJNIB8addBNCjQx/Fk79c0YKWL0hfl4mOiEgEtZZM6y/1Xq
OpNY5/Xmv+vAGTTNL+BMzv5RkNg3tmJKlZX51g7d/sjFwbwC0Wm+FvtNjDdmFh5yVtATl/5nq11S
paXMEiBJMMiY+XSI09xCZbnA7zx3AG4iKCGndN02C6RRh49SXsRZU7V4oVykpaIzv+G5tJ44fLak
iOrF/XR4f2ZotWga+/c9oVl0HQV2D9ZClEBakFrYpHZ8Df1wQXC8clrdPkBQhlBSddrF0vLC8Ojb
JxDU4/O4ZZthOQ8WemyJ6r0aXmFL6q8kKHVTR468RAYoxeUiOt4C+WznTS3ub1dtbtZpirWRrlsm
WA1It4kQPzGMhQN8vCZihTymoe3FFFOGAWfOwtraDxvDC9pPYG10NdLAALDQO93BUYc3rDfxcR9Y
eeAKq5iIJnbm7NG4y8FL9rxP5uTndW30Cavd+mycBSKn3nI7rAHprfIwAIMmG/GHFBJjDsLVmycz
G8VYUEIbhPTEJLtqFszzW0qUm5vr8wfpEIJGau0wA/PHvYnzratrRa3MS0swHkbAiJg+1T/flVIt
yZBnTHltwB/X2qyApni13JJ2kQ/F1L3H/4/lB9PxVvr281kgZpZtbiMg8vrwqeCRwxlESKS/Aktm
XX3ELRwwxPJe7v4S4ToU2aSYwacXKOfwzYMmu6iotg+5yJHGZwzq8vjGhYAEmyn/GNyuY0Vmv25B
niU6ae4gQvd+f69ekV7urTLRDgetWpue7NdQ/e7ZiA75Ksc6rpafEsCV0KGPg/hMZ2YHlGXo8Y7C
6l+CpLs7N9KiLBjHot5eEsCYfPlXkfn/FRjxsXwJ2zHm/7Z7qIEMzM/ZoR8TeQyIw7++7D4c2m3t
z40RzaUDR5089aeJJ1RpiE2VRXR0p042v7R5mk/Mvp5zwfnF9rmyGG5DZNCO4Y28gALCn+SuexDZ
qP3uPieEJd1BQm1uSv4gN3Nd1Wc1TjQe3FQa4RSmzRWBEUStLCpl/CntpHQ8JKFoYvqvRsYD4Mo0
2LJtUs1QTbuOV3USlQeoEtZBLKdIyEVjpOuIV3U2iD8msbLOlt000+GWm1yLTEukCLPGJS8P6TgM
qrV7RgRdeH8IzQxurx0eT43zeGqm+o4JP2ZlEMqd4qCQemNl3rZIExRAQXirf+6r+LrWcZZpD2Jy
AUohrB/nOeK0xJp3SvbWltLAaJMN+WLk0XdsrSd9Qu2VI2Tg2ZEQ6mZI5XTm9XUGg7hikPhbjrvS
i3WRNKgEBrUp+D+XcV+HawdvAD6YGatR46mJSRmfr8trx6hlivmvMU8zeoysEwFHsevjEmJvWlpW
x2sxCQgQI/tU/Q0RRYTn7YNQ6H7SFIGs4XPnF4azBeh5QL1DWcHpwRQeN9rpiVCr8UichKfLzP0b
eIZHy/uU7Z2CyghOSWsqEnRzkNAo8etkiubBSo9I8DZJiQbxCdTrmhO7It91NSzouMtrFmUPyhHn
UmuqlE+3s3Dwizh6pSQkNaNuRNQUIq5SmaDsZ97b/yxt3tIcuGO3689CGmuzp8KdtQrlUS3/9Ksi
+6imvI6q3WAY0P4t/X1wnSrXJRAbSFJkH7C3ZKXdE1ohvfeV9J0nkMHRfv+jAj7T0ni2ZlC1uuDP
Ff7xa9WN4MpILtPSBIthfjrnqVSI19y6K153X/4CEPOVf4sCfuKD93e1JwxP+h0bej2AZlbdjyBF
j3qiBZM60vpaY6TF+ogoPKT6ChIwDovcYSXSPYdiWd7G2qKEspyHMtRgeYEqdapJumF9fW+yM0uq
4aHHaCb/J4m6yGKzV2RVf50T6iskdxv13xD2VzS3sHgwRBP60JRy4yCKID0m6wzrkiiOmI8LRp0U
gkNfdlJfa5i4aNXCjaKMMhVEWbIzPFd70Be8avqAJxyGDQ3UlsgZYCRzctGmqwe9TuClcKWwJ+gg
I5mcxMvnw0j9Zf3t5eoLI5121y8ZbXBE7eg1G/ry0BqBxl3oj0Oy5f1qm6H4QjR8MHW0nym65rfg
08hjZalPW0YE1haWZ+mVZMdecOL//m+fJOeeB0rsUfb/9oExCXZkfNmqf8d/O6upAqVQaarct24W
iaXFl3SI3C3XollVJuFPi+h1974BhzbM1kUdkB3dlKlJuFqXWsPTl4hpaN1BfkeoFRBpihihFNlh
RVGA9wrS8ovYFnCAO9xZ981Wu/QJY4vUTMc1p86TboqOfX32anGsOfoJGYwRVKn4doK9OK6I8WIJ
LLL9Z7LeEW5zp9p9b3Kvmv3yIlPXd42r/tBoquRdx8qlecxx6OdRzUTy8xFSrDXOw+6+tnuywjm3
iSgfpM6SqPXxiqOEiDxXp9xH2ZstOibRIq04GItpULwwzp+tqkxbm3Gp0QnWoJxtaK8WE+GGy0xp
SzbdKdslvMlyLBI3x1PtaeXqIDbykKQtFQ40/ieC12DT3UFRd0eUlesNGqb+lPJ2ytqrB8BnqCZF
zMg9Y9YbPa405aZJMtByVmHBYyQQWGSfK6gzcqoXN6ZNE4K5xhScHbO88g2xRYsM0CBzES133EbF
c/+UzFVk+YSlsJW7BYz8G4OgY50mNYQbBCg3T+y8MHETijXXIaG0qANeDWOZQD8V62HDzh9z5w5A
W+Zn1K4yhnZ8AQ8Jaj7DDJ6m4H1lzkAQ9k2r7UrWUeW8dtH9Kcou7DD1rQuNtJ7GGBxQbVkbVTXk
Eq/5b6++5N11rFBn2AQqX8/VS/hjcYYlVoL1vVuVwSKGu/zTzx7BQaD/xbP2P1avD09G3g80tTu2
dIeM6TDHVU9AWKvWTdbeopNTkFiTs54hAFaeby0caj6UliKFyUulWtU8FkhI6g0u1HRuIRbKufW5
ZsCjDv1fHgcf+xrpuW920FkqH8vBXCMm4og5IKClthgHGSsClYXkUx0AQLUOWpoGfM2be4t/YduM
/qoHIZ1SfJHPXYDZ+uUiMoExi8m+jiLHC1o6e/MaM4b5ZU+FILBzFHIROlxzT7QZXWpA1su0IWrb
uREgJtGohuL8ixFFIb522u2JGuL7QJF9Z8YvhQjOxTA7o3toOpYvCGAdFHbdY9eu9wR0ouPUVsam
30RZUHMYFY85g8Yz4CXwx9Y44bs57gYv9rIHVe8x/RJTwt7P9zhs1Rz87H8VnivCTKCsgDeuGXZz
+g7wRfd3DRsoZF9BIffCnRZCaS9lFDorvcOWv+lrQpNYxZepccqm7yZjj54b9fswfD/2tvl1kg7+
DD5i9QeAvHaq6Ev65C1Bm/CN8T3iroYVWGcO0BL/NPHMO9VYLT38rvIBPcan9k+JRaEJ/5QWDnhW
3h2W0Sa/9jlOJq3RrgE5O9mEg3rauLom6tpvfn1FpHGnPtnjPZZ2qQg/WF7LNz9vhvw02pF+4VMv
x7t39516PxogzlfSOlezQhD2jjeKVf80cph9TmfLGf08k2Qhjub+DLv6SEFWxRfZtTywwSp29Y+c
bSn2qpOiUfTNW5ZIegEQvo2Mq4HY8qAQ/zb8QFeWDx8fWj0zRe7hAAm8EsQJ2vfI/4NRv4WFVby+
dWgUGBIq1GAKwwFwxhv/4ca5Vvo5m8l7fat8qcMrmT12zUY9EIp/A6bSRLPicFrhqiYZh1wIi4Yr
Mpn8pgzLt0UKz17ANIGhUsHeibb5ot61TlWGZ8dWE3mpirScLv25cWI3lB6L41Lfe4mb63B6NwP0
d32eBbQN4xoHhmGY+LJ54M7mL1RuAmfV2GkyCee4QxNLpEdNJbVWD9IInNbMW404SGCkzmN+r3qS
YYa9mT2H3p4qcBKq3ZBlUGxLoCJRPVieTiR2R0aM8LgAtOht67BvePDssNoeq5ibYQKVLo3Zz72S
ATsexqwFiJxBLp9KpaNaO4y0YKfQWyXOSyeXjB/xf7F3B5tLy79n6Q2fSal/1FCNcSDCiC1Un17k
JOYgLDmW4ASx3Yz0Cqs7EHoGoMLlkdtNylr/BkBYea/8COgFE1BCNXYNcI2dHWj1yFQ/+hMkVtjC
XWQzkDVBGCV7OydQrOwWKVXPRFxcQwMc9um4M846SWG/NVUjbRwVVm3YlAaMNgMtJOXc9UDKUa8V
FlT+EQZFMqf8zlvJfniK5olFTz/EVLr7+Jh3ttcdmIRSI0PHSzat35AD6EpCiSSR569+H4QGPRtk
R0U9uhp9bJFL+REkxqQdnBS4YLea+vUfJUQzDt4rGnonePRLY/y17cm/qlTt4N+dOmgdy0RQucCh
E76v73PKbp+Ip0U8n54B1Z0zd5/1pMMbJL0V/57eBpGkyB1hr9HmJhMjyeosv5eH6ynhqrZQdW9m
Ijfy6zckvgQv+INeQXOvP0GRWsm6egEO+ckJ4UnPDW2bO0FKNOIhyyEafed6PWZyMQB845g9qw+C
jPB8Lk91vtxLAAi3rJgARTJVfYNUQTYbHEbDAh46hRU0VlR1OmqKHrfEGGUIl/+2LxEj0m7nGiXH
u826UCWticbJWhWUrhJd29/9H5bjcqWXmKtElIQHAGWE+ejq6/ko8Az3qdwoJ68CcZUp6vWFHj/z
iUbghY92t4PL/djjM9reru3/it9WvvLjAv1OM5U9SRHvsCPqJxSJX7Il6qKMqNDn3mSY1JklDEDa
Hmij2iUswEVh2BVZA/prJ3FEV9JGAAdzb86IWILKKIdJksKschTkwub5euGjuKVKDbYPqhuR5XRT
o/YTZQMxiJ1LsPVYa9N6Uguu830yq++/w9OCCq/YFYv1ilOUg+oPVksMCrN7e27H1rPSG8vCLRO1
YTpJbPPvNwPqhubhmoXs8PJJtCEvJ2CCfzsIo2/dljIQRzGFz2GdrrQ5rAWp8u57PHVSCT21gTCK
UvMDTcrie8I8esiCJGBmH3nLnOHJERY564JM7PxEfnxLN5W6my873MRhqOQa5S9G3TAAYhAnoAAO
MqZveusHVcmiQqVcdaHLGAUKXaUETtrWBRcFEtETQDOSsDc2bS0dfiEDl5xCkaZyGr8Ut7NobnYP
z4BPHcLwvMU21iYEcCB8l4QI9D9A/lj88JEq3z08e9ixGrJiRdrtYxH26U4pfiS/TBWIuTHNSOoQ
P504iIfKQ4WIYrsPyp0hZ0n8pIsVagkZkxBRQiey6q/oJs5MLvMjkBM50UWJzeP9mOXu19xvx4Jz
9s4JmzgKZaHCluS2D8V2RqxPqK9g400bRFztuZu5yHllFNFvvKpyn94HBzgWeCslBOGvsAdlLIJv
6EiySW9yoTeL09JKpQ7AYIma+ftvLdJTGoGRPImHe4zrzLrEnbgd4AW6bTvC+M1/z4SKpkJDB+Zh
VxEfL/NTfH+ujIN5R2ANNGTHyPqPqmthEWPv46xpSXrJq9LFU7mdagvMv+7z6Fv32ZD65SBe7eNy
Zeukto1QUwCHv9HlWWT6FOJpYAodA04L3W/VxrH+rbMrn8DRyvQJsAP+NGT96ICMpboOJGs2HNq9
a1mBcj5bHdQyzx4PVV9oxNvBYRYVfdVlqvlqsJwhXgDHxVzpHkCiufiDz7HONYUZcJQDIySOydLh
6HLnlmKA9JexjITbBq+6sa4ZX5X9BaRkN1GgzFIt+KIJe4JY1My5X+aLWaaMFfXZr0S2wRfwIca7
ii87GN+0epZrWWXhRBPBTWBcWHHDttLq0acwIw70e6/9Rgn4NHb8dRNM3zn93AXDFXExGgUB994+
m3flVRtCC2NKPbKr9kas0hFDA12C7VW1ir0BWSCJLsVV6VaRlZPop259Gs7ErHJJgul+8AVs+vk7
+90wsMpZQqEW44KkGOhhDSBWRdsBUCUvdJCu1UuBYMZzxEtD0+k5v3KQeNoqTfPnO3TJd7ECa7Fc
DhHt5LEzeDUFx8XyjFsoBHVkVelIsQXDAzg0prCsCFsBfUBMAz0FV7LU3PbGugNtCU4TGk7+YmHG
CgnBhsaGf4yXT7/JkR2+zdUzEmONWSJivWvcHSxUjJZGsWBZTZT5DMUIg3zkMCsf8xfs2rE0oxuM
wJ6Yd96MFsYDUSzRz2+BcRgsDcfSH26pryy9Kija0xUf11F2yZ21p6Xl4ImA+U9Zd9yybwtRKOwL
5hAhmO2raorNovQsU7zJIkcKR95ZgV7+Am5oT74j+0yQZITlo1uKipHBolDJ8IPQka1df0tGVltk
4LaH/eqXYZNXAbxUsRAZtoI9oG2665XPAR5D2Z07l1yaiO3V6U4Wd3iYFwppBzvqpdFYjd2uN/o7
VU9QcmSYsOW+1a8E9EbDAbjMt1nDozqhOvZBdfgYK4Lbnzxf6JLpy5pjMHPb7Gv5O6ngVj4RAPXe
HvxdV9cdMWGXbifZ5f9mlht0mptTmqx7WoRzut47JxwrMFRJWbuOKSApFrimoc+b8f8GPtk9XN26
mRSAcNVBsdlvc1tTkbxL1yxu0VwBzl/YenrZoJ9aUiYv9TIoNfbCCXQR/qHf9dA8xgAL7OwnxI4F
JqaM4bBBWHknAty8O3lB+kwlAUpjxkORcv1OD1hvaXfKXV1Fap1OCxEVP4Qh0mVj5ocA/oyjIO1b
6B3aaXmco+3qIml5cGfraejsbmcHXX8pVaYUUagrpvo9gFNHEQsu/Hn6ZZQQqdHa60tsqrcc2Tz1
ADS3g51YnhalEAuU0cuYMsnruz1w11rg12Pp17UNIkZdmN9PmRacGgF8o/u+MkA8+cfct0cw6bOj
/AmeWXKDXxjT6KjU6WyqiSnNwTbzarZ+Xaz2QA5DXLYnv7UKzH3+TihSMj6AqRGFvw9AjIw5QErT
HP7/JhUZwgsRLlpdgBgcp5qZbDl23utQ+bbNeSrhk7lwlON2Raq4mJLuCVblrDo0Zn64iZNHyYtv
kDJky8Uj2t0ZC9EQrxjME3A83xmxybZCqyH3dU8i0V+OP0EVKt9e/+dymvPeLa+PBYhZtpJMDv8f
jU2ciS74Y9Py0WW2HLTwuiJzzlMLexJJ5pjicVNJsPYernvqxMbDUvlAJdFeaJprCP+bdJmipPit
tWLYAaDkxJYRIxGy1IbDyiYl6bpLXBLgROPnBpe46KVKIQm4h3D/aQ30xKCRr5F8Dr5xb9czRKkN
JUQO1JxVw7kw88wOVBW7aNL8ijLj/Y5WWSRTih5FgMQ6P/IEg+bLCw2snrjjImfzUp7fOrMsR3Vu
H2uI+idn7oBzZmTcvFCxCwQuyislcH0ksfgezaITNq5GXuO46ttWGvYaXe++jqhjEmzmvMDrXcsw
GLCZAERzxgl5jXC2mhddq01yevE860d+G/aiXp2QmptXWVeCvF9AUHbf4a+vOgG8SeERO+l3QsrV
meDQGtqgzeda6JtTgMv5J8GsOxxmqgtuCY8y8uBwtK6ohsO1UBVKbvBn6dqOydCF2F/5kODiUsQ2
gLV899cvZ9FVbLrzK9yUVXN8mF8b7vFsyjrgkqe7BJqNFoK9aMLnpRcvR2QEvabVbj5y7FFa8uGO
eCXXgn0OkkwlS0oPSI0cyVGDsN8zJcMDHQ06fl0WJrBiY2lS0tBDJwCddgj5cCXibyzF1WlltmTn
0fH6QixQdEcCL8lXh1VZJL+OIt7f2nkqo0AzmdP/hZPdsHBNA/cWVBOXSBE5YN1NgfezrK29QqVE
V5OezixLcOvRruAEwQKQgdDElyu2wgcXh5LRuXJ4K1Taeyr4VQt1E18IGKJcukwIxi6ODUIN03hf
kSK7z/JywyDIcgT4yC1o9niabZ9IGGoCS4qVylhoydLdWM2uv5SWb/wq/4ypetB0CkqZJ9wHFb28
zYF81s9QJ9sHU+lhk9Hj22ETITYSzNCe4FvGuYv2hG7wvcgw4bXZaA5VWiGj3p0tVWNyfS1TGGyC
2mzdUeQ6OYUz0XL5Iqbq/VdPslNWhruLbsxtrHVVZWusXfRcZm77F0Q4s8Br+zymo8yyaoBIgwjg
vlS8lKcz8oSxZUcT++D1L20VLGZ67OhQo6UBMGUM9nkB4ndZjrtqYaQu3EBUzW2EyiL1Sif1xgAk
hgGTagG5b9d1fqKEzobOiCgOatYhsJYop0y/NYZWkL3F00RZNSj50J9oB4ZWJr/8GyZsaENVBPHy
xYdrnFXkcDFc5VwUhAOGV/uFaw8bjszLvItY5hKCFhUI0wd6M5zqMnjHLJS4lCTP6DyBDaW7GrI2
7zZy93UzbkObgP1lO3xjRJfkZWKgciVbc2OUF4QUD7ye1J9R5Q6pBgg2lu68Rq2r5ANWTqOxM8xQ
jdnQ5miFv3bNZEs/8eTCYKCSuCqwWt+TOQyJd8oXqSKpBASPqb7KonOHJmP6Qtp56Pyu+Zg2Bcrv
b049KpR4r5zm6EC/GpCWQJYNF5wvXU2dYLM41wJUgahEb+dsvWAOTkZm/g1SsPCSPHvTIHviuqaX
VDSLWF7uGS7fEj1VmIyCVEO5jZW2cjo7WZKzGTfjfeMQ2XEbLPUlSgCXQaX2h1ELV5CAfMMNTaCG
yg9rfefIZ/xsQhrrKo41ye1H1jdeoSMpNPv7Ac1KKjt7gum0XJBjIjyM9eO39C5FozAQ2jitaHaV
AbmxHGx/IbvLabCXhdAZZyY5kXWGtDmfMTX9duuM+OO6DHks944oRQFwXox0zkMzZFgd8tXKBQoy
+n1tguyyxDZJhVz95Xww+bdroA1GKiRTiTXgSj8TfJa5RWRErmy2HVRDsl0LxtcdHSxbc2Q9EwQ+
YlH+EMVnLHYln5alnNZDtXYQ2k8vu1oTtiYdIK9LxkHEMLy1RVyFn8U3iJqtEwBdrM7DugxOUWkx
NRDsNZcmNsh1p64L9ARafX2mEXxhFZUzM2ZlU8PfI+KliHSq5geYG/VZAW6hhFAaAyxOcg3qbK0w
2oThVQXMv/ENfr2uNd3LOFDETZyClDYznTTFpkLA9kc6uzSPipyRE3ocG74aeUrsfQjRcd0QxnV+
CiXM5/j2Kz1XP2pPq7zQyVHAjYfr3EPIWPYIh/SNvoTxXl1nRZJhODMtOrJlu22fOYcph6d6e3Z9
EMgsGNSt/wmcUOkaQyfIevOiZSDz429rxI6aJzsIcOFFJBSu0T+tWPUlDBeUQrECzRZHJX3fcDPO
3y/pFKGCl0wZCco6Tgxnxu/h/F2E1nS2TOfJwcMzRRzLGeJ6XWLCAg9Xq0xL47tucGbMU4br0cul
yMRpM1ADoU6rV7XLxj8WvyQjtSjTpfEipdjI5bdgyJR5r7GoBRHrlqXmgk+M9GjGbawFhhdapIpI
uJqtV0CZDsrKmhaEXCe72WvJUEQe7PLYYPISXbYQd6DTQ/mscoO9/gaALhwuvYfTjBLMj6mYn3q1
EUoxUXuZQnowSdsBGqbsm0ZnDITd37CFgBNO7uqH2x2f0088uR2DIIDzU91LEN9yjySIKPUGUuMs
QM/4ZQopWNGpLfrY9pC24A9fdfab1AP9aHqxGM/dH7wMZNOYVPPugRt1aJMljyx88wFcwyBNLnKX
XneWGZYQBC3TsAhgaPhWodyHoKdG3pHAICm3eqvosyOveB2ztxzspPu5tUunuBGRnYxRwuzvdgK6
ZZ4ZFnMo1hLR279WBPZS9KDGU7ArIiJOMVOsiG+tIytXvJMHm94E1hPhHOxqi6F33nShIW7FFiMN
+EgM1QKCeMsCia2Kxmm6GCGVU/2r2fQnOHDsgC4Idu1ZfYvfzglvj1zG/hXzUzT+b74FyDjJovzL
N3hSu+LC8DW2idylIyb9GFXBqM+8JA4kL3FLJNLfYo1L/farzVY5+M2atTVZaA/IFbNkA+QvyyTl
V47VNSYzDez/OSkDV92P4ys11QVxkTSj1xCjfIKOoXHXczsu245vtAeo25R8Fa4AQmreGiaPcfJd
s7DDQpszGrVBf6p3i937we+9wAi9mDYLjC/Ij7mUXs+dhiSdAxj0ns1VPPmA4x4GeO7BB86OGYO6
v7mj5gfd+PSx9X63ja+FsqdKJ66nkplNWBEAm25SoSLz1GO8DeGEtl9ySsugj4acNQRLrzIgIJFV
NIj3nk4TRTMK0NsyMC7pQYj7J/XRgrqzVC7AjJYK/YtFcb1ozeYqkRsOdU2MnJXLo7ZLwOCyQq2x
iTo+DzjDTuq7SdYPLt5owZQbuYDiHdB+phNIUkI+Y685fO/Wmpq3fj9S+BMR71qMQrsl5wxvMCTf
zTOhZa8V6BSlsjD0IwTeNH7iAcKwrqmCZWNodo0L1ffv7iqoWwqnyj7iDE3kAjd7oz30L/X36nhF
d6fi5uI/N4JX2L9np4ch6LB3wX3BNCI+bTFljsTCeW+Q5CCdmbpYXPloH/dxMseLKm9Yi/0lVUCS
4S3XZT+e/qzPDvbsseYWPkeXN6QU/Omk/emxNerl8I5LR7jiuK3+/GqEtIKo/G0CEycsmxd3sCQJ
9aKggxMgEQqC+9qBvns+gKvGVh1Q4D01eF7OtjDkYDSatrKxftsltQRZIS6r2XaG1P/cwRTfFmTf
vx8foqGHGcjdd3AG5Vp3N+SOV373JNxC6/6r9IqHVn0XvF+nEgoV0QGD6a7Fwov+rYKWewMfI4Zj
NCzPPpnFNfc4HKhWrKu1RpAgfacn6gZhlFW9NKEHT/F3UeEGoyJcjWlmaQ+YTiaBpm3jeALXk8BY
1V2O03uTZoOG7sfNMmYGrA6x57dL7IamEB+xNoUS3FKg8QlJg+EdBe35KfSOmnnmglGHduJlXoxC
pPTx/DxgVmOsG0Gd2YTtbZbgPKtDn/qB8Hbu12C9LhlMHdnfBTtFNn29NHFdo6yzd1L4YD1xoh1J
5EhgmlAJHHQMEY72C8Zx/0rydzQ7JkIlIUSyeDM5e24d+GJiXx2h13qcvAm8OCsBu1USofHZe7kz
4nzmhHwOPM2aKA0itHoG3USJIwEDeb3v56ubz0pqLlGqP2bOlKNltI2YD+UiizBML+fWI6yQ7lOs
3kOlUsm9gGwNGe47Y1UAIpCEcQjyGEN8l1SvDQt0RLKz6tG/XyjlIiqzjyU0WR2ncz5MQzdwhqnW
gu/SyCtEpoEYMkFKRTwvYvs9T2r081sqEq3Xyyt1cOLQ3pPOxaS7f+ASQb47srUkDr80IdLIgqhb
JQGDIAtPsO93/TSs135oiwrHhoyDOEuyytG95zrUixp0k7reCGDX9UptirwFhE+3/sF1MXQg8E0G
1Aa1gVRjD5ioxIQbEEBYkgbCxRMb2LwzOwleb/lfd9rKsMn59A2Of0npS7Rcs3mMM8gjmlpR0FgL
7245ChciHL1OF3a0W8HUwZREuqdrXFKmGQgNdeox0CLwFdYLn06T7YQc0a6PWKgSD6/uheujldVV
/VTG9Y+8HGLHV0PqlKvP3+OC2bPgfgUCgQJ4JaFKPg6C2HC7fweTrWXiO+rq0GE7Qsf/l5eQwjeJ
J4wf3SLfUT9TOflRt/2C3BVs8ywVVRS/ws2LomE7ai3BblC6RWeuGp5Ebrt1ehVzzkuOs72g6mI+
lfsBa5rnaCyATHt5wHYNaS8Z/PBczfFyNtmN6fSDQ/1upOdMvHm/3RlWB+Cr9J/g/U7UP7g4i3og
+19XPNYmrZMeNR40tv3I3lGGMwJAvqsbdT9bvGJGzb/R4C+sFreEWehUkGP1UgEZoTtecODHsrC9
wmGgmO9erPQgELfwC8T5NalpcDXLfefHEOidFQMXGVzQ49Q5hIBnm4zK9Lve7X53W+5XAf6HMC0b
CaIGZae2wJBWsjtAWvuPT1XJzx4+ayPuJnZYHrMHNBwqrjGaIEpJIFNEMwZQx43dAXtH4NNcC6oG
U4Vu/vXQwnXcwgPsQngoBYhM/wst/Z1O0FOxkOChn9XKlkN0P3SGXP/XiYt1RHQgtA/UxyfTMyop
cQusYilqFyE9Q1X5yMRUdQ5y76+KbWk/IYM3yfjIS+PB4ujh+GeVEB0e6Y7Z48UxFq3JQ7xgGXua
JRX3U+BxjeB2Tjon6RogjIJL11jpryEk90p8KdmOLi33jndtbtIs/srW8YZoqs0tSR+6C0loup9e
7qcUpsX3Fukraa+eFlHI+MJcRwU7uOPgoNOFDG2vts4+/Bib/iLCQyVC0kXIKPQWWA0Og9VNlRVK
BKfuBCjulKzzKPyBddiX5UhbM+KwW+h+LxW5gRi4hZaH0W1JyNPCvZcPTz+KiAAKjrhlsBlfYP0P
MB5Su4BJ3sUimbmu/wjHyxGQX/OtWv4ZeM0DuP6UWqIkak3S985xiIsiOLi9WRTxKxXZZUogsN7T
F1/MTMIKenNxZjkJQlKCIZjD3xEF7EXs4o9ByAeTfbTJl2Fh8u89zNNoZ03VmAy/d4h6lbJfAld+
hG890yBgHaMz62VSJfFlHZAvYwjvRC8Dxpnwqs98igltSHsMimNyYElDb/S7t5m0g2TWajdnoK7N
XY5aQ8dB1fRldCAbk4/uc7lha82Z6z1IV2dtn0It2Jdefjc4jGV8C5pKwZLWMm1IyWXSP2EKSnVo
vmuQZSPadubhtd+IRaMfBX7Y/eRNmqxsZ9yMCGZsDcTH1zZgtE3bRt18UAR0KID5rlv9wp2Mm4bG
6QT+qWGzCYFzrhYNfZLDwspzBbLNQaxKYFv/vsXastkNvtfEZ6Y8T9ZXp9PKD9ttpPIcdQ3qeIQj
GVSExh4yBldNqAnyLzEkcyTa62HRVvAnMdnExlK8UybBLXiZxVbIWsZYc6uFvJSWBtQ2MoRpqCcl
1i3Ms9teuQ9ByS/Gx+DEOtLVviFzHV5OKtB5c8MFkEVoKS6NzvZh4Vfcljo2AIz0EsVcP/ZdwqJt
g5pR+KYS2A4pJGjudIOyEkff++0m/pnG2FIDMDa7ObZEIijZPDp6AFz4DZ/k6SX70d7EEaguSp/4
DP35Ny19hMR+ZDJrwIlS1l9D8IjvvlVGGWk7y6qdCRGSuTNsqkkeH9Oc4AsoSBbT6Fpwxhyd7dC9
AcE6zF9Dken028AxiGNx6CxlRtyWGyqt+zY6oPM0re2kW/4gBQdLGH6oDU2RqiVF/8xirTO6T9V2
vQMri0TI/RtmzS2ZoFcTFcWb2llq/PnSDNaRpCnAqGcoOGV0Np++rjOp7TAf++aB6MB0scUWnMrG
ykXtnbLEWBCO86ZjQj45yWS5Q20O4eTZfNiQXVUGBJzu29AuzIw1nXj1n4w54x8b8+erSPWGkC/K
mL9tZ4SbwvEwG4UXMCWEvM1npS8RPY3sPOXZSrtiVDelSKdwcaVU6LvqIH6rgHAP6nV+/F7/+3EW
w3ymY8tKlljDuc30TqWVIxK3MfaUwHsEFMlRSsovVj7smt08nVF9IerBQmXWYRDdXHWLyk3iQ3WG
yXu1xY9qHz/a18sEg8P0M3iicXCpsHuMq8tbzikAPbFoxX8a02jYv6z0GEXeP+Ht7twodxmSclFN
USLPBXz1aGORTTT9qm8A9z2gQM8rOBowt8QyxFWFivyWrsS0yLohZ66Xz/4/uGndcfKAmBTu6g3e
VBLsGbm5ivqoiUPJXSZGJ2kciffpzx00zZ4jEaHjnOf7yRaEtRLe1WSMN+fJlwF2qmiRIjyD9x8e
0hcxJJcBK2vRKZcUhTyGFS+ZbKmgHxBzm4GdqeiPGTaJ/0RbEkOkPTig8LvG+TzbbiTzNVqjlgTi
8Papq6vmpSFAi4CyS/6Y1gPu0k2GOQUiv35DXlxT/TUkD3ISpRyTnt7fsQJNSPvRh+xfhyYEJRS8
k3I/NMyPR91j9mIMrncXAxwru2ZV1rjPLUrAyse9qUfJ9Ep3xjWx5J81GGyEo0gwkqcyPY7NYFFU
nXzGHRIRLMNNuyM15VDmAUTcxh90ZGhBidc4X9IosedN85n/9A+CYesfGn/IqYvy6rLqw5aderDK
pqZPhefKvQGu95jGZgrtsxItrpXVLXSfTgHek4sjd7R/S2RaYgOfaRuikpzKxap+iIs8gsfj4etk
vFXuDVZmE/PRegIvqKCZaBEZbRQE/G2IdBfMLrT9TbUoA9+0jPIYaXm8hGrOHHtHSGw0fGmkNWU/
8LwdzoFNkftnrzDLt4ZHzvu9Yedv+VAoBcje07mZSdEUfTw+g9IaMmP0xX8h2HjTa2qEovkOFUc0
4RJHBcsVHQ2V5gFIj7TpWw5oiRbWrtzNR8XOsZFB+NpKREZTckY18Rb/jxLFhB4OrKBm07E3i938
16QPkNsVvO01GnpRqn+AVpTiSC9ldVTV/jeH4f5y9d5YwK+CerbBAXndCx1LXhKNMTXV74yGdrZZ
P7M+alK0bxmgkB9FncD06rUd5qaGIa02dg4inKLrObNHpBAyo7WaFUICcwKMn14UFclxW7uExnAK
k1ezqu+VHLSuD9nRz9ooNHkC37BHvj9h8doiZ7jQ7o1PYjIFkalXQRATPRhbr42OgZY+5mg+iFTU
g9ku7K5nGE+LGcQ0pzWOy0LxvjJFjRv4qz16+gRzR9CsexQefFsmeoEPaDv74R/Vr5xrZQ8RHi7F
huGqEuwTXfPYkx27nBZzVSIHr8jZ+QnHOiEp+DwRRMA+NdascOjN4mV9hlP2QgpURyGKtNOQBh7M
5oUgurPCWYztP0cJX/ARjOfjz2fh16zD6VR7dRmW0vQYP+ALIgGXbsS3cfr4V51EDStj/HYzCF8C
ohaHfUNRf6nckE6ppridvcMYJwCdETDGl3shsHp85q/7FhhwkRKm4Ujk05wcMcjhWtc9UHNhkt1U
r116TuJwKMGgTvlBIPNn+d3FRu62lYJIJ26lic6i9k+QEjVOSuoUPRUr1KKtklen5zHALF4a/Ju0
mMX9DeqTd3zxAZHUXaMh1me9O66f+vbdSsCHcGdciU0+0Izm0gqoIrE66r0vbWv7llfwXVlq8H0G
cmvVqKr9zvN3JefmVG0Z8FfEhJvTaJxu3MpLvMyN9+UXN5T1Wgr7AjO+yR7jOuoJswK/tYqCwsNF
d6dXgvU9bJhrbzngOxubS2937ZAEwiQMbAilojMoIl6GKbcVyaSv4vFRTJsbHgoHSBr2UeXR+NEP
IvRDj5HQwlyM8jezei+/reGo5I5aKB576849oyoR/omjSqkv1AjwSkNOmeQ7eIpwcMRFeTuCFJjw
G4iL1BbsqBffpAXaL24cxPh8XiEB/1NoYQizBE4YuMxaxtvG0gC2eyiul33XNk7SEi1aayjJGJQF
bTj3X/TQ/XhDnv9qY/MrEk+iyQSqCFpgQSqY8ZYxD9FOD4x78s/sHqiIhRzdMOd1Gq+tkpdW4zln
T82K6KtJVX1IbPgdS4549pTdJlBqC94o4QFmgDTyFnLZsa/8cSeznjHXpQDbfGFQjjjsIFzlTA3l
zk/Htj5XV2A+msroovtn3akyYVi5swNbdbNOMUsDWiBIPEom8S26tPL2N0o3ZH8GVMtjlXXAL7v9
ky26KqjTWGovp88xWmVQ5CZ1rmRBspQH3FxL/T66N+IQnVgX51hWJrx1g+u1JwTgOpeuDAk/GixK
wxiO5yRooA8gMTQ3CHI+hQZv/+ZAK6jqQ+HxDzJvUR/0OvLxKHS1mIiqP57leXuvMi4I1i5T+lqZ
a6N0nA29UfeoFhh1PK2nVyN7deSAeXi5uVNvubOelTC18F3mHh8rjrPR2ANAkunwq461nRupISzR
PQ/opMDiZTje4WgMmACr/9oEd6pTJA3SFJivC5gcYRWTYku2aEYKoPPKIGPZTsV4VM9C9Am5gbnw
CAZiVS0oVbKIGqv9vuOmI3TnYSlLBVrXkJf6EhayEiU9xNRsjcN12FXwOqSDmqkHTWxz/rv+BPOa
FYLMKtcuUoaKMzMcDyrBqWBr2xvVFz4Z1bBbUVGWW4X6oZFc4LrOwgcWSxyX3ky2sySviK+WRFUz
EoyLYFcKMv/Gzca9frNSkaEg8enLQPzFMaE2XiXL0gBF0aCeZMe//vtrtqiHxKOUnmEEwT6mJzFV
IiEsU5rnN2t/t2ZEZO7EGJDQYQB2n9xppnQTIOuV9zrtUbOxgafkHAUqQhLXx3D5DFWgeMRqPv37
5xuNtLyVoGlM6LQGCDbRK7JT76qNPYNFfKk1sVXO8UgX6MLAvP9jh5MvIDXRajalMAUitAQy0dhB
CIS/UylBbNSyfBgclmUAwZ5BgyrXgwh695qmrwy9E1J78A3AFHrNSswJXol1sRWn6oRblnj7fpyp
QnrwJ2RpHs7jswVdv43KkToRYzTi1HKbl/QUGN3gCFRv4a2W49exLKiqh3NouY7asokNhvF1iuMC
YC/cMW2Y2TOU/7wH5+dzUloVEBn6BK+McoiFXCc+sDehbn9mm/p39s8CA3bA+CTHAcODuDuMGpYj
Ar2qEJzuuRx1ExVj8Fj2iL+HVYz8E4ykCCLkb1G3tnvNqpHA/FzA1Qy1GWapJQKykCoHMiJiVc8I
sVBbOSY90epQUnfImRkuCCYOn52oLng40ZKELhd3ipHK7h11HLu/SmpJTnM+e8DIqW/nuLXa781l
u8JsxsM8srNDvIGzR4Ot+ZgsVuR8UiB6q7IEk4mz+33PEHr4Rf9ZN6elYVNzPQKc1lVK04QeVuv+
fMu75OS4zaSpIymT8cDzb8tkcJKvA+1uVLnjZJeAlzV3Ch+KdqqRdzgSevp3kDi8IHMwIWSUs1Pk
Zps9fm/L+6CBIyDGsVcLbB8iqyBatthONT6RnyQHaSnAEaKtGR7vW8ZJ4tl0XsIjyqeRLpSkNYcF
A7+znqpud5bVeTbZ16DZcm1WxedN2uExndTlUgdEVl7PEsDj1Ctj0nCc9uvT+xejCdrn6oXWgQyX
oErMo/pQmYeQrorJ2Ey205SVDCMbJ9bOHQHM8lp2a22+BTj0GHYns52tJjqAnvRRZwZEQzDjlM/P
bPzw2jufhIYsYb8TfjK4xOKX+drV2pXJCIBoiD+1E6hllmZheq2VRqu3wefk6Vf/wnV0mE38VdYl
61wE0SotgV9gFRzkyvbdfSBJNbmljPCeRb2QpNWNqZQJ2yLluH0YZMsjE7lSz6SzM4P5Q05CTpIq
r6TeoLUb/sZ7OORaVUPx2x9TaLi/6attizQ/nlqgxHs2H6ipEfk8osxWp1zEsyG2gltZqa2U8/Qx
KFd10yfJcZ/EElQzltJGh9uASVkKZ+EC2m35u8gp6S7Q11eRpBiW5Us9r1w83BOEVMi609tHJcdH
mduW1UjIBCs+bsr4Oy9f4gEpBzNtMVE2il1D8wak+54FIbs/TW0Zxob3R5oPPJvHd0ZAd7wSVTRN
4lhj/BqUtzaWvIqMnwVz8WvRdvotN7+8KRDO1d3nNq6eaD+wXxq3miqpXQfOqTTZEbI26mHBnSvO
G8UULNseFJvd0MMSh4n+24yBueqp3RbhA2/cOZV0z9KdH0BEK2kzHD7xvVSK2kE54ddnCruS6l9f
UECakyIBMWOkQVQ8umv8z5wQ6gtzQCn/JWc8JWJD638JfjvHZQnw9v5OOrgTczFchrlywXmLvXfy
pNp5mf/Ms8hKuPUIE1lOVCcQPrVyn6lxTZoHe8RDQ17viq4XTlr9PiBATaX1gfw6WGDQ7x64RMhM
xJ3yM/M5VuSSq78R+FDo1rC7PanKC15siFyuTsKPyQ8McvKpxO7e2QdF8mGv8g8rl6TA0CoAuG9Z
9MNOMD1YEfX/UHpHyCvyFbbzyN7aSM0FvOpcIsqZJcA3GmLLUphqrup6F+dFZcswLchP6Xfs4rwP
2wN1/8alNPV+KzwryIpCPu53sASyJ10PZWBBsI8OYFms5eAFZUUXTEFy9t/IcFdiUUT3+BlGD+mc
bTh4kXiGJKoddT5oYx/PbGEPNg6r5myYYgKBXe7PhvwKx5y6supSyx1F6R0+xcogqSPnT3weazHD
PkvPB/6WoOSqME/EgkoXyZuXZa5ydV+vVX4mCwWgZvq1hbE173Bg3tlRpwWmml5Gs+ds1pzp0nvz
wxMqmGYSrdUZGJ0uSGB52af1SCuQhIjz/KWMboAOs6KQ5Uzh66FIeMGhjqXm7p6Sy3B4Ndp1LUVv
3keDxSdcQoVTvQK41wyX6G1JThQ0s7HFsRfWO2GlG/CGARbPPK6rc1zGQigfx27FDlcfKPRFmlfb
uvLsdwaLz4tpEa3twvjXGHA2SsAueMKttvmEAjVwf40MFkorcXmohC/T+GnM9W4bNaZXau9JhCuo
vcWwIoFLt9JEkVYndQ6vjBN0lyPja1/UbpHjrvzhQbRPzo+RQ3nUYUx+YknFPK5HzMa+vQcZo0xn
hbnR3H9YskX5iUgVT6t6o4RVQeko4NRUm52eHOkNa37MSmCNhdnCtNf0F9lHNosoORULGj6FtOOB
Vi6dpt/hMidUhocd5BZ5nnkD8JWTV24WioPtvL1DZeP/j/w0qCaEAi3hIlP/iQj0CBc6gv6wMEgV
GEfcMJ5wo5Joy+dzfzZKXtepAuVPcqsFN5bWuVukU99fwhPrXmoHP5BZCW+MhcY7gu+ZHKEKybOm
A1N7H7wi6pGqCPMFiu1k9DL2kveWOpIYPRzvTAw1/sg4ameJf/bYf8uFMZvzrRSqbbad2i6F7GqE
YfNK9ofISWFFjbfzN455SfJQ1gicvN/+eaP09FXIHmbujbwiD98wRF8SZvnR7b72e9XDRqMh7agQ
L6OulDxjs7ag6kUl/mkaeW7oL//iZtqOIH5WctxVDeyRazyLBS91Xxx1Zod9ibwm3Rg8gOvwFrCE
o9frkU2Qf+pbgfEGbMUZiFWDPqcX7VsFUZmf88ctUMce+B0u2bW3zowAJ4YrYP3UXkH8PFLm3BiC
2DIJpazh88mH6LYDjAk+VUU/hrtip5avcGG+KYr2EuJEsjxuD7c5mrebcBQOY0eF1XfWOi3cARqE
YVd5K4NQ9ZMP80iEmq1b9NaRNUAi+0uHnAw0ShFQcRxpYF6yOzR2kY8x2S5gpUPY9gT2UGdVWbss
NDhWqu0GypsFTaxbeUVZwAqaw0udsoAGq0BfEF4jCjECKSJhQoMaOCv+sJCTmnEDQgbSv91Q8C4s
SlJW9Bo7f3KyvZwpJe4Dd/LcJ1CrIEs4ZtBctOb2HID/w1DjCjKVtDlyEx5fGY1/yCirajoTVh08
zBzZ3B5HEhgrHE536s+hK8o8mgcEKriOgZYDBAWLPaSkphDkyP6YRh/7A2PFzlvEzHH2zsYnakzx
F6rPkAzNGaqTsfMIr1m5fAJqt3+L837ojVodlXxtM4kODnACNPnDkgZLNgu4n853X4LrF6T7Ls1C
azPp4YWk61b+lb0dDTgvm9P0WZ0EalZCHWW/GAGqyVt/xqeYJPgyjuNVx+k3Ii6Bs6OyGqM/aTfx
OhnV/z/+sujeamN4TAAu1xWwPGUq95mnlsDobGitHt+sepZnE5y5ksQyRmXd4NVCSXbHnrrRRHEq
HCnrSBGWow75xt+c1ifGZyNb1zud0/FCzw75JE1s1vxOfDchjx5DGksL43P7UpdeYkVi/oeB/ok8
+P7/1vCctVjBxGgDtYH+aAnB4+c5+YDxm1jWQc5ltNRU891q+q5B+1de+4LaPQR+BwiKyrGZwOx3
DYBZ86clocCa5DdAzF9pTQbMK4VXh4bY9H8tp6b1Xdlc6bXkPTsTtxLULAUgu1ogi06wFYbjui+o
FQ69tSTLCQuqyWzSg5bbdwzENGm5d3yshWuEwLRhqvPQw710a+wmN3XpDvBoQKnGkzSMQmfnSevh
QBZxoT47wWHF393B8o+1Dmn5bOG2/tBho7KXR0/5j2sGfJI9CWCCHoapDbbGmu3wYYxAUBEDTlrg
agJMbPxmuC91qbV4HGeJ8xjnvD3x2EARqF0Z5bDRP5ytisnqeexkATFyb1gaROKQNJOrxebEPu3M
ztL2yuu0oGGNOMUOd76PtRoVx3E+w5ZPUNP+RIAXCanTRBjH/VYU+rbt9+OEobN7jYmoOXTTa/Jw
wXumo4nQb19oZlAYne5yzfRDd78ZnWl41NKvajBXesGtiooyVwfN3pOTU7HwTEC4h3dCsOmlNs0E
5c8Roi1natuqpsJIblrFmMcSuuTbKZgC3bDotRK9AxGIoNQD2VbKbkjc+hbi4O0c0BQ7AExp4NSj
v236ekBKfpGcsKdj38mhzlKzoDaA+QRo5G21kTMcOBH0ywobNyB3WpnVVOOMAD6QZ+/WoTGI61f7
Wphyw1EqdAX+nOL7NjQ6ZpUmTXQmNXQwt3pBMgEOEPxxYsLStVQl8gWBDWmKN42zytT5iwJ3A14P
7lywpMZx44BNRTjO6/HqjMj0vIRa708T7DbQx/6+JgjvdvRwGAjG8XgHJy5D+TXWQ25YIfeO66e9
1yzZJtJ1RR4DkO/vNGOPD4BfWjw184LiPU22BdhrrPsoBsPmZJRbFfxKro9zJklVDMCM4DbEdl6+
omgVr6hbm7lo3D7PytIyh+AFWZoFn2S4uB4iN1R/QrkAhYFHRivEyg7x0uFW2Cro/MEERBOkpAkR
FySpifB/qEIPkxbhds4b1SIQcU3RsPyl0FqlECt7ozc7GOkMPQfLON8WjcvuyCrOXcz6qT2mTnt+
BMNyJ95qicYKWCKBcMrR7ZsGMh9Yus59OZ/Jn9q4Gf+UIKVvozPrUMUeu0THyiB1mdvmtV4udf6L
Y4GD7bpapvF6Gei2xQdJytR1xO0Na0lW5Q3yXIaC6srm5jqC3e4lI9Ue1VuVOXAbk1wKKEWMFwtj
ZpjPLILqSdNk5qb5w8bQgWH9mfVwG05lM6v0TfbVy7JI0HFKN++y1C0vCvDFNDx2VBd8JPNAoCo+
WKdKZC/xrr4RnRHer/9NB7AY4OjnO4PDUSt0fWzaj+WjTLfyLPvxob9oz9N+jHH/HcCBADJ7hAZp
q3QauLeC0bHWxjS8948fUCKlaBf5kMismuKbRh+GsWyZK2xE/Yq4HVGJiAjTkAyV3/c3+GaJQuXi
lKMT8JcRwb4N3WEXBOo/53DF3VsRu8SKZaHEONtcdOwzcwyMDi9cM9U3YESJ3+0p9lcO+10nePwc
EXVEt7kOXj6MlK0EyppWXe0KrshEg21jb+xKBLXFxvEHLlmc2szl6NbdwOqkjFXkS9owbPBMoAUM
7N1pnQ3GHBIbLWedRYKP58u1KA+mdGdA9akBFHCY9W00vfA7Rr48wj94ck/mesU5rG6vEeialZxW
SlD/6UDYe1Zoh2+TlxvGkrYeYzk3NtbTtHfnjARcertxEETxAl7yaw1eAVc0SDjUQUYO9hCihyZ4
5m6i5ULD9azzA7BEU3xYLMmaYu1pLg8Oea1NJNJXs32y0LvzXn1iZ3UYwgqY6xhbZvRHqxBafSMy
FCuIv9P0lais21qVXyqvd+iuOOdH+0spjxfX8U7LESsXJGnOf27lrRAxx2OFrO2qoOrpmwo8TYGu
Loe7yquD+htrEr6cxOUMSRAg+7KP0kgAJUkO5aED7ywayPiYBbKDPvLmn50kHmee6n+oJoPLtb2z
TveG/Vo/Esh9pgDWRS+ZYl3PSRbMcAyeZ/c3tTixxYuTcREjNoxqNT5ILyilTwdNHjlGpQqMEANn
8qe5g3TDkgHIzUyGZ9rtyqspallIxpun114stgrJmmmS8LEHWeXMDW67PdAxAfjzQ5fq/UAlkS18
mh0f7OTV/UeD2ycuF6RgqFnvv9HBEMeVcsVUbx36Qh14cgM1SaZeWLs3DmdiTMwIHglGHRVmV9Bl
C5EH8uDF964uFK6//ekKNFKCZaiDba/5IyegTXiAFKeghFcVpnZB+a0x4B757SAjTITiqLpTcJwh
s7Cty2EQuwm0aH+txjCjCgt8qaaGJnB7FGlq6chxjUI4iNBv/atN+WZEbfjYPyAU+5vGwOpqhoac
aRMIs+wwoPyyua626nuVPSNcAeimrB27ZbHYJRO5LM4TCHtjApv6DowSA3eoFTawMrHTLo4PiUAQ
rtbGlsIpgtVtgs6xXa3ImgtwV9Um4AT4fe1sxZeD3gvqit7/uADme2Yg1RmfGbgxVdGjpWgzDQWf
gtLyaOZB2CaQ5G1CEfFJAQdTA5JR2Wi1dplLC1ukCGppHzRgiT25xUTkLBij0tBoQ3fIivW8K/2o
YmQ+17YcLdh7vMqJPvajpPUwnOEWcOxG9hOpiaXxSqR7DashJs8AwYQdYCm3hJ3zlPr2lxiFNTX2
7UMWvDuRph6R2QWHCm0h1yO+gDW8qCXXczvD2rSaVukcQf8Lb8otHyU8tyKbWzvF/RI9bolsm/4Q
k/NiN+Ie0LQ+4FSMcVkcZH/WCVL3hAMG86fjkDzx5qxGTOv2ykQKN8lqTEJNIbbwIEnrvcEe0Ik0
3h4khtPnzG37U5SE6tt/lZ9TGllvm4U3pb0YwO11BXscuCrUoDCJqMEfds7RVU1B25ToXziahSwd
JyNzhLGJpbcDNo0KZOdTAjLr/5r9VBIuSFL8np0+OqHvJrsNcfessBRa+FQq2B336hI1mbXaG9Vf
kjhTSHcEazWcURt0uNm6+yTVKxwDzfm5XDSMocgDOIzsDsQOr6D5GPappt2iaxYi2IokhfFS+i0Z
8sW/DdjgGqjC5vD0/DixS29LVYkopsKVbgRc3dovaIYUIU8Z9EOdeCxfVS2oHwUUjF2v7/lFq/mf
1QY+4No4+4xUTRV5/i3YzRoSLndffhmZp9S5eq0frnLFk4aecnvaF8IuemSGbkJkFSykufMEDA2T
FblttBmPcQ0v6HA4UlDO0elcIVYAGenFYyUDGU3KfeV2AUv3fURt/kySu39j1gcpVXAtj9fp3fFa
VplBNPJbxUBvxRbDJ/3kap7O2YffJAGlSQqTo4WJ5OFQ/YnpV6JZpciLT5QOniYveiaiSIxOztpN
MY2k17nzAqSal1XKw34FOPBaZt6R+FTvZYJGJJ1ht9QfNMrNixP0/kerL+Q5TSDqFU+8Ufq/PBIJ
cBVD0L2pCe7m2REQo7LtI1qOydD7M/fwvIAUerpQ8iAFJxL60mcla/qXzEmEMjjBgeEWFbeNnisX
gpbjVxkVO2TI/EudcwEbQaPW4Ft+yr1xRCfeQFqqh9SfQmUDsN1Z8hqZl/Kzh1uzBYMjVSP0MlaY
QolIi5CFrjDeLLnSrs+AkQBXyXpV3M//djZWytjUGKDzbFB1PJsX6c1aZ/+JqpkauATBEcRQXFmK
ByKA0269xY8PrdLe5dUizRS0Owp/VIe+0qRgoh/6mUtfPWca346itAP/FIbxMw9jJujbVTg7fL8I
nsARYRLfNN+X2MLhjAOvLocecl/e3i3DLLKbcEC6eA8rsBdLZoqp/QxahUiXiNHkUdXqAkXnqt9i
Az2JoAxO2CC6/RW2BHNg8637kJncs60MNBErzRLpawTaX3QYS/X8Ut9EPICndc47+Npwc2Cvy+WL
XlM0AsKMg07Tvh+YUVi2E1FCTb/khxcYXFw0E32kDaMEjkHKXzreJtLmc7QZ6LmMLjBOjwQsMZy3
oftfPTtl2XStaDnc2WkpDsj27OsEpDrpxuXTShgH5vt3gXAqRgOXWWp31gmcRz5NTlDRIo1w1EMR
y8BAF9xkfVl4o3wiKtaIZu5O7su40bmuCQmgIc69AN6nfVZgxCYVKGOjxhq+BN3rh+7Q/o6bqhS+
KqA/zzDzYQWjtlkMA8RCiczz+KBRjgYDoGWQZbBXs6hTpK8kFNt1QVquFQoZVgUV9ZAwQ3VP224q
/xEds398yfZ4JZvybOP1+UufHEOmLYLEeclnj0Pnzh/j+u5jKe3SVUWRHCX71O4G97hXXwGxg0Xh
Z/hl1h+1nTfEJtBLxXhEDjRxht2QZvPiiqY5Bqk+aE/u+st2b/xV1cLm9QJJlppdPnC+5CWn8wQG
BnhrDlEehZkbx9qaf7UKbMrRMwXQ5UAnmM6XllQ1O1AqyF8uqO2mQSc5QrFElAEd6+hEbWDWNK9A
PGERKOD1vTy9AHPtahD5cm+tuan6KM5Y8eqYyWOGuqmu2sjLESsLmNN50agsZ5TlnamXCiSH8EhS
TDnxNOMGWCfzF29xaYWowGv0ZpSDmIqZbvOtz89ddygTJcU2MOw7fj7WOMqmuFRI4tkNAApEisO5
hOgtBkjYaEs5yuirsg9u4EmLnD3C46+Nc29hulYM/O9eIw6op3L2RlRMNR/jUXspWGBO/9doaocO
Npl8HIMtBSGhKQuUsbwoKAP6TQHxj3pIgSMasxTACR6AOny9WquQ0xUycLALI+yveTXrJ+1Oboss
7JZ5fvmfL9299o1SFOhwyK/B9/7M9oPgss9WHe4mv88r8ON3/UPe9r2xX2dxM/gPPkjTPGQsAg0A
rjNdktf+kyKFGzKlkyGtv03/trjGZGLmwmAFaUGXAgx6oqg5ybAU6QYyebiyciPqN8RJ/aDTSipK
f8syp9gStzybY9R4ovEyWxvnsQfbQz+/YZo/0+rfKd4gyOr21DhhW6N4yh12rarWj/DbulIwiPWX
iwkzl2Ia9i1xbBrmeDvWD393YD1aLXHlAj9+zG0XNPxv3dndUfgSXpkGkeVsIU6OhNAqF3e6ifHc
F/T43Nk+Mf1x2Uoizi93RCQCy1AlHnd5OqA6RuOXTaFlQVU55ZqYogmGvoCOIMScxdcEY6JCY0io
6VsbLGi4BfEF6bCu/zUdZ4WebHOQAoyEG7+DixZ1AKGFdMrsKk5Kj4XIecb2rtOm9mjMx4lq4VAj
vnCNq11vN6tS/iVidmu+YQbZ02fdzb9Lxa/RDQjGsa6UnHNo3XMobfl3IHAzPeUwkpJOzI+X666/
JFsH1GCVGx28nbr2tosWEOU3PfEWhU5/8Elzcay0IlRERHQD8mINpQeHMSkm6i72nhfm1fFdyoeO
3keFcU/w4zL5iT08whtcOBPnXORQExdkQB+aCE80azZ8E2PZeC8PHTBv8rLUIS+XwpHkqKj/9SKC
3ae3tX43JJMmJFxK4hMn2beOmtGTE+QQwddNBvz3ZTBlFN9dk5JVuOG/EDGBqxSlGxV4G+Z1Nc4Q
fJoxJ/x3XxGCuN9TTxTiVY4NlbhXNK+PDSekcY2z1vMxz05Fw+pmK5wIbJW5afVowV3iZk5evghK
IrBq3Byt698Bhc5cAnMmOVkr+Damdy7pmaptfuIVSMu7hy2EdtMAouqdSh8sO/GMkGiULE9ymIym
kxCdMaTs4I9dS7Zkztm/MhrFNSWaHxN032ZZzlNdBi9jC/gylWqHGtyjP2RlhMDPApTLggQZCUpg
2sSDgn4QEyquj8iXk2YB6ud9VJGf493j3FoPeR8Yp+rYgrAFKJpsaoVWFW+gxXCWqMYYTthB6F3S
xDZA3iyeqJrNSCJWzfNKwWlzPuTo8pkhpuAY0zAP1WbfV+3MlcZj2wX+KBoC/+lwxim3L2C2dzYV
TK8zRpL8rqpYbnmvIymdxGXdrLDDX9TfZdo6MieeoEf4UTROTQnmCOwzjOaC4deSbxMMZpDZ8gQX
uHWjhfJSNb6TclYIM7V6CbpHJfgYaAQ4WNY+fEAOKdx2kI7cjrlwTYY/MdK6xXjHkbo/5VKmmpwx
CfDqZNQkGXKt2Y9qr8VwyAXYNm3guj0UEMn7PlUYSnbfCU1tuew8xaoqxXXKmGvlKC0l2F1Q15bj
Cy4TB5It9sRJNNkfNJFORoylzp2OJP770CvySR7dkqm8t0BHe4VhSVZvxqxkvKPmvIufnnumWVhU
MlLqBvLLd0cyv0MZHEwqCytPliyZEgRRjoasEE7VzUCW9fkkjcFlEUbxwOT7uI8Hyqju5duwgFBA
4NHEIiMeMqAtApRURkPj1Qe7Qddg1z1uuPBSQDf4HtbnXN/uQIMnbpHzhHZYacx4qNzgABotm21K
e1+8LYR1VuOPB08Ub3E+kI/WCUKkwbTpp/V3ThW6rS9wFrs1Pq+73seK/biHi1aUam609FT90bZX
NvqKCoOCew3bjCZCuqQBRKbWbQDxEJ7y/cqYPrrnU/qzWf38quGMaNle41tabA9H9M/bhjoqQkG2
mp8cnZ00Jdik0tvG7ZPHo9jwx2FH0pKYKE9VGnOV5Xp7ZgImEuqtjz+qYJn9czCxoN8/E6GSuroq
TiZt44LQMhkEFek3vibPc1ehbr4aSKJ2g0FeyLwnLCclXC7CaajNGO+Q7VtPYIzWIspCcep/NEtO
b/4yl9gv275N4kOpA5AeJx/arB+IrFgDcBxVwQFbq3uPqWr93lNOAiv8stc/M8cYWw8IbD9porK9
QbMr/C5bJKqSfwyR/CyzZ8VxMjEceE/YBHb3Rx/BYG9BHQ2Hgm5rzry2itXz+mYYYxP7Kq3IRsaz
YqXIdgBW5Na3/GEwR6NZS3WsiFfqYYXcoeSTe5d01AL3mIqwgAV5tPPqz8aFNJwimQNMYPvNN/bA
cd+50/EmT46SVAOwKYeaVtxDLBv6iWpDze+DjuVexOfbdtIcxOO2xCckkAIQFjLoqck+mwa/CEWt
C/OwF8mnC4eTjSygpOcPhpIzyq+H4AyracUK+rPhzZKnjHWAuTSCyLPXHLe7NskwMuUJ0rAFtGZ6
AupEA3SwWtjn+WU+f8H8uBSUBgmU/ZUGcZA24At0rUW1jqbAWP5Q/osiU4cTgW7/DjH3JwVAy71o
cCKta94UDckxKZmxqfDRwWwGtf7YRdiehitQx1q383AicLtKMnnUiw9c5yn0RcopD+EekfJosjRP
ZIDaA5/df1qxNgj6epHnj/8d6dy26RiiUU08HR7a9HrKmnb7Ft50S7uoSC7v7aCg3tnNBLMv1XLG
p742gL5pTkxhcKsyaS4ddGEZTNWJvjHBNxHBIvGybYLFDgf3cq+2M/oTMt83yjhOoiNVCTK3ja9s
sOkPSB6FWbIygvc69DLgsa2zTL9ffkfUzUcFg6jovZ8CHxqpvQ1Khdh+dimDs20fybvNiOzmM82c
CaoJantM7bN8aY+Vah1WuVGV1+YCmss2agwnVkjPkR04WeSNdSTkLidmjKZ2V0Yldb1RpKzGGLEV
BUIlwh5GcN7RG3bFxeHl5InjA5zvCnC9vAosks9q/QZWZQvsa6THsllmP+Zc61Z1rIyH8fBDkUvI
mjQJFeOLjdQl2Cy8cVPcuvpeNVmhVdq9L6RVSGbiF8EgglYCcodKyKdYwYDT555q/Tp+a0vY0IDM
6LcQBF9iZ6qLaCv9dhGtzlSA309qFpFq2wNmHID9RnSRLsQrrOKzmKKmMhC3NFYSwXV1OIXbtrsk
nUDMyd22s2a6uShrafAF+zw5GGbpk5I24dXxY69Hj4GyPWtpN7Xb+DNT+ZBTPXCZ3PijAUsjZU4P
UE4eOFwjGHPmLeeKEsAeuSa8tAZdJ+uobManqI9nzoyFHOIqhAuJkBzIu0+ugUddKDJdH/GsxXIm
+SLJPhnp1/PYC5x1g2GxBF4vLGNZN43kwJOMa3Le8BzYVCVa2z4YHM9xatnZJov/JMi8beDgFubu
Qvtw5vyBeZMmVoYL+mjdFdrYmgJl+bxlvUvTRhzszyi0kixTO44zl3QB3qMC4p+uFMVsK5Def3qw
X47f6QGyr1KOG9A6zCLdAC+bK8i7dEzreUCVspFiz428R9GNx54bcx0UE7hkI5ffDBWpYUykDaus
QLPm8lO8Zzjy0Ow5qJ58sqT9078I0pT6tmBPeTbDum/05zAf9qGgLQrt4s006UO1L+rQgGiUlT2V
HRq9o2cDMrj5oov5oW/mRZRwauO8h5LdDU5tKqoVKgMyCAOmUGBa0+l9xi9+3DIGZPf6qLcqNFpP
gYze1m4UDNOkVrQ4/h5EG2UGNu4QF2zSlXqDoEZFgsXS0g3NdQaqwxBJg0q0jYcQT0t8mcmK7m48
KhRcCesKmlzCdzkIXLNPZZLROyb9yU6FY9qT5IUjpo5OifNJW1hdbd2pR6l3YnkR6MjyQrIacjO+
euA4s+/lq2H5Hq/jAJQQ+AuQhQhbhrf5d5BJ9KxK+pUojzONA0kNN0fJNVQzDFboucmha0Qb6fS6
P1JtrU1hxQSwFc1tuOg1qMX5gZsw+w8lFmkwiadyLT3fQwCJtNk4K0phUzjKsz6hh9M+6JSe/YuU
imWNo8M5cJjfawNLnaTUEUvnZK8+oOvVPQqqu3SCbeXnOHP14TdFPQe1JsUzIE+dUh75AQqSy5Cg
D4nI7GD7/udS8jHTr1QCrWfMUo/buNFXyvZ8Ky9o8sczoXSh5VdfV1N7sk2+pZzKW5C3yIyKE9+g
VevR0cd4IIeKG97AS4Xkb4orquREAHp4I0W5MFRWzRR/bcvX7zvsGEi8NOdHNdHs3c6gbjpOjoVN
ta2HSz03GBMeVSiuCuRM+LiHj9bvBFfnviZFXZvlpUinGAPOaKfgMenE/CQlZpFzdDIoe82adYYr
UfXwZ9VkbxM0IBegjEsvGsft2Gvli+wQt/ilVLCHGx0/FOlxo8j1cQypbpzoN2AX2puSDrQaW0bL
ZKmn9sebR75sAOe/Y/lJjBIdcqJwO3D/1ni60VW5Eq9JaoQDdmjBdY9JMIzKiCucXH/3eeC4P2wg
9tUIXtJ4TAexXsXobS0m2sg8+vxg61Od58n5w2tslAZ9EF7u99pmhPTM9u/Awsc0v2q1KmcecnrE
y/ltNWYvWz6UtwLu+IkG64bhig31vF2Gg02P72vR8+wohka9Mc91Mi3sJj0o+CmP0Z4aSfu8hqKb
H0EpynANLYcl1ISgExj5uNQ6IQnXhE0yMVLIXmvpwVJD9bHwbX53kD9Smuv6osbXCJMbnNEaA1+k
2qNlN3qgyMCQsNFICUzG8tFZc0eh0TwUCzU3qkT5+wtwntX9YdTemEAXr4aC7UdXeLFn6gnSCkBK
C22WxIdFUQ+jma4Z2s6IJzkm4m2DaoahnpaEsOGGess47AiPFKheuPG2rY8c49+YKqrD1EomkOcx
1Zmw1lxJd9Awrve24wdk0A50r+m5yUXjDX5jPMz1X9+kmBYqi5L8CJAysofkKUP5jNMpevuQSvdr
jx4stk7gGWOG0s46t3g7OjnyIMONU4jI2saEtmE3qKxmc3iOaEYdkvHETXL1ltpPd4Ar/O0OgJDY
4qmehk/br4PlBuaD7b43Hua5ecdtf14TA8lGGkb9/+Cb4OlYzO3A4a53yNTrwSq7rLvAOhxZ4MTZ
sLW8oAdxwLvsOqLWNwneKE3p3wN8Rl1+L+y5IcJn/vYHQtLeIEJ7k/3DfTWHZMRzuBtAJIh+15Ny
YTIcb11Kcw1vOUROZyNVTFXo5Zd0w9Hayl89ueWxnMosb6AidkM+LuTTCunx8LOcctMqHRRxVHoa
lDtCATVj3FHCtWb4LsrauJLHtp82sTwaFUpRwHf5gc7nfgJJaQ7sASusKBWcgoEKxrJdS6NtuzPT
8PTbGVVgDFDzxuWe9KO8VnUu6h5sKqd5GWWC5g+TMV6lLNnF09l9Qu0v2Tgmy1Wp6wPvKVnnaMjd
wa6240ja1iETqK3KfFY3hAe/t83eq0K9HrbWQpvmKAAlmk/ZBmRinOkUcaTuHNP3h7PBU1eOxJP4
K5UZrNFjChWnpJpzJIv8mS9BNZWbK4G9O9vR7YdUh1Da6DVo9HWHOG/SzfVQyai7G7seXRFtvgGB
fo7EjUvu73+ABAMQILH8TaN9WcM/EUc0hHP+91q7wkmNBgC11wXZ8qbvp8v5VAG9sXjBNj6PMvX5
yMBl6A2DW8i3NtGU/5X1BfOaRa2hwx5bTrxl/w8sjQfe9XU3B8pnnhSx9yoba7u1Ui1GuDSTKjhK
vocBOEvnU2Q/f6YobR0mPp4V+0a7vLyEf0rPqLVNo1Gd4Plnhxg/Mn+WIW5j6R1S7cOyTeyP8Kml
OX+bSucXTHme/0SzR5cfyZEEb4Cv5bgNVP/ZV6hsYf7x3kFmkjQoxCaDkNQQvfaC5glddrZZUaTf
WgVmXYA08uiyN1YCUL1xQJ9D4i9w3JDPesMJSJAe5OU/LiPykzt4yfJdaH+m/l/2uMMa4C2oO/Aj
VxY9SAkjN84kXmJXhV1SSrBk9NffvPqwjQCe3ZxTraxNy1wlN1jl4fBzHcnuzzczrQUT9HCC7MPQ
2A4UyeT9jT4zl/2S5+dmSPsT2+jEJM3S1DbWBBuUylyDnH89iCoDo6vZVRMZs1UwlUapc5a+SCPY
k6FKmhvSEZZD+fkhk+HMPXtEyqrPxktHACB8vA6TgmSgQ6t7XS27bGRIR+zTO23BOigbRwl+St8f
dTZP3CSVPyFF3K97AsMhwlJlEBGODj/pnyhsuGzR8Yg8zovt7Ds44E+isRZhTKz2z+skYLQ80+MX
LDx564SMGZY/bwBgSSVLGr5kvmleg5sHe9i7fqpfqH8Bm1wgRE3/Ao+J/eKk0xLpaVyFkIZLGfTn
VsyAWqTsu/FAD8cHK1GdBmRpyeje1g78pQgyWwTBUIDLxutakUEhRi6z9IX5IiU1iLzrveFjlpi6
yezriHc702b5wnKRwNTZMLEhpnIGi7eWpvVFsXU6QqY2LKPDT5gQIZ6DIb2F+xvN3DWM1n1692zG
6Bn2WyzMOfQMCGDj9pIMHyCKpLB5T+FpgWEIAGwx3SPcKKvNWdymRK31Bn2xQsL3LDSaHmhkABwg
P7N2WY1o2SvCkS0grP2pZuU/G3EA15gT4Oew7o/J3YUjbGI/43l5oXWD2EBpnGv1OZsnn4BZfkNg
vfmgYGOU7OgELyfR0UC+xSJrFWLKDcTnQaIk59tg3hYV/wNoynoRSPt9AQXz9FEAzrLlG7u3IxkT
ATeLLa5LMje4hN+y90kOAQYHzR3te0Jl/9HSpJhXKt58HxW8vUdr74ISdKtP+sfnk6hkukSxcjyG
E/CPqXjo/PEyVhN6NqkxzmW1jjkBE/T3eOltb5LLgBKCun7GhXzCnkgwNJPHAkOBCQargAPfZLMS
5MSJ2WcoG3252C2dld3JAjLGSHlH+IjoTHSN5MCLvf+18HmGHxofqMR37JIsOBHhUlA6AnOctWk3
jF5A2BHHHkOV19ZRJZ0VCYdkUxwYpfFo7fNgkCNzmih31KO3l4C1wIRFCv9mUOM3cOlyog5WqHaL
z+RGsmyjPuDuYfCvtIQJpXANTJ+DqlTXY/GxYpqGhLViQ6g5rI3LxlG+EhpHb+F6mUuiXQxdtjXi
5q3Xs/ihn8Z2WvA9N3pqDOMLgIJvfNov+XnYfl4t15DUPqy6CisJdwHle7kcFDjnnFrOLUTxXNE9
bGrMMJcAmjMQ5ua2ugCmydb//FnLwRcb3SORFTa/99UikKtBF2KUp9AgA0eQ0aJ5lwPbfG1E6mg/
ik3/YN8afPOVd+K21gSz3BNjRVHuiRL9E8WFDMQ969bl3ZfGD8GedgQKYbh2PqkHXrLMJSLGCpeQ
LEzw8WGL+7pSPimvmYnNb3Og4BZK5WrHluDk0FZ1VIPXvDWfesTbsmNUMAHDXMZlTFFwcsG+Yw05
z+SeiQSP3ItvHO+NDk3xgsZ4RimKvGqiPsVuF7PQHaT5GFX06IdwqzcAf11SGGtUT4Qd0Z5LbJgc
nbtFMPUUA6wajgdHyDCtKPKslPY9XdqQEnE/weQO3nDcANxQb/iInE80aowddY+fi0A0vQnul5lY
eyUnA9waBRWqphjOFsBEdsKhWtaKbUH7gaoVBW0zYEWOdPJwFyANYE0Sw4IhxM+M1O0N+T9TZSLq
B75CUkQaL0V6pfhbhQxWpiw9xr3sC/UYvV9qHxyYt9tx+L7quohlVov7xJvmvi/4BOuDuLdOzsir
YcNgiMiLa0MU+w5RcLwJSEbFUN4pLtMiJrde8mdoIC/nCiNXXJaUyDhHZjY5BtkC6CP4QMF1GTiA
IFrvtR8Jcg4GeTIIj8V43uwJ4FNFdHkkEhfi1lvdMVShoTFgx+I3IcKS/a7fsKypUpjeJBV8Z4zT
O5NUVdIMVWk4pKnpDpHlFSrKfxM0fzugjBeBVuRCc7M1m0WI5sXurfziUTPQjkz/Fn/StWGRs3RK
QVGCdV588PR2YDdhOGPaKs+Mm8nQC4bd7exWObxUlPQHEVYEfoxdmNnMoIh687Xpno04tvmitgNS
vGsd8B4nDweSKx9SA3+XraXB8UT0TLv8g0qBA5DkB/0ifkM76R7CW6Eeidi7DZowQ8vbPh311cu/
ZBuDZB0vlNBPKfQgbe8pG5VWQM1GqRRkEMw3m4ZPB7TF+R5BNyXST52voOHl4jn7RZndOymQ6BVf
Sds2PNaOXs/9KdBU46UtBPBHj60n8CF0ilnqnFEKdlgG3Z9j9kvaU2n0rdcJvxGCeGWcpRcsx6PZ
h969ozoQk3kGoJInkdA2id74tZHyLPC1x9Fr9DqsYNw1442xzo+XGrx+RKM7Oa47fnM9chcLwMeJ
NWlDWlvp5jYcSyZvdQo6uZTF/t+aFcV/2+aRrH1iKWSW6EJAPraNvZjY25fSoKvcMvRpFUA7F2tC
iJkeOwSt+cVeHhTZ1Yy5TU2As89lyvGmaU1nKXKzc99xf0onld9EZr89ktiB57m5sz1HmMvTMFpS
cMwq4qHQDfLa4MlS4Yy3VVjLB9qSL+NiriPB0hh4vmGUX2r68cy94u1NTjbjUnNiIZNP2oS8bCR6
RmA1yl7wJmAbh3ax+2kTOcai6wV857m/6Mv7YmGdMHcXdnc2webKJEokvTTfmE6iJzVG6pRmvZ22
SYsAvz4S1Q9fnRLVOTFC1lPw3le1Lb6+qe4HYXoyzxOqcW+7Sra0tK0auzUdzFcLm+bqoF44plXY
V6eDap+JHqtSQbxpRaEOxBgKwiunD85JQ/oMzGhdvuSvJzjXKaY1aAXqT5YdUds6CdXPn8rnr3Hn
f29BKgt87xBqVbZMo8TN8KoDwoj0DSSKCXv9SuT4IP3G2nTVasCcA6bu08aoJ24vdMby4W2HyuSm
7DhncTUNKfFi85DHcLsCksB9fTxpDjlWKilvvXLtqVjn7ZvB7Yv8+RivZdcdoh9xKn8m5lcULESf
Svv4ITT46YNae3vKyZ1Z6t4+cutYwNbRmwDFJFQXpPjsl843fq4vq0XzcQTxIYHLMLkQzYlAYNa8
u1F/7d9D+FViUJC+X/mnwLkaD3lvw71d/KQBE+33iGvPSYZ7u7t9ad6eGXgJ1jjzFQ/PvR8WbXRH
bcO4EOa4Vs9NqaSPPvAQJCnj95xidfWpCBJmZd5VusLTXmcL/amMRcGTzP1PaEOB4mN+HdcxEuAR
G29/Mnd8GZ0p9+p5hDjq9oqtU3kUPK8d2oSonlNGMV6wAurz177r7mpkjL+HEjb0gu+OR0y9W+A3
AArNZ4Z1/26M3cVbzMmrSRnmpIifnsUY+rhENxzV9t5TQ0BDAyycOco5QR50HkDoeZAG37rs3uDW
75q8zHi9PlDgHYn8gxg/eMltvPRVgcvhSF9S5a9ZbNMAaAjZqN07It76xfrDF1M9Xz5xcON8FOpS
BnFwcYqc0usVO7erblnA9JoEIJwUjkYjZ/ktLCGe3TJV/0zIsxM8JgO5TYZPpaSneXerM1SMVWbn
meOICdQRq+ZwtWp9hly4mto3maut7S+OELuj5v+aXnwzXq0PHaU0wtlJdnzFV2DmrKkpv8oeiJh3
qnaZ7hLOEsWytZcbFQC9OzAr7M6PbqqI+lwYr0XWmN7/lVfyb7KaNki3Yu9KkEkoy/91zZ7ZSBcZ
/Vu+xaWrx9FI9twuvM1KedY3Iwjn0EKcEPB2M5e24BHLEb1oFVCdxbLZExJ6GO6aumlWwE/TSF/p
2OEbHY0j1DNEyAhh+UOBl+jNRkiFFGE6CQjF4/+oD0V7U+2AIIEgbxQ93dAjUDda4DIG79/XBaBF
JPh2aoilHqYnN+evhrk7Q1QFUARu0bsuyvnFXrHKNvxHyJbI6RJE7BEapLhDUvUx+0KqpqEMliIy
pTqgw8UMgJR2RRKXArqhAgF3MFkre/DDfTZmeKJQt33QYiXCGzmTrFflh6HQ3s0LOnsO20mr5crs
CoeIHqLTkeTTpQVtRbzut9dxCZWU9lVY39305FIJnDNCYeVONl3469xYfrtZ9GySA9T5ux4tpTxF
nb6wuP588YwKj403ApCfGWdg93Yky5pz1/6mjv7c64vuwJLapplH4zr+YeAF1d2FJ/X1HNn8zJG7
qE6mImMuyGnXhEh6EKuhKRt6P0GMsZSu+63o58RPB3/e9jl1WgB7T5ojda/cLJlqFaoOdAdPm9Og
CV4N0JbQXspFVA6cTRoOglTdm/MKYhdHg5/fDH9tW/VWdbOtyDLPb0zLKAosywrjEoFYCcu7VCTE
IrpUXBqgGHMac9uLa7FNTv2c/on7fJ2Sv/n34aBlE1kfYGgylY1Jqz4ZR78ESHetulqwDXf+3sO9
KEPDMr05Fpkk1t5W6T8xFCt2uNrkANjSly0ohy2EJi27s3J2nhoOMzgoexNtAuaOFevXDQgwNqrq
xnm7l40g++xgjpl5wVcJD0i9RIWL9oQc0o2ZOWj3m5eA6ufGrLVa3DcDW7YiPPhARatjMfHfXgc8
uHLiatGa8XLqfCP0/TJU9L2aQCaZ8sCbLGeL1Djk0VxqLxJahecnfmwPrG0zxLy3aDIY+MSdq1S+
2F6BcUlv+ZhgH7vxhMe7xNSAroMOznueM1N5r2Q2xSOOJJLFw0vZEH2vo0YrNh8ozMKU1PamEfqp
DrOwNbIV7seumQn/ul3xgH2tuevqwfO0F/Z0emXJ4S7/TRS2R96mpJ9z1a9R3WVQEmFpOB3KFZDy
9Xh7BHXyP4iYD0A2R88ILjAjl4vy/Gub0AcqQpFoEwlB02nD6MHyvK+7jGjJ8P4zSFx/magB0Plp
q0f4qMKxRFlvSV23HTJdayaY4ujkEgsCCUMptuuGY4GxgPtnlZzELsGJXr8vzTMDT/R5BpgmsrlE
goLO9lfQn+3aWrwRJ801pBEV7xQAV/IrZsp9tp5Mh3V3gJkvwD6cb+kuAQWQwtaCBiO56qB2IRhM
fbwytdN7JICs4LZGm9hDIYAmWo36ySF2nNDdkRqPAySP/ny0KuGMGYHvIXVEtcZuQZIwWmxMV5Pq
MG1oWq8vRdim6AdtBgPjU3ikQFH6WLJQvS1swMqSoD9s9+Y44U+BbElDEXn4qtKmz0U18t+uBh7E
KUeFJq2bYRMDmUklUZwhHmA4bM1cbuDJQ4S0m+TC7YC6bUnLn/4cquyQPVZLrtB+4rSGwjKRALvo
kfyt7NZXEGWPgv05r77wUZJhw6cklylLoreehOBZXqJjbCI7Ov83nt3QaKmpU5g7xjIoefPFZkzS
52+vKxltQjiWPLf5NFzqW5h7vv/M8CvxM+EpOADmBp+GhvjkcmJuHdT65poeP+lPbr1MDxfS8mzO
BFtP3AHaSoG187CspUJDIcU95ypdSGoCnVat1+ClgOMjFrjRgUAxFoMD/J1c0xwETmvrXGYCeufQ
xGCE3pnTbaER304llQ4ZL56Ch9PEjTwXmWicJIecKyxrApUIAXQqmZP7aAFq4HP6/9TSBh0pPPPg
8BBYPWNnkM2FznkkLJu/hUaZhMe0dAeB7OwMJmECSQRAZM2LTH+2LOGJzxwxHf/O6NWpWIsDbcrh
j1UtdqeSE2Aax833S8dtSRSiLqwgCXTVNh8yaQQ/b8VZDRXHT7Gk9WU0yIMF/PBv9ZGIkDUHv71L
9xJKTedSAMyGgvh42Vr6ZxZNM/zItE0GSy9UFSfH7Er4eKcb+pamdFVJ0MHxua0Y+0k5JhAcWiiU
sdqthCXI4omi329tdDASU52h9UtITf1Lrg5HIoChYfeUW7WEUew0sr/pCYIevw9p6H0OAVo/flqa
BjTt+lM77EH3gP3RjnRcmm40CeIhEpa38D+EgEuBixm+qwooZI337QZ1cjG93gXtCyYzhJZ6bCfK
u7wsiL5TTs3nGHQ29XH5u/27m80cPAg4fqKIru7cIaYiUh+VbdPe9ASgVZAuHDYf7X1pugHikyMU
IxLfInpI3gHG+s1RU7vLz5PoS/ySnsRtHHy6ajUhYXpEkL+LrrTyKULNfpHRcU53s6z+pJGEUm6J
WBWTk8Y5OC9X/RkdFOZicnKuKuraAWDljlqCABkcVkdwdM8FUipUJagkVvSOyNniorq7birwEddj
jzUVa8qz8ixxKRrm4a/2Helpt+uX6HvipzXeKZ0Fxisry2zk0uJQWEcRFUcJtMA0fgwIHKR2eHQa
IbvByxD+9fWMLFJ4PaI16UFAqDi9HS13V3Y2yfFbKbQhVQsVE8D8wpA/LwF99sh3/c+7PoABcnME
eqmh1U/2AK5FE17j6YJ2MaWYNQh/iuttvcvadX1ETxo5BtbzkF67vC2DykoovZf4cuvSZajhloUy
EtT2kBC+DghQ4K3JgR6b9CNIuGj4/oZZbkyLVYxP0sSFrWhpLkY20vbBpEnLwxASL7ufFNSbOWnh
PKL4H4Kj49yWK77ulfGyvRjw2Zxe+k8dC8pAjhlL9K36cgNijwc+Q6ptckRRSAuBEgaYFPW+w/fU
H3qcTe75MSivoU8m48iLGjCqgRZln4jL204ZUj4aDF2Xg01qn0t18EKfcXJX2DpENHHESd+JkgIv
6NsjdvKsm4MtTVpLGuKmte3pSThTsaS487TnNICrtizAGbupyo2YEIDAMmoWLmyxMv1V6rm4u0H7
AxrhEneCemQaF4h6/ZdpDKavqb89q8FpWcQ/e/z7BIuhnI9M8lfLV6YOS4Zn7K56UiA6gmYTRPWE
jCtWOft6bZ4lteRYzFsfACYdPZJ8F5WgGupvcITgqZEXs2a6q1EfVG7pvvjQUjk7oMcxGHfNfJaR
TEkXHhWGnUlHwXORVz5Berif6eJvwYTT8BbtKLPvq+wVlCFd+5YxUSU0mNKvypTbqsoK4jC95OO1
9hoc/EgmWprcnG9NInc1zJiyoFdiP/YHB0vo+pXRu4WTWIvrHDBYnL2m3meD3U4RAzwcYwJ+pQsd
sGNCRDmOpRb213G2P5kd0l0wwy6lcKC2Gs3Q0dx7b5FZVFD066q4BwgpvT+QCDbGFs7OAD2RMVPG
jXc9t/xlAj3tNnZIVKvTN6u1ci+RpEAIaRQr/u3asdlSF9GzphieSGrFBRoDa2gydYyOB+IHACYY
eCC9ACJ6T/zENnrDPlfY5CpGsikRd3IppKg2r/prANwPO2vfzFzLvfJlwaUVBSk0wlhqaaSuurZ4
Vp4PfgUYsFzVxP4t/K6ac7zx0QZpAL9SDVRsyvfycv5oFXeHcEFAMAaSSvLo/SfuyWlmb5zis4hu
FNJG5W7XWD0CleqzxmmPiOoB7/AMgxzqXTD+49iZpHeuHHfhukgdXIub9QYmYS+FGXentzElcnsB
QvNqqVk3/q+aq3mT2NErZeIcZvXJbGrucm0IkbX6iLhEsH5tTlNMk98C5JthHqgqRYjcaej6mcCe
DL6+0m/LrXAaQLUSvFMNfPUYv3OLghlR717oEa3b0u+FE08ebTo4immNYU8c02isUTNnJGIyoGdA
EhFEeOdNZjaiYcqNBFG4RgijSkhWSJyb4qJR2qzjq+/vaUjjVS8hFkoGfUadVNa4NQhY+v1Jjo+k
o4LXSWa4hMnGXZPA/S+0rZXQd1iSUiUFv6SotwEnjx9o3CwXjrdiGbZlYoNUAoGhku11SCUc/Sfm
7gXH2BMkknk2WJ5pnjfSQQ/gqqNVXoPMINAFYjdUJSFYi2IDsPsg7e0x8WCTj8fOoXwTKpPM/4wx
UGfS+lHS3KDGZkZmrZWdhGIorh0wmq32noRA7XDMI6Cy6poE4lBbDow5Zy+BZD7zsastb7Cq4FvA
wXVRe49fgXHa16ghN7G9uYWOw2aaRdpVgyuKKY2/gy9AL2AZ+jKaibbxiOQaSV1EddUlGPv3IAEF
1BQ4JffOhaaFB1LqZxpyRZhEJ9NXtgF8RohjfIBfRyNRYyRZTeelgwhEBVwRK37q5FKOJT9K36hP
LZZyBr0PPHPbeNl0YE186Vt4hXnNPX3+aT6Aqjx0yBENBWSAWJLi1YrkNg9R/YpTPnaOrLVBWsRk
vOiyDQV14gXuqB6hXIKIASiQJzoB8yn9qtG7D7GizI4mPIxoiWfTlIrMM5qayXRZUJwikxrlJv9y
06Ku9vJcRAuczG14xExDHt0vdnlEOY/CR+oAMx2qkGyT3KCdloR8pDW7mPaJhYdie075xgEnPC6Q
FwLND2uN8UlayMWCfgeiW6mUxDyypyIsTIeLg+NsFJKLSEToKsGNqKJHScrU+El6M+m0ii181m54
0Qp4Xt2yoTsN228qeAg5+8djiNJpgkuA8exIIc6zLhnVC1IcAft9Ho3tLNKprXBVD2kXpIDTY86H
FDAi6HCjz9/R5oGeXGiLyDbxghgQedDUnDT7ybyF3mPxEZqlgOkKDHWet/HbfdUmVHnMFh8+vP6u
Vmorj4nqMVrAgs4vejsGF56vwgYqHwqToYZdNuWLnjKThfwGIwx1bDEt7DqyDNgfgbY0C6T6wc/F
1GzYJ4EK8otP9+Mn0244HnzblTNG9DVG6qxhFOGEqPGDmRO7ZZ2ZuX5rCSGJt39890Spya3ta+Cx
dFLQOGlHRiSbESx47D8UqA38Qp4jzzFPaW7/teRYau/NRHlxJWEflcrD6KUeVOOCR/84fPoN5aP8
MvVQR+T13h8G95rwd38uft+9C4UecvjS/z5IaGgpX+KejCK0FGysel75gVfepMtdjFbtOF5SCklJ
DlRtFJQCyCo+1la7HFCbvyKSHmrtFBK/tsLhKL1q70svQoubICcTbsKKRHOJOKlEWn9e2w3e8dbv
BB2Izcy2Wbh+EBn3K5J+/I9AzGVTe4IoVRTDInMQUdKABZdmzZfA9WuLX5+jy9RKDAUh4xisZgc9
2oAJMrO+NOM7j6kyKae3OSaQq0misWpHCSCcqvl4iC+8wKNAVzrp+1+UGo++2szy0B0k8Gn5eobs
4QKJwxttu8LWMA0+IETUDBDmTYLcZUOTiVoSrq++2WLGeQQ9Oqr8Y+Ke+xCiDS6FzWtcZPMqnPLf
kCKRHMrg/YKkufu8jaBaeGn3i9TS78ThPQ9TkPuLUn+iNXCn0P2ZOgu65GAxtgaDUbySOp2Hmj0g
qi/DC4ejB1PalIMHK2LCrkkbc/HNO6W3DbVav8VMpejoSaTLSD3JHQ6IV7RlFqoYDAyjEUQavnUK
X+K8Iv+BpCR7tZGk0jqpDcBFdE4Uc9wmZ08XLfUhGL54aBce/XyW/3UIx6A1aLRfgDNdJ38SCvVi
ZuUgrjYB+40LNh8Y8TUIgkdNTsiWal1xPEDLpRYXWUBCWm1mKuB8VDrkdKlhZ9t/3/dTJbwUGZ6v
5JQZ+FfCxeIN4xhyFZoAOIaZcf4mXwYecdxzjr9aOMFmiUOMMiV5MrDBMwjum0mf3qR5kWowoZve
0agS3G0WpqDaMWQ94fdNK3tnVD7FHwjVQTino1RlXOF1ZwZUfBA++wDTWyFbRmPSn0rqm2TdJAYA
5RG3W+Y9r7coM9x6gjYrRHWuCkWlKkr52IBYOw/dAcRgtmNnU+iM3+llIXizJ38I77XGHpoEBPrV
wxOxRFCnQKMqs7U0jLO+v0B0BUzwiEIbF9LKQzniG7w3D6JLKBSH41lVTbhy5PkYfx9XqusIXGT7
GsE4sLAz6vbYGyShopAbJorSMwvKQENMC9jhILWgkiCDJSq4SipE+EWaff8FICNly2xAYyZFhxQh
39vu8QqQMMBz3vwdC59Jsvt9qzHD1t2UGpT18KSI0s+8AUjy0OvIphUHunVgO5qkA1HRg5HWcWtX
CUFZo5slMGogee3A0qy88pWd88/UVDlOdjPj2FUnArUCx+92gD/VEshH/vgsvO80T9ohDLNuGyFR
mW5yo/56cn3U6fKupmWIIT31pmY9UAhpIr2fOb8Y/tZ9aOZc73ge6B8L1DmaUIRAYasGYEZB07KQ
VVyuLedbGFlwxsr3UCorcbazfNq+zWTw4DdR/ApNaQ9eSwcP1BXfwqVbXxIG0mE+SPY3F+J2S0EC
G3T+CWEMjpWmGDSjvfhjvbK5ujKTqPhBi7+Uq634K/QXLSyQufrQT30tZZC+Db6x3yXoLp4K3fbs
9mMOYOzB+ZtB2nWYdFvQdyMcX4I5C1/6uLzXMKptPSVX3zmWr8qnsSEA9IJfBpLEhNf/zD1SFsdD
kV/HAcKYC0IWcpwFiEuz6iqxT2RnhrS+TZ1NkJ6155dWmXneS6xQqbki6VJa9br4vK30smK1wImI
aVCsjJ+fBywpZhLVZpDxNp3H7z+wgeGoQny/WemPcA13LqR0wIa9dwLZeSGVJd99540DpFo8k+3v
9dlix8bpmjXqATch8GEOKXnzp1+ccywkd1t7oHHTvE7LlIU/RqYPFyXptYofvka70LHeGI5e9NCM
1ykEqtroDAAdP04fBh9DGtg1w57Pxf2vnKb29F1e0kwyyM9QnP1sf64E7MYyFujSsNIUjmAxPxVf
PR8r5sxIrePfiZ9XBMSdu5gBRP45WBlGbq1Kf2VaevECBQP/MD/pTXIpbyQpQNErIYzxQY/ht9a0
v8gT7HRDnz1coVcNYsrV8Tni9LTmrspQKLNb96M3VE5B/3tdtur3DIsyicBl++zVdmnfdu5j7Eti
DPBIsM1QwZ6JbCAM/UQLsfQgfq1scUHR1OEavlC5auC3bv4tO3ICR/bdiqqKfeKEuRddV2k12tPa
Zbq4GyTx5ZO80hqTdXPi47mNLB5gy6wtf1ZQp6zcKj3RPhAbA/hg4pNjAsxGY69wk9Cqn3kcM5Ds
tbafTN5U7/Sf0QbkrY5BEc2AnHItITVeKr6DCsCOPDL6zmP2dnm8AB4aIMnL44sCKOc4a1eiOYqJ
zpzke9UmW7eAZ8083QL/u/jI2pMoORABNEv9O43dJaDXYCnSo4Fu64iK37QzBmJEhFfid4CeYyg3
EQhgqrwIw3fXbO2K4vvR06qNjOKdtiK8NFnpNamcCUJv/G9T/eyiLlIPbje+GrUSaoTxopu8CLdw
i9CdRJU5GVSPECaQSF44W5fWPEnZJovHMEGFjADRt1Ngti1P63YhrzUi5I70nr1IVFbxJgxlnpCL
embkr0itYJwoP8MLYfOoZI1dKubYNYVq0V7WQiSICbgB+9tog3329DvFc0MOVYsBP+ZshEScWdax
NGpb8dSOMjeR2w/3QUg6VglJwyr60/rSsFx146nbFqjmLWZL/3Gy7sjUFeLppD7uhycH2D+KlFeA
7Vh9a+GZkXI7W+CPJMa/1ZxalvyM7pS5mZCvdROrYgCPcs2yuwhWkARLqz5RyegjShLGV+0LgHiA
DI8k91fJty/rbTihLm4Z2rIr2YDaPi6p7vr9kWi4T/pDaI6eSffy2c7NHcdRO5hPzbhubV/uOA9s
9NtkPO/ES7lQyBKddrgz9yJbwO8VTWjnPrdU43spZMKibzgUowXVtjsHF/regrmvMroBXc47CD6a
IDHlYpoAWlEt845iFU4O0exoNPJqJvnao6MGnvWwFBkaM0HSAuMyOAKP7WuoV1YaJ9inmS8hM58t
O3V0ULgUe45toZWg0UNlSDvaU3+DybqK/4Y59raYgrOmH7esNBr0CWvdntmhjn2mXtKCF/d/861+
gLs6t1cA8u9M6Q1VmDdbf+M4OWp8ONhpjgfRpKfjks7dSADulQSMxcW+yF1x/bPDSCYOnL2fCvF9
bH5thMEJIZ1ZTBdTbyZnY94Fly69Ymu7nBuf7S6OIHdRkCUP1vuZTvQVmu0dsfhUnl8cuIX+qvDn
oubscmgC/V5daywr59w8AWz+i/LqSZCOegRTqMlASNhhQsKV64nM5iSJSE+IwEUZ7YtOH9Pae/Nd
mSvmJ6zQgdLSp40JmmZBdkVI/fU0iBt1jxe+EqJXsbedfoOva8W50xN1yc3fCHu2+Ph6ZtHmvjA9
Bqup0xhVEu8PedP3G+lXlqgZ5w899g+gfVFlJd2JKUiIR6tHrXTRtULs4F7iB8JwlYWvtOYupyiW
/I6AXyPRGrK5d1AUzEnikhrW99IqKRC70/u5y+2Eo1LvoaLbigjgDUFZAhVXBX8rjBhEyvWsDg/h
LKAbP2LYNG8ycMvXvmK3JK896QGLjeI6IhMTWVUjzEuyg8ILAFp0rDcUk9F7MpKW/5YXzL8nzM2D
ldjdxNVAaDJLfvDtBFDZubx3WDrG2P095cHf9FM8E+SOR3Mqxiu/b972RMSK+yt2W79cbsvEBh9o
gFtXV4kqFN74q2VOYzAf5nhNV9+yUIPw0Ni2wI4DRDCjRXAuUtYzRFV6N2ocdtpkxidfaHahtL7K
TiDaZFeTu6r5X/rC2AsA4M5G56vkM910+Esptq/CHPnjauHGlqr0lGMcG8VNS/BSLskMVhToEcJ3
5rolxrpXWrE4Viy7OtbPLnDbkyswxBY22191QAiJSqEFsDDkjbrBtRN8BQsfzL4SEZf89Qx9rEEd
Ko6CveiS3l6XUwLkpB0ZZ1ivtPrYwTtj2iw7AhQncOQ16n8BVepVNpxVjBErbPJaFpDnLBg8PKJ3
KQ1+h0wGEZqkzBvNvtwusxB6d0qPVfz5NP/yK0sJ3lI0npLsJtj3wtLNQd1+CvzZCCgStm5NCunV
OG7s3oG0O4Q+ggctct60IUl+ERYr5Y/1XHbQpydNKegLT5I4LQgKmBip3aFPpaEMG/MkDD+nw5jx
e5K5cdbGaojQFUV/WqbvwA7ZXDimPB5deBgLXm4qUhrMfyC3+cZFUG5ocjymUyqGOz3CnneE4P6y
2TnqpmTYqc8yrcjcdtzyUEhZZ+19MHey1hh56nUutMr9WCanPgvULRI1UBHGKATexDQfvIpSjygv
hNOlNwiXqGgnomP4FNeAb5AYHgdCE+CcN/UcIfT8FOQhdqyFQZaOWs6TCO5xWZtg9+dumSs7oFc2
VRvfTwX914n31jDlK4PJHr8HjUzh3J/JHJsykNUqv57p4VP2PAwWplpo76EK+Bfh639OGFgtByl1
UAZsX+2zXDkzjVvEcS6NeL5LhvYraQJErZjH+0DTvOb/xCNesSJuDbHpPThPVzjs0Zhn5kDcKpPC
E/321O7TRaxj2dQjy5NIPOYoRy4iFTbL3Im/bC5Jf0RWg82LRqWWgmuAmdQlWoKSTf+QZufJ7iDr
6OpL7M2OLFN79/xZOOaOvPF0O6zYYJbDIHbadY8FaRiVbLp54s01XThPTCg1Uf3Z3gLg0v5hOg6T
XDvaNvr0222aXXnPNfDLTNZoIe0cXgT3F5devsDL5ZkNuj7jTmLvXQ6wrzgKT7hDONuYiCH3y9h5
Z4pN+WLRzp/Yr5jCaCGXN6cSfJEwJj2+S5p1nxLsXW//isvzLDqArMGh9JX0/t/1MHUGdUOQ+hlI
FtM3fz4SLOTan6pyFu//hoXMxg2S68nEldS31Z06WmwdXNyWZpoJXAYxEvEa6CUw6HJZif42Fq5v
Vvt6K+4lbOD/6ymkIeu1KRRzKbqZ6cWu9/1mAy7/jJwtJ70o/TtNKqTgQLNNDIvOhx0vcX7NVeqx
h5SjIn4pGRAh3Eoi27HaEyQf5NXUdfU7aBxmTbvkvhFU52zQN4617jd/hXY1H8750+WtDvJBPcPx
WQzOt/BQSNjFbUXSgGUR3w8Fu0wiGm3GDws6Ol0MTWA5ziNNhNGErhKD6+UmNxlaBivS7CiohhDC
19YMDKxl3e9Gma4E+tUN0mTbJOyj0KnjYdw8Cj+6N9g6YHcsOi1sQWXg1ERfy9v0YYl9qJchO0k8
SD8Xbb1LEQMU3JA3csljo94UL0HRrzol/ZJ5w2evtMujFO5o5PhdluKULFdTxX9GcQJhhG71CTZW
USlvSEX3rO6hrp1ZNLR5G4zxHYXhxdNx3Y5//JkZLrczDkPOkk6DEmhPg21yyLIs7x9cC3W6lo/r
pritX0iCvv2IGYUtZurbsmNFd9Us3uRwd04I7UVfi+a5pCazZUpgixaPnZO+IokCwAEVGjnbqRQI
4SkA8sv9cttSonSzF9NjIS0SOl9U9EWzUtWfXpxwDjRS7sXbTCJ3EBHkfQsguEM8nEjH8ayV53pG
uLgIqN13pKE0jCwpzZuquNzV191yUamXiMPP0VAB1dgr97m6VmcGW+MBvvhLVaXG8WpVDiBxWg+o
UTOZF2IJouc6FVQZT0N1bz3q1WwP7s5+CRoxBIqyEOT0qQNqlCpKQjv9eRfHxuOG+HDvqC1NVrqM
k1BeqB4LmTuKbvjpLWK8QIG+kMs15BGo+aYSM0WNDkfVta9fzumKwJ82Du66xWWfFm34Ly3i2HOH
pIMj7yMN7Izpq/fEbovYRkMEigBtvnrtgfOEbRvXrry/2EQMTlKnlFH5rJRkqHHGsb8XWp0o49my
088r2YxnMTXUeTtf2sgz55SVcL4dNlxeieEe5xWwfx0GoiGCLDyKqEiAsTrXTVlB+OTWZ17Q08Cj
EHUD9Fevq+lRBMHqbf/SgDJ/emwsMfHn/2xFvleTBAuYBuyANCsqbR0vIEqaydW2D5SkO6tnapZi
tHY+fuxxe9qdOMi7yKND3XTfGqJH6LNAv25gwIu4WIfbC9F/DB7wypp7HYFh7ZlT/t0bgRu37vfi
F7hXJBFJUdSc7lbADFMrk484e43h+Wb7rbnc0wP191qNcQ/7lnkRkWfWxg4EWR5bXpLOt5xVn2Dr
wtSNv0NXYhSYh2logkWDrLxT1FX3nW8ph0eLByGzgvQ7ww+F0DCJn1wEQ4/pFn6L9WHcmHOtBnQF
EojIiGRU6ms4bDqAquq2y++5QEWdxU6TSKBMh4KGUdp7Z9fU48GVdc3yJF2LfFHdrOp5oRYyFJHU
qmfH7cMERYNAwiKQenwJy+YyYS5D/D9ZHWStfMOFGR74fLUfL9UenO6DkexfdRc3lf6c0IGIUO9a
pybI8WmKPzwcENwkEGqw+a9VKLa0tigSAzWLeFw11lROse6AQBpAnvP/0lx6YPMXsmy1ycYL7y89
uGDYC5dQaH4s1bFPEtBG9OvYfuC6tt9AYUCmF3Ll9KCSSWQcF/ULm+Z8x6axzzzMNS1tRzYRKdT7
fvVI2J8QIGciqvgRE0olW8PqCdsv0sfLzkOlLL+SnTHrCShOhJX01GJBIxTOauC1M0DORW617SLv
Cg5o/otfxjgNdl3mF6ZVM2S9QSSvbDawy4UdWmstzE2YDejM7k8rq4X3qmf3YijH0j/Yv2JLBvB7
KBnd7Qnhc4CBfl2g8m28d5RTJDn96IMPT6E+pAoYsjLFFk+auQAjnH36TSjzY5t4FHi7YKCpIaTb
OS4WBW/uO5BJafKjO6853d7kRvjdAjT5ixGlxSb6/Ioe4Zv4/TmzFwYckhEQGBDa3oY9nIN2Pgw9
WlVyloZbFtkUNNPcpxkEi9G7UfOWHnHSRaD2uNeFATpMM+BXOAM8simrwpdjX/okqlRezy+XXT+N
G3kdqCPh5yGJm4bzbYR1ZIHf0hGVDZ2SU6TZiMLLCLbyE4pvTpBhYhqVLjlFemnrymXcsvlkcfjk
mwTOxU2PPKXrLZDyxER4TrpTMWa2hRLfagRye+Zqon1dp6EyOsto83H/EIQyDjLdBql2fhrOFIcM
v/qXcZhJarCyHXPLAW/IvZbAm0djiUd7TyW7Nfu1WKaTtrmFg8lIoEJANCtGK+a83q17XKyprp8E
iZj1kY9DtMvXs68/dcQ94EMoSWAPzBaMbDVd5OX4eePbMl2bEXItbIDQUf/H3IMQ6YlnSD1xVJ+s
UWPXqLThE18hTIQWiEK/zxo2/slLk8vdgqlK0KhLdNhbc0DKlQ9Gn1eenfX34zIjltotzO627aOn
9Pa6bxpvokw5096hecvvOGDaqlzc8NzVw1J956y9Xd90/1mHEsgv+GW7fudiC8U7K0EuxqkCi/Lg
Kbb2HIA3o7SSCZVNujyeu8gO91VZ9HWKM8TmXf+F4HDoH3KPap9r5rBCesXolYKYYeUTeKxuvQbk
UEMQS1OwjutTTMmtBiExRwnzK4YhLgAi719hQ3/kDaEDct/didyHigNWrCZp9kx+rE+e0QtNt4Sz
/l+/cfb3yysVMMNblmoSa5xBcUrpTVw1CMPfYhZUS5S6zxrYPgM0mH0N//l2WhRQcfuqp2ZgZkWS
trtItDDP9OGVhVzSU7UmjbIYsOvZjk25RVLxo+NhGLjFXZhKKtmV85ZxhpOIYVSUu9Fjol0+5ZkS
LrBa9lBTd4ky88KYfZAFlOvoDiZfx8uL0cTRDUAEAvqKtz2yzv6YnjmA77fMYehM1zaA5iewoU7o
wKZ6f6nmjW3G7wZKZ8ndwvDJ/S9SPnKIZDuaeJ2fBLaGWcgtS7u9e+7AlT8L/YEUk4/265g4jy/p
Va+oG2PI7e9L+SjMTIu7kBobc+pCQay/69+TCr6LQ/7J0QSiZZHINa+fb7Y9ZL3CNi+FDqtfxvC/
DVtAVo/5dgJSI9PPKKDL/wt0TtV0E/QhpxPGyg/pL8vrcJzt0FA6zTI2aV6/5OYfGESuBOyvOPtI
iDEtiw6upnNLUDHKgLdAuVrZMULr6EVjmh0SNwEHSZV/dd3+6AWynke11M99Bs3z+P+cxmnu4xAK
6i4Y/7utoVOxClL5u0BqO4rjdRybFtTh39LSzArOVtvo4y5k17PtAUgaIkgleoBjP+YlfvgxonVB
6Txva4g1rwehElJPO7DXsZTVRtmcLOeyFZ1BoSKi4H1wseTP6lRaj55RWOqE30CxLlFr92aUosOg
afRw3MHTc8ZoEbcRo8HvpMDavh/zP53k9YCv1i3dMhYrxeMW7goEhz/oyeU6/Xj4nrEs4wxyWxLg
FhMbAKi5kbNhU6iHLkvVMZrzv7E0D/W3br3uPcq9/ur+fmT42rwN+LTm4TuYKWweigkhq1+yeG+i
DgPlU+jEzeTXRi6JtaMSpeevj4qUoarwmJJZruFKZKH9tDi3ixDVx7MRMdn86+vijS0tij3VNwx8
tRr2/bbLlZOXGqoz50Z6pzkZmIGEoWQX25lS+itCoZLqUovNyObCaTA7qZ/k2IRsB7T1APIWtC5Y
Q1d9YTQC9EjhE5w0Uysataa9XIevohB0JrXV/zDQPl3oQVJv1OhlNgrqKNYFGbMJwHB7wakAai1+
NtVVpsjRue61TW2xN6H3oly4oz/bX4tLieMkA4yUhBPd0xpdQmiOMZVnyZJ5XY8vodCQaKXdAgno
DRVs3dJuWvjoIfMd6FT12/XV7P39e5po6O0Ok+1ENcCqbZkgPVSnC4z9/yltcP1IMHM3s2VfCWnv
WUCCZjtgHuwP7gjHDpGJ2hHeU236ul3sAPAxaaXqjFf06YFCMKS5oHmjHgwuGWOc9t457x+ux3r8
fNLlvq0lK1GlCx+WuO0XOrZxNCbLVaqmfB/0UrhsiS2pDnjprP7lXvTIy/HwN451m4CJy9l+bYUU
CnHPf41O4gXTTy5vOcN2FCnBc71n+/yZDo+VcdCtbWOlQeNT9dKV5yw4idRcGxrclnEzyvlgpMnn
/OYJ/88rHfj5uFF+xmhd6dCSevjRP5Ih87LqJsQD2r5wf9+iX/RhgmaDfsvWvYDO/pWoxHVuzCl9
cSq4FX0Bxtq/png8jaT7DLA9fONdLW5yD3VJo7BbpNiyH64FcaumaIXMAJqwsyCWBGcqVpYA95Uk
k0oIUB5W/Ng49CMuwdnazWBxSp7Cvc8DfVAOPc3e30Qfj2GW+7iQHvSBKC3JDMhVGOYzoltm9+3u
LWym/DGbHCOS6xpAlxycbjB+a/f803YmbDQsVgWq9xNWndZBKzeSp9OLEIOgexJL+WTFOTtzBf2n
HKgtavRPYXTFjf+dIvSbIc12l+dzD5p70UUFNUU3PBVQ74yL9gSX4mk3fTDDDq0ykLUgHFVAYI5J
jbxTDAxw3kIKWjkkMUUMVQER5JIjx9zRHmyECKsktKjvV79uqFm41qmXPvFb7CLdFpo+xx1Qz2sF
XnOuQjCoD70z2+n540mshcg8j089rgZak3oZcsLX7yQOXKX3/QI/pmviAzqJ8vuIfNnFLVqifj9y
bAFkr7FtaLJtWNDuhjOmVNAavDKY5GUrBCQqLYq+PKWA0nM1weUwxc5gNnQ72gcpafRYS6gu8HWS
kWE16hmiZtukpgZ3dnM8JaChZEm5/RzMqP/4nj6iClsKZiIWI8+4acn1Iw87sSl/ua+WCpU0QA9L
nSMK63yfwdsl/VJflVyStU97C5ggqNuy7dhMlo9ElMwNR9PUQUmCfo1Jf/tQ2OFSCti+A85a7hX0
eRTtL9GiI027daprlXaqlWREYL3raiKLGMtcH+A//pubdiR4b1xwZH+7ExFQIl0CTMIGwSIrBHNX
q7GCbxoymjnmUmaSEent6kEu1P//5V7uihFv2LDbIw+/dqmSUNDPiNRQGACG0nUgpc9V2kP9ZyMa
l36v6Xy4iBzLPCs1EbqIqVMZpNei5dUsK39j5h66BbWNWj2vsOrr2wq7UJcpUxIoad4DKecyTbDy
TtbQaLMNjBIDUtPihS31Z1Ng9L6MgTv3SJ8TeqEAhVDZvF8p65jkZ0/4gaYuPFKg1xyyHoaLYPoO
rofZr8ef9VGVFP5EazY/GV9yY3vRwmvRQWLaI7KScihYtMCAZvQbLBsK04pFaSJpptUkvqLH7fQ5
4E+k5S+EcFTkD4RmxrnbLlVgMmiq0M8MddBQFfBfFq3S/mSsOf37B/fOS/0UH8WGhkGZgRurC227
xDNYSNtIeZAQ4TF/3d7CRrzW43qADPbWlaxPT0SQ0SP5nRmZamDvSyhi6dE5nPHHCjGp/vtx/F4W
RR2dpKqeF0Al0NSvf1rGhVBnmhbPO+RPABbJnChlmzLm95CISanhinwUoj2zaOdnSd2LhPVUrK9s
oOxiqBAvlBacWhtIpcUuHgAnqP0jD2pWzKaUlWYpco5KIZ8z7Tf8+VSkPMCzMCBoU+cMT6vHnFfV
MkvAdAV7+Piu5C73ExGqXd/N8KmPZQb2fj7JUtkgNP09xWvjsnhv0Gc2qo1Xypqh0MrgVlrgmt4A
VQ0gku/2OHyeWDFmahoMhzpJ+IKFibnC3JtETqPs7BvlEt4jeky9iN58q8sQprg5eT/1yxodhrL3
Ib/g0uU8mMgPdt3OchPb5gyuqWsIJ3BGoACEfR5Rf6tEEmmSBKa5SlZKdFqxnD0/ObUG3pNSRowA
DzpCWIWW/1W4zdyb1sEPYt4YUEZv9iAJ9Abo3EKUNjFSCbP/Zx1MqUxC1JJCHWvAjXJUizO4E29p
ZYljrLHlox0D0Rb00YCIr7XK9qPbZ1H39KYYcphvKbSuTohYsgy+CvwvVrMih4E8rUOPz/5/4lbd
vAeaXXQieE4klwRPohCi3L64jFwC1FH08rONqP+/0LnWxezIS+U70Oovbd5CqLaEHx3/qopinX6I
8CY4Vx7US9OZ7sCtL6FDMXU5lz5iiW0U4kQYai1vvLgW6cryGVW9xXpcDazwrMMqVLZmogo+ZMgf
p7ztWhJdws903sNLJUkXvAUsL+4VoFEfAXHzSUah23tk0vo7no1Guuye/6BZtueNHxD2mheBip1P
cN2beTfuWbOl6sIkgfKOv5V6N4PBy7l0/u8NKU8LLY5uCXI9AhhjFsAeGn8YZAarl6ir1V8bWkXL
PvyggU+S4uXWmNggyrXyWff84ksMbrcoU2T/0nOxmyEW4iwv88iZSVd2iVzUH/+I14jsTJfOioF6
710sKPEp0YlW2jXk33oF9uZmFuMKQS8JcYyiLmOuRTXovToq6KHcv0ZWVMKL7tZoKqJQIca3LqKX
a2gbOuBYCrpoEcKqFG/rL/u79y7jxICyJqV7135LhkYYtjFKjKHtVG3fxBOb88u++EWs1OF7+faH
qgSLwUnY8bdqP3SslISptJ5TkIxdBe/K1ilpEygK3fQqaLQU7x+KDffXNQVguDE8JFmXOh0i5u5e
47yo8Ui7V9u/b5vUfdd/FzSHdUMS7V6xLIQLG2kDGivL3aHKxXa5rNVEwFnz5fKmH9gA8NBfPTFo
giGxQFgMR7ZeB25c65SwfqqKRPfycQ15pVwmRAqoilEe2mGs/wUuQ1smpgmAKv4RV85Kz4mX7mFz
q/jdLlCZXC1qiXl7xn23MtNLSzVjAohfqZTbJopnS+spuvF3nM6QJmkdj1HfN0Nj0zrFji3nFcen
+ZiKgOGZQADF5HaZeJ1apv/0230vz3d2fG6GpPf5vHjDLDwmd9/wqOr9akWL1t8TRCvehCSsxDTc
UWw8JDizvnr4DL8gvSWA5UI0JS60tOoq+D1FsvrPXMyP1YinryQ2bDBLLZ3833zpE1h6IuXRgWj/
0VHuHBPc+VnYOslasLb5te6vLg3sGglr1nRVMIjDERvlaLrdmEvSEmFbA7pOEhkgisePNMGNFgYF
61jyCuEFQ5/1Mrv6JeDv2m6iDxK+MmNNRXF3JT7NCfcXPlsAQDpfz8DDD3+S9zRv06c4YOLQDux5
IqOOGTbR4GHTtY8cBcne5nGARt77dqPcD+swBmaSbdAfkHnjehCZ1PHR7YT4DqmKnmb+erbUcdH5
jiOgUFI4tidZsZ1LD4zf7MMsq1lfWw8954xgTnfZoZ0oZBArz8e+r1b40eW0OaCoyZEp9XANGs/G
jSN1YnfXmi+vluIFTIp6og8RtbAfxjK4CWOoLbix2fiJ7EIC9ln9ghRSl+JGJQjqp+2suphMrO+E
wG4dGD5QEKCYEQ9F0Kvt4EoC1Y5ZzZg6RAP9KB/jePCsurmv+A5Xz0/zVsTxHQpSNSr0cdSKaSCZ
VXuXY2Ncd+Y5/jqsPXbuGapkxiI4943VvdVuPoV6ZhlLrK3ffI8rtsbZDjCllupUHLmV4JAA2chD
kxuosIR52DERhjUXD77scyFQkCTBhhwOjWfk+NcTW/yI/ff6KXI3vVQmR+6AHAbyCB4Wz4bx5eA7
Oa9zTBb5vtDHBKbYJqvCLoMQGge6dYp08XDCxV4J6uCQtN2Iru/OOdxhJ0B0W+EuWoSkfzT/6/4u
ekg/Vq6DGlHY+LznftpZ3QtiC8ahsSlHwtYAwCadsxNMPIMfXRZuNU77SXYPo2aN/BLHI0smymgf
MWMbRezYA4P+5w+/tmPiW400FhmClo64fmrA489qCGASFSgoMQeDDQR9rGNdpLna8w1RC8xcyIoR
xaeDZszSt32SJzzvTRtseQtOTbmi2kzH/gj79S58hTSt2JbXSPwQTCMp0Tv3UJBrCGhIt3yLCge4
uEM0df4Fn5JqCvzRAay3kjsu0+6fAtjEVnmn204vKUOqN+KZdZ55XDSFWD3FrD4YBm4zn4xCitCG
Ts/Bh7B66iDArwCBkOEtAlTLi/ibfCxz+CRtzeSa7ocLMS5QlIZ2i1+QJ3bGh4boZE+GVsV/uPKS
X99OjTXiaXRGKBgswH/yc8vIYRlAioondCQA2cQMZEsJQXr34v5555hbhDX1thM4EZ7Yuo3YDces
zf3Dx9M6eSQk0Ne50k5ti2GKymFwxjrZ2En5HCCc550OMTUwW4S7pO8d5s8pnT+PaUTB/ZgJbV+O
5CbMILhnv6THQD1s7hSFFSiBqSqArbcbcXfnVFzvQdSKx2/0at3+HVdZcmfVRVQt4Ta7f4zF4H2X
mYgcHOpn8B2eDuXkci8djfDnumJfBBPo1HNFsaE1Ymz3XKdveFcVJK6Qe58H6U1HS09YJfnnaXmL
ks5K/rW+SjT/9CQua2xtCE7jEOhiq5MqojoYskFPLcK8tVo+G/99T2RphCVscr9/ZcsBIHHeFJNp
BqZKCPOVdbwAgmS9ULEIDnOiAbJ8jovYLqXOilBxtOrLRrOGW9ipEdbEzlxJVYcubeXpf+2q35Hv
aGuLwMY57Nra73QVX28WMA68LSrczHOxCaVgRhC2ZVa1+j3h/pwkdfE++E+vxpf2uNqPe2dGoAE5
u2HYJt1paVJOKbM2B1oUs1vC4V8VedmHIdOuQcVqj33+7lArugFm5GU1ozUDkXh1rMPzcXQCPCjw
fQaGwvTLtF2JxlsBxlvHBdyfqZvP6w9mfl1dXcHLxZ7W+u/L0gBTMc4U/KOCuwgMluOEWIPgbfOP
mQCcVGd46Nhcsnt2874cC8SG8cxC316Unb470C8O5P9QTVBP1JbV9u2b1Jz7wn/8PwyaFnY8+r4d
EeHqkutWRC8kC9rF7+Qbazx1y84q1Mx0/us6JZnmzv4AqmYVRIutLYp4w4WL1vhERmcqcT4D4TUy
ZnBmoMogbx+SD+3QvzfdeBSNzPYabe7YzUu74pILrxUMqeuQFq4QvWfT4WGCWrGQmt+MdI49oPS1
FOQk7YWeoFD8j17lXs2jgaI0ZqB/VMyd/bwXuJF9XqrqLyBtjTGihK+0wztIw/Jf9doexQJmmZfs
as/QHWFooFpocO6S1Ob7elrY1xsyRCCcIwvIRPd3O5c6C++CKvckAPKjrv9v7evx0i49SUOQ9wux
y2Wby4o2zbMPa5LsC3+LSQ4JvNDA6NBLF91l8Z7Ru30cBlm3WWL1foxDAZr912G/5XJwXfcXSN+7
c2qO8f5/Z1zde7HbHpwdKVAGEu47X6SbAHJqSqo/kuMVWYPS1sVSJ+AV7G/8ZY+Net08PR5ecG2v
J4ZBDseTnMoW3yRGf2QQVZcgK3ISJvTsAGkvexQe2cmuAH/oReiJhRTYsFxicxol0hO1R6DXZ90A
zSgpgrYRwIiYEtz9CMzS7DuvxD/lHirfp/0xSY/w6V0++KUJ0BH5h482SunEO0mv+iFWd6Ta1XBu
p8BwewuMkB6jZakyhQ3Z642w0yyTQzsOtwyB8fQHETe6EnH068YTD+5qV8GGnsmZEUiHaI53TNB/
46VsYoXNScYtodbebvv4nhhL8ItL1zjh72dVO+8RjolNT99fzHeqaMkyxoZGoWpPsVar0oDLKwR4
Cq09eNbDrTAYy1MPcDDZsSP7s4FZofiM1BV2nE+v6iXltWNhiKoYrQZn/6t1BmKYzyEVyNR4Xtpy
VHy+BwowdNM43dYQZUOO92pVSHpFur6yE1gTe4WnUoHeIOlubv8ZhWX6bb+I7yKjYQRJP7T9wp8w
0mC8OrsoNYLiZ2jsQEJbw0KKs6aXSSL5uDtPaombkaZzD6DhwOuCIg4I7C9PGgr8xdvpSVQBZ7k5
HZ/DAKsAKNVDyrJ1xdMuuYmMkONeJfELD8x3ufffMiMFt7nit+LugXh6rg/8aGinsaDriDEwBQaD
JdmdM/sC16dt2HY+X5QODkg+TxSiFsfgtrK/4yQrCeYbR2Rsy6RO+jVy6uB14W18dSHzcdHP/uSw
R1EQNPxPcF/cZ9e+uXLY35F2yW0ezgKUYSvVh94o3fuZfChmPy6eTZtmGCP/nmDO66Zu1GB9HXqx
W2x3CagjfdfbNvCttoOiOqsdU/Uw+8Sp9KluJTDCQPHiJiytybu5qs24MMBWbRzgoiWaZl4N8Yh/
FHf/VV1LzLiaNPVC+r8LrhhiYVEMf1LkvAtu9WOStq8DldkbrtVKzzQTRycimu1sv3NggUJNswkE
K9+4OGiX/KglDKKRNBXSY13ASMaszAj/3fV+I7DBwf9gRR6QoF49IYo1MCjc74UKMmogphuBgioL
DEMJUpXq/fBm+3Smmmgmj9GgmKpoaUQCc4fuIh1Z2/jFdRgU0FAmKvRmjlPI+FIHPWJ7D1ozHpeS
V0fJLiqARUOQA1lM0riJpkQUYT9oA9E3p6NHB8MfgzN9bEUhQcJXmF6mUCXFkyXMxmNlF5ufG9E+
hQp/aH/4qq7dVY9BFBBopT4cfWdW6nemkm0IZG7r5Bv4DKjSn6N/iNT8lVt/ERarn+XBws7uqt5Y
fIB8CKfh7xl03Gu7xL6YsGPoG8LiYbxk4w/MQsomJj5JRWvUI9nhb/8v8jzFq8uyGcXHnmUurvXd
X66SmyQBZWDC5of+wjAKGsZgmvgey2v0T6R4MmbeIJ2c+oZ1wJ7bqPitL16G8/l83y3H957J9oOh
VOG9YtY/Plr2RjuOQoSd7ERGRtke0hAwaLx8GQSqjxFIhU1ItQoPTS4CGAgn04v1aRPKOeADkTzW
TtHVqt2+IBSz/PPIhDCR12/0m4L398mBgnvnxHBnm7fUQpUQ4SCcm1RsjRf5+NRf7VSKwFZiofCF
azdgsqLluKY6EsrTLiOk6BKs1qpDTS4tT0WzPSUJ1kBT73ODZnIoYdw+B0r+e5fxQeVKyW+oZQ1L
ldMW5q9eyeXI0f1nfd75gCwCFYyAUMHjnYemL5P+DZ8Q7YIiUZ3DxPo7E/UCD/cXk8uTkIPw8nAs
Yj9TQEsKJUWaijkV2YGspHLpTxJifHwFDfxYCFNd/Scqy4oZVWk07/uTgudEHayqqTqy1al3ENN8
RpbNtmpl5GdGaEydMlzvQBFDWjixO8MvsQWOehurspGf7lJDPJbZowxaWwigBrbvEnm5adE5vqk0
RxErOibRw4Vt7triytueEjgcGjiSGUrueku5c92JL9QXZYI6yuJV1nLcDt5UQnUO51X96HJvRIym
hP/a0C78RxYQbJ7+4yHb2FrOeIF9YXqL5nF9rBXbEZvyEDnkjdr4TiVsR/xVzUJg1Um/F7lRv7Io
SDmnXauHBXbJFzTloYeXhBnNclmjIfiztcMlTd6FPND5YKwzt7iqXsxZ/SOfeSTuYletUEROYoWt
da25SHNmPTwCkROBCBnKHlt7tq6cOsaT5HzlbueKiK7e85xg6dGM32SclsSx1PoxD2+hIxv3bP1L
21V8cP7omAuff0Rt/E4L2KdqnGqkymY9H25iHo0ngv/wzWf3xF0JqNKhHQx/PKTQ0QvBbBDg0aV2
kYMTxoemUsDMiOPFYSkMGxTzxHR4caNA1Ugd8xgDAWlohjodkqXfQdFrFEGcdGG56NQms/SzR8VL
ptdFN4OeV1n87DcPAOaX7wlWjAk4rd5NqbIGBqy7jX486wgBbCTM9xL54Vf2Y9oRoifzAz7ar0oM
EvbDVuA0eVbus7zJl0UBgcHg/lBhiNGjX6IkWCSELT0ncLDC1z9kDHhwX7fNDsIe60jYSm5Nkc4x
Wjor4cHJsgedG/EzoUgYzKMESvOlfiFRTPb18XMQBwZFE2WkdWO9Hg+Cj0m3XCJpzkprnwRTnfK+
TZ6nE9NCQNyYy8g0MsPBZHRh9qy118Na+PIz4m7qYzI+RjI56xJIrYLFp2C6H7J21iPiwAmcjOF6
ogSFVNUTlN0nm5la9eVpvVk4ygS28KoOit+T1cs2mLgyJ26csX2A/KyW8eV4tqqQu1AO1lkaD7VF
Z97L6bSve0jRj1r/KkLav6isBgHicGn1kOh+uzYBdcrYK9zvCKtpfN/RtAczs+eHpAxESwSthqz3
R40mdNVskxnXq4utKi4r4xFcijtA8CaZ2NylmfDpWBYRu2Nj5crEeg2ZgkC5UOdv3t5X8gkK7Ox9
rRKGI2+GME5JyYuy07H0VCVayB0Vm6wckZLs2NkAkh6aXdoQnKVFMyZDrGCBLhTkRxenvg936c8R
33q82aPwq+YCzRRwmcGZhRMoGYCrAkrOexx6YsUMQKD/gUfBTW2q0i7EDA2iixG9FN2Dkua/6cLW
D70tj54+FcM9GqG7SgdCBTl5nsOim2w/KahbBY0iU/TJkver8W6rIsxr74IEUOVkxe9yMBJRMEn1
ooDJs/FYnvkdzuQQGFPkoQz6vDlvMC6GozG6Pl4+Vlvw5EPtZqEli7p3EJHihVxsnj+xruzlF/3S
x/5ii85SJAPgRoIhfFR5eeI1AtgpfeMKXWIe5iMypWLNdXb9DxeGh8GLAkwtDVRl9W3M8HEQSXbZ
/eb2q5Pr2Klsr2ZbYvbYbMmbbYtW0aSOQ9OO8jjDdqJVhrlb4uvO2dAbIyHeudEDwPce7RmL444X
Z6sEVQFM3vchuFvnkIV9whzymITP2jSggb8rcTJr0TTz7FRSXuFH9DCQJktRIxa5dA5xnhL86Hax
fNkUxqkU1h22dGrgHiZcPOgVA68infMKqaEaguswWSkQI11dxFw/aaD69vwQCwghVMiKJjuurKFp
4rbAGmYpuxdkm9hoD6RVHlJhlwoef4DnoHQZtYPU4akLBjmyeXUFLio7Yr1IqmETGxh1OdPkPHeO
eC01ijxkIOlIIeJVLuntnc0TNprd7hDwh4pEIj/ehGfvwqUgCGRIx/XZ7UjX7gFBLkyuEOxvh0xy
eUBVs0/UrJKCnn/n7JRHxnMdjFnnZQD5oHcwB0LYAkZVa0LpZWUIUKxNfXCvxTs3Y+dKdpc0LTX4
H41Ws3x/5slErHPwUan/S90IQN5v4J9Qy3sR0sVJBe5QUQtlVFLUbyrk1ak6aGmDBKTg7qgPcVIX
PlgGaYcvbC/dkJmX73Kh+v9I6dlXYJ2cQYTS/I33e3iv3CyjvSzYoKhYwANk9BpGZr647PShF4ah
8CX+flm2i2FVX9dxH4JqI0oD0J/rVH+1Lr62+qGi4vGsF4/uyZdwGZ74BkNfwPkheE0xnbDrjoQ8
+Q9bEYm6UE1MEyZWZRMHZxxtX7LB7LOkm4edj1nkMfrssukh4IYSafA1j+N175jQLV+vDdTKHxrm
aP63ZW/9is1YTtedDiT18uj6KpR0Mjg9b8JFvzuKSKMAqAFgEY8W9ycDoiJGyoJoemtX4EGRXCD4
UO8ljkwCzzV5pxB9mRIumwdEOu6XbDRNV1/2IdQFxbguj/pupif9NfGQS+TQqefoOhuCnKeeL1ft
zDZbWGQE+g1U5rwJnK2eTbK/7ST7ynR5hWMq9EdC2BB/RgrdAPuNZ6LUtuacmuYojWcZtZwqPQTg
Mcbr27E9t5oQJKoI+eaG9g3BlEaB+XArb/x8pCkf7s6N7O07TgV/bcfmGEFov6mi8QdP43tZQ66z
f2JrV3NzGKeBTHBEX9vHGwpDsi4ecTBQMyL3GByWhI18G8tvFasfNKCUb8RLq5B4vq8Onu28ljwT
iz9oOz3/xMqH+dv2cuC6IRjvgZebaDkqmKZLonjdnjIeQHKZDLDaFr+0tzFZAc4LVYHy/CrkKlNJ
Y2dxHdpn5cb4nzoaXF7DRcc1/d2ILLrRsmEFJjTb6Mhw4dfKXf+W6pvHed7lr6oQrEMJrumNKdZM
P9pleSwB7m3/PBTWM1gllB66Dg3kTPcmBOP3Lq2xB7ZVGJjzdkRCLxeY+EiIBCGQAaipFamEzJ7B
BVDf+PRJVEbViILkipvapkx5wpp2wfjaQE03dcoWsduUykUnNl6bVxB+G2Dx5t02d7hgYMKdLDT2
QLX39xnNv4o4BeQAD6rv7W8QBmet+XTuVGsaJwAE+SNgdSHhTaCPK1O+5qdCfF90rX+IZJhZjtAm
Yt0tCC2hCGby5C8/01SmmaYrmobTXym0o3M6GysUzfYTztDMu85h0L7+taRbduKOSLk/KYO+tdVE
SSctslIAQ2YWJ4zk6mDVWjwM40mvBPWnWOxKRCNRB/UzoUB0fCIdILEls+yVkRg/AnlUkJnCVUyO
dmeFQUyS3/OXxs/rkTJ9/LbM5A5xsLkIyjUKBLPpBvHEMU3owziopiH2cL7op2BCpR2eMYwXO2Bs
cZt+yoDLUce1jXIpwDsqUIcM9lRIY4Of5zkRc3LjHapj+3uT7x8mgSdvCd708VVh+Sm/zMX7v8BI
2ncXq4clNvyNKUw72fE+Ts4Pvz6klruyD2yGI0qYVmVVFnahnVyQ2n/02eEuYglvEjRZXUsznZ7q
XaBmkmjRDf+Y0ff6g8Ky2RQ3g61gDfNioGuzz5HyINTZbzaMGKIeLtN3gScgOCM2pxU4dHOM3aLF
h4LMpG0N8HsMxGqDB1Ul2LqviKeOMxtwmVCcRbxhYmlM749NKY61jEl886uZ9I1m5fBx3S9Z6pji
l+lIgMBOhhnqPA1Vlo7yQB1+nSfuQ+KL3O/Fdv3j+f/caYBJbosByKEX2yVdvvSyjrOc3g1IJx6a
J2NfEzNQT7a71CbEdW7RULlSa6jV7jnixzdcH8uEwrQgkBuz3qgMH8X9B/xFmZnwMtFIpmCrF3be
wlJfbVwMz86p2HehI4/M3SiDEDnI2JRUJBxRumrb2h+kHZLP9RzCzifgHw5yGKaZZ+8KZtW3CCWR
FHwaC8UXPNm04+y8nQKV4zXXbsFQ6hA+XDhiFuEq6bwBnppsQqN4R+ugXN56ZarIdJVBnj2PJZUb
R/sgLfh6GbPYyzzYfXy70TloArEo0ZNwYsnpd6roMjZ2OJ0j7bpOKsfjpdVurZQ9Ue4XLphavp7q
vg9qWDy/CKOnJJgt0ojr+xmh3JViCnycNrrVpKOn5V74uKbwbVZsFq+CGHcjywdVATaoI+62rGOR
PYGKfZMrxCW04QxMKdhT5joyyJ1HqB2VA4M9QVsDrT5C1HoICOY06kkt+5TmM4Ptg+rMdxSeaKjI
s01vinXGp+AaDvPXqjWZpArBuvsPP83vz6Tm7BWwnBxFnI3KAEk4zwUXnlXvuwa3EYTgZFLJCdkI
1/0VMKSOdqVnxOHHaCwyPqDG5zs4qtOjAC5aFdaNQXUpvX33Ek+uxHs01rBMltbeotxQPvisfxCW
G7SbpMD8fBzN+5LeU6TaxJGlt2crp2kgtx8cN2OXDbRnGOiOcJNDcyQQFHfnAYQdjr/c00zOzI6/
l8w7nsvyTRtO1/zhX638ZeXFdCkfSMtZ/Mlq5KCrL+lheCv6L0h9H2iO3sj2VhU9CwBs6qfU7LGZ
mlxz67mm6JARfdyW8is36cPGSS5v26KNMMhwNZVbFeRjeBaAbpkuT7xnk121l64P55qUZt9ujn2O
tUfPHyuFawaPhrmNEJud50TuPpPnBq/8a96rPImfmH7K3v5qe2WrJILoEB+d3/eZ58zX9nTw7DFX
Azjf0FzmD1MJLsJOxI8HYReBxzrkFIsBNS3+pLloAf6GzPyVQ+A6TJ3hofkkPblKSrsZ/1KdEsWV
CGZZpKcDKOm0FpphyNa5NBBkLaf+JSP4tbKdmrd3JS7dzlS+IFGCKrBnA2KwLnxU8gz20xQvDvqt
sA7YtjzTXf+g6KzWSAckmqnVZ4K+bbLk1REXL7DofhDwmS2qUgrT5BbTfWPcPoFBAkIzXI9Xd2oI
hCtFwcMhP0FjjoAqbKBh7FSqEBPaDQ/SaahhOWBGwVAnbeuOlDbHXicSinINbo6rBjNiC4vTi0B0
FVwMBOe/SYGXnoDivNYGNhQnxjRKY+mrjq4FBdi9E2nj8EgiFfBh76judtYyE9TL/ZpvL7hggJBV
ugxGKA0p+ubr5iD9dpveJ9/0YhocqWDVnzLabmvgwW6Zh2q6LUM7sBlTpWmW2/fgXzJzHBaglEq7
waw/3ZCV4QEkV6bL5dFbX9H6nH4SINts0w/kufIP03iFpygzkh6YZz/IjhAjBRd//O6QX4Ngtop6
KXynALdDn8dUNw2Ng4KqcgOuRXnmTWI0mLwd5Hw1VigG7qCtWnc3PNIYTAKsh2Hrkxf9mMddKmGv
v6m3t+0YYoWyau1dAudbL4b2Zr2TiRAjkZcKStz3fIbDAHgj7vGvxBeZ7h79icdvIKVIMZBqunay
awL31AtDxN+mdoajKouV3VFy/rmE7FF43AKLZxNcMp9boDSI/EakQdBAJHzLdQ09iy6wOCB0Ru74
b3297kK9HT1B8g+lsGN0x7hVSg9QSaC3m3jIe4eXAoKkYbRIM64uSB6Epp3WXX/Fuc2lM2o52iE7
0yDWtklByyaY1nmYTVAGRg4V5Ku0ccMZadGbdO7gYEiqhI9HzMW0AM7DSknGZvcS+tZfEVq0XCFd
zzDQqLeGY7dnqnIr190xb85m15Pz7lIoC+T4QM/94oswoyEphCTbKu0a0TwAtIHbczjl8eIESTy6
q+T47h+e98+uMCPJzUUHMLS06xrOJCRYB9/NCKhNdKN52+rkxj7vgXFlb4LBt39TmZuZzy8XvVDU
ckIVpRr3Khb2f80/sU0hyDaw5IwtHxuZR78Js1bAgUH7LwjWnf/9AUgYqw4AbJxWXl1POkHZV4ZH
NWbGv9GuNDsdVFike5iQCXiTOVXd2WKaA4+HTG5++JhAYmphvd/FYdXt1OArSvlTt9LyQXkvV0Pe
8BlJsB5aLZdAf6pkN20uL56TstBcHXPh/0jbJ7H6Sfs3n5vyRzJWpX+mzPJqZUwXyunKf702gPm5
Rj3nyWT+nbxn7AdyZ7ssLRmOTza0IAJ6P065sCfLKxxVyu8f0jDKODlcJjOE00qwv9BMDJTpkaYM
/nXMTSMOVqxUteRRMkyr3vo6M3YCSZR5EXWuPqVxOpy87uBU0Dr1weDsHjZljTW0SDenHcGBL0V8
N4zXyOyGj6DMxbbWUKBL8inv00Ri3Y5cu7eSGiBNHmjLjjIS/80gzT+nnt3K35NCBoRaaybyXQQp
xtI23vuU/EjIEubXtWSn1/eZokrA/xmRnkTWPNdEAUMH6tUBdyzKZ6ZBeudZ1Usrb6uG65upzUd2
9521Ax2AuupcYmlC+u7YU0rNdKcY6bQZiOQOrv/ZDgAepGt+ygzgDTEwq15yUmHO7DqIaU6JACxq
8u2PROcqm6AQVEGTu4HC1VvIKLuBFHjbIF5TmdieEYLzcBSzSXkj7jYiJRWY2auiwB0/mruT9FCL
ODrGb/KKNIe4ksB+iGF9ftp11AyEXyDQSmUxAtNWoMxcrZxv8eVQwT9Cn+0yw1zIvDxnKjgcSXx2
I8kZo5+LrV9vk7aWuDLnqTvDyzdsPUI1AosocbkWyANTO44+v3eelfP1nTH7iEscBlXz99V/LFP1
K2dtatlSEsDysdWfSecP9RQjB64eRsZh4DssdYxE+en85V5QkntkUCbYaLky5UVTyFIt1gauwr1m
pLgsLUwnNML8nIJ9wo0WdmIoW0DCmeMl4oSbhIEz8vpBPbv8hOXSqKH25hmyq2lB1/gsAfHwZhWz
EF5rLcv4Xm8HNvof1nBUfLVsSF63tTCQxsUKECZU7mza9CW3w1EUp+a6l42jkyE6khFI/QdXbpQt
9ISYO7FtISWOMWlgUdQhmChF/HTMZKS2owDXDImt1G6vfYsURtlrijefHeX7dCjbZeKxOiOfS2P3
Y5DXYKMvrZw2cjtOFdhAkX+Ja3Q8o9PMpszf1ZPhC7WGUz79qVALkODgGwWTSawN3OIx9CfXq/c6
Bu5DJ1a1ZettRbJgJDApbM73ImF5pXaLATSW86AdBUk7VYt5ZHDQiTmT+vCyI8iGM2A916OHhnoO
PRwwM4O2TnB8gKp48rbFa+1ON0PlkLUBq6BG5a8QQGZCiP1q9SF+tKH3k5LprUSzqab3yJ7bVB3B
K8fGj1aDYm/zIAcI9GH7EbR1RZgUnl0mh9/fFA/hMFn+oI4ehvj+WFoRmCusJRP2iqNInquzhyTz
iF1as7VNHkeBXQaf4hD/aSy/rfSflAlBsiyloFfHnzZ7e7Ud6TothTUQ2Gp9WWaNvoiLj29TSSpv
dGAonpOO1wH6/BtS5LYpqZ2tGrEfP7Y+URD4PKBMhmH2EDEk/U079wuh+1DRpJWORLC4SYCq28AP
iBGZQ2taDJo8CGt0H384tjfX0MJ4/IHcSKlKbM3KPd4oXQ0rib2Sokydy+yynK2k9yOyUAlMeH4a
9h0A7xXJYhXkD8kG9CgOpc6leH+Qp4rDNrQW5fNArzexHVlB6M0TlKh4VMdqLnlA/LcHBOY29Wjq
Im9AzAeSNsvXis5uvkrbznJlX3h3sk7Mxio/DX6zzHKGS79QPPS98siZu0MqWpkp98z2LaeCbvdV
X2nmSEBWkUK1LF93e0OhggCePOUFru1gM9h6RbZu2SbhqH8tfqJt7mpvbxJq7m78OHIRyXhIn60n
KX3Y2lT9KeaEb5u5mM3KGUe6M+GYetLkglGqsaEgl3Z8FCMSpPIESLzfPKDONi+ehhySEC5XNB0b
JTle0hjd3DujeNgInHbVZzgLGqypA1Y3Fv4tDx2boa1m4Gcmwqk74xqub26iY86Xe+EqWE0lmtOP
UTUaPNrp/5AAlv6v3Z3xFtmCD6gQQHo3T0GcOXo903PruBvfBB5tRRlF6vF0VbNouIFjcvVcRgNc
f7fCblqeHaQq3AiHEv90koCJW6v9zIgoM1lLWx0LjKamGf63bR60kXDkb7kdOdD1k6r8/S3gcTul
P9zb07H/ptD0bP//FLFNVM6FGHuzzY4ckNZNGbhfN6SXEdLa9tv7CwdHd1+GvpFsWj/AgCE80ylQ
whNRN6Aovy07nf+HxedydLyGrDz9eznzmlLndJqPaXbNcB0uesj4wsmM46jfYvSNyU+RoNrDKltw
aFjuN7tnH6+War7BFvzbnNKPnDepJKJcMq1d3Tw6MoSb8DiJc/JQggYv+zB61KO2ZO1Ugn7NYCKI
EkIYOzn/2ZTS9SmdKQX0z82gdTMmZmATMOkhqAEoRvW0zzn8oJFUb8PSQMMMp4mHclo6wlSu896R
2LDJoWOLP3TnfEX+4COZfzb/1yeOCYbLzeJQ25Md3XtJytEYuURuocLjZZrKM7PpKOlYSjYc1aM8
rOVBfgAvf5HubObCU2Ku0pMMWGMmgCTH/SVIrqcM4jVGvGondM9EGSGstvcWFATimXIMTf7yuuZw
XKd1BKUDGST3tGSYuNdIJvj0SgM/eJFPvbaSUdvGfVQgvkOTP1/iRkjL3y5l2DXs1RPA+UDWmyqG
w3lKDe3539A5jbqCQL0bXcOuD1pGnElaV0JI8n+rx/QhTzporU4s9VoxMWY3aOd9tqHj5ZEpb5Wx
Do+Yg3Qrbq+EYnhYBFdCSoYGsUOjUrpyY05TpBo1WvPNAk4SJIbG/0/FaY8TeeZeTBBOtRxRJADw
yCJB3SWxHcULL72JCRFltyf404Yiy7KJBc6ebNdue+E1y012FVcZ02SLZwH8uIzVLkELCOqGa2ok
6SZsxqq/+d+BC2aTxcjv8YhtaSc7hSdhfII+WCC2601Fhkdt/mElbiTMxCOvcpL13MzBJ0QUDxW1
giT3GEzwuZDGoV+kKD3O180Dlu60FSyR3RIOiO5P3qyhvZG1ZqqFuR0XRW326/khdOwP1kBjW9kp
WU8asACIu2hWwL2lVr+LMHKn6W3Hz6EAJXvC15tlGCuSBCX1BJiAH826XflzmT4yHqUxPUBpTrcf
kObzLgbq2WIDOmGRyO6ZIdFfSsHHxcx23a3PzToZyKntwxggOnlDZeem8BGXpghwOHLTTcdmRyDt
+CjksqAbjJ+BNUQePTZ9d14xzGc9eftr7e/QZA5ROUXvHs4/UeTnEZvtKRzcJ6/KYpcES9Eltrct
tefCsr+di6M4AOr5A+XYOI4n1wb5utaFU+9nbYnk14JKCikM6z/TycSEjXQ1f+5fIb1oyY6KJf8j
eN2pXT91Tf1e2CswDfsQtSCuc3xPyasUBRs42SlwjmdQpiFPNwTA6IbQ5lhamjgIc09pre36PVO3
yg+P30RH8xzgvxan0kPaFG5rYnOJnfP79Q7Ak1KoDPTC1ofHCrFdgtZcLT5iERmn9EDPOhEegSZh
APQXrZ2Dozfojd5FaCFIMg9vmjPgZEVbb9yUttqFwJ0MxZ1qy2vpqA8V9dEPm5TIKvVCT2y237Z0
j5KvQe2sjy6gq2eoeFWznJxvqmTyFIvHn7bMKb5DcVVFvi9Hl7vtFYirZZbDYaV2cQHix/U+pQtc
IWVehZHuA4qfLZkLFbQy9vAY9GAa84CGmrA6sbDIqoHBQkGbiwyNLBVQOq2Ug/qtYwlTmqL4MaiN
zM2qDKP5c7m1einIdxeB7ork5aVlfJ3KI6NyY7wIc1l1/2bM9DuWWqGSUQe0QKHuDdGhIFMlKBZh
p27qwY9fFV9WeQLlFKpW8Nu7E/njsaOqyfpUh16Bc6ANW69r4WiozzC63PB4yIOEkMSLdQOkZqdI
nv7Eur1BUzGw5bgxmQQMUYt+wNkEaf09os8aSvcB5udQlyyIVpDS8cuM3XMx8CAjy2sOTHBcc8eY
oUY4xvpYt9bL+etdS7G+NbdyP92jEy+Dw8TdDVC5Urfh+8rjr9jxE/WpL1/ohJFg8EDw6Od5Xl3c
CALF2XgEbJFmlA2CCvsI0mgFJhw+DaoDXKDmwNu255bGbyAmqmZyneVe/Fsz2DzWQkWiv80JoChk
2zfI7pEsFS7++NFdhgdFnAlun9qWs0BlWYYS1mwhM2oZv1/ZthIxm8BJgbA8n1aKKqDVnpxyThsy
s6ShpqwzTaVjSevXtGcbsdhm+CfK9dlpGYXPdb7yASdAYrT1Dm9Ijcid6Tu+Y+uPOfYySAW7Pzus
quyxI+2xx/F6KvRwEiwIjYMeyfbRh80GKqDvBrL84rvYuVT3+HctXN6w6S9Fcc3mEcJtFuxSqAhG
I0MePG5dxSoVJmmdSDd9kQghNZqdVN/zwjtXRiaeVe1LpLeEq9YevtZfBDPFdLbuNXV113kKsw//
kwTBIuLp3RuuLw8Fdd0/m+Ne0/NmGdhCVaAqaOB98NWGg9F+HQ2/QqbmfL18eE/HlEzJs1KBUOcC
T+u1hZ0k2nu7AvdcGnCzBKps2EuVcWYLb/woDsFY4P5yL7bJSLcWYUUJMLyhKZsgkxmAxsGl9rPW
1SgahOoCmeKlLlTuHvTo7cDagQ5PIDv+c/SufOn/hvfrtt/dDWc1PKvSkagTN1M/yFdkvEsky/vo
/M8Ro5poQzMhsQp6bQKvrrscQw4yVXwR21a8jeyevrVU76OHydMWGDWtqPkrJiWTTJPs6uakU0XS
gPFFSV2vSqyGDlkVBOC++KMWhYZ+3RuX1m/G36rTMVELWz3lP92JLalXXz2qY63KKRCTpDI6BQmM
/MjvEnDxSSThhNy6duAdnTIbSJ+V2NeMXDdXgccDfesXyOsz2lvMch1HIe4UC2MD00wM4vkeNAB+
QVFSPzbZw/ISW5bJwp3ydufyHR3Zfc3C7RzUllN4I/4H/AwlrXITkBsVt/uFYdEBhRl2I5jxkcnf
H84qo0U8fx//I8IF5sJKcPTDSO3wx8diM9DC+IW8OcuDX0DZ8sUIH4FA9GwZqJXKFNt0CVUpQ3L/
NRIKM6K754/5dw5VyOQxVx1mYGPOaq2+5XijT6XgTIqdYW3YAaCE+Ji05dryW3JAPhwUS+nIXZI3
cf3qg78H9EwLHdTj95EP0CwjcVato8ZZ6moMjtbfUlHxEYFLEKtNLu4epvZ2Uw7Hbyifo+TU7k2N
ef8p3P7kdIIFEAEWJLEuEkZPKyj6ebvAut0xwdt4AFBoOh+W3DCkpaTHfrWBAOYt+vb2fbdjIgVS
GunGOFJ0jfhNdmjDZxU+Xb9Gqnu9+uStz10GehpxRhEBdOmDB6NvwZN6SaQBArK2aCa5cW/QYeKy
8IPKpSAPg+KSf+6lI57lR3WSJ9TGYHvEDPaUybB8esT7T8oLMuahYaUW0/9H3XXE+kYWNfT8LKHt
omqQuwlAeIJ9DrJyr0oHK4TdHPyCn3Kd+ca1LdDziLm2XhT68tVY+GJFY2BPXwB8mQiHtc8W2Rxg
YV0HEZxveccYWIw391FT6jcmx4tvGUw+B84zWxMxoc/XxoghLRlZ8Pa6pS0p2YXsSq7tcuRiZrID
a0K/QMpYu/Hn0o0x00Zktx9upBOGKUwMMHQBDrUSZhyLtpgplQDy+XS9RMtV1mYKkvvmF1M7+SIh
Wrw66NobH52W96hKsY5hXl8B8zbhWQFsBoPnDQJkv93Kpzi9bAW2y0a13+MevYJJ0aloZenqeFqL
OmlBJoNcRtKmwTOQDy3HXYvWnD8NmyU4fg/skEmAdWVwP3E0Pxkwcy4PsKcaIAHRixx5jq+k+qNv
bj6L4mkVp+S4H6u3ATBF17ZXoUtJbAwGbpSbJWKl1d55a5ZfC51SW+1gao+EVOEcpYgFspoyPdOM
o+ddnE/fIDwUsImRDmEJCKiaCQEZL70QwYPVU+41DjPZjzFfzNDJdQ/oJEDNazCb0FRNS0ykFcLk
vGlP5WaT2AnupxWOvE9lHa2BNLUMbfJmpgrzKcD1s8UayABrRckldJ8wqzYKe4jwZzS9zbHTLSfW
JEe42wUhpwkYDSu6efpaVpj9T0ltdAuw5IZepPO+y1q864ZUPqxiIZhWmMwE5tmzXp6Tx4tQDT4z
zFOQLr7UZsz025e6quSqmrd1k1qfCMJVcnaxUe89tPOHvJYL3p112nkdD7OyMWlsGNHK9ClYKIzK
tbHQimYoOA/teE2Z4UQPEQf2fYBPWOVJ6XowLOZwB5X5EVYc7Za/yE9y+RBICdAukZQXJqGVYcA3
BGj1v6sizyNeaPugHpcnv+RvkvX0heEEDOoqlDr1BXRvxO2oCMPbN/SHoeX4qluFYtCJt3Nwzajy
cLKtn7kgMBEWyCLKFd9W/dReeNKcerTt7w8T1DLJ1GonKMvVKJ4up7q3ZW2s+SyyxNrFGptt0eCT
YSGkUZ5+gGch/1rSCf+mLTHeCq1ST2P3RGD9mrL08WNrmE20vwWUic/udw1znQJNUkP6480aL0Yr
FrfqOVGhM9gK2yn94mxUHaCrV2GF3N/0ZiSgo5lihVs6v5eUbwVC2Wj3J4+VYAbCwWRnfoDuRuG2
FFz125F6KEZw4qqwd9olBNMNNjalYrE6oLNwNYXob9rr9DXt4gKxfVI3uGBMN8p83jZJJlFFsVg8
k+DUSEytlJ3wlTpMB/l0xdLlDHiH75Xnp4sIeV6/U/RArMFLw/JwHLA+TCpLCleu7i8RVITmGwzD
2ejOxf309gFL5d1T66s5/v7DAcacmEQYJSA5wEHCphySF1l0AxAlvxIZ2oBuq9e8nTuzX0oWl8nM
pxeS38+PYIPKTierflvQrnpMMZeQEDyJjhEjO+TDXEgYHiqj5ZC0+BMl9zOrSsR/c/SEUxpLO2ej
ANO7tONG0BIBGpq9EhbyuOQVgy6Y7B5cbPe162dmyOfgnycSHN82M8IDcSpjqAeLOghXiLmztccc
jXUwJOWlcXD6y4zOjoDfMi9y6+I/SFXNnC8L1zAIIFVM26o6oipsBGy07+DCXDTpbsGXZ/aBg1mF
FzU9NFDyLWaFux/DnUk2YfgJxiodAr7P1rFBymcTnbx385WjEd+jOqezBANBLXCi/MBV7NbhTRoM
eLlzk7PVuG6Wd8zX508C4xzrhooBFlcxpqfpOigPRvW9rgRPvfvpheW/34yUAH1MGnOSQwHENxZ2
YKU0cvRSbwbe0WxBLwN5Gu3rz/myQmCI1hkmva9TaYIYOCfWPKWALInSOVdQWwQX22MyMojH0TdK
Zfrwm6mQKE8sCNV2oKssmmmSfFn6Z64KmJAR/r/3atBSJIGVMw7CUQBey4PEBL3abivz0O4cUDAg
iJQ1s4Ienl9SLx9uOu8jFzSMNZ1qEgkDtlJhpWVXlS5Jv66vaS33Sx2mXLS1IpWCQrFYAPYM98nn
cRK2qHsJ5q6+Y5R9S9kuIGxUWY82rrxmhlHhE3BwgB7im0VuTm4UqkislJFnbrp3YZmW2Dc+XXOu
Ss1eAHnA2gux9QtqzCo6C9AnwObuo5wFSER0w6QTr13Cwn4bVLK+DSYl0YfE7D5e7TsXB7s3tQxi
+IAt/uQwc4Z9/C5lghQdUuyRVnKwSzzhfLSEgvYtDYkQkydEXh/wkoF0BizcoaZzZVWuyIn2jGrc
ZDtlVmohmM4Im6htKyGKvp5rNWErMoWIYNuYDkt9I7+TD9uTmFAMah9S3bODX3rvvb8dvI4GF8Fh
X82WurcVDkPWNRf5UBkV3JvT6CuAj1BaLFfKQPsBa+xnUQWm42Z22eOdcMSZNZjI+bybobyrWpAu
kGJ7WxOxuuRGWf+BANm2Ov2aVVBfFVBuLNNVm5lBMtI8GEgaj0kkh5pdQJGMJCRsNpfBJORvyVo0
We4gRgIn56ePUt5v2SkIGEXkPATLcBG6h6cW82VlO1B9irl/BIq74LDgVQC98RRuR5otxPygVi8R
KbPNYAZEQuGBRD91V1o98lODRYiserEqMIqDwEzwS2bsm3XIXYSBuc+zkiWVdOz7Kw7xLag7FnHC
Yqf04mteK4vUG8tRiO0wNE/YqVgNeaZqCLvdVAPU5Kc46hQ5E0ubhyiIw6rQ+xllWLrtg9xGQN09
qWg5ga3ZJiatIa8dsVrsc+XXPzpUlH6ffQ2JuNfeSrHbu5sDE4LhfU7bYtmmQ0K5pQChT98NUaTN
GgtZGf/bcDYwq8WE6H+9koOGnYXfmGdCG1pAQFaVnIgQ2l9sZY7FpWuqw4XHq92xctrNz/rFbnSV
nqb8PZcU9n/NwsbmAaVM2jlPWYGvtOTUDhJIU9qxz7fdCOrQ2rqez5ceXlL28C3Q4VfjlOWWxDe1
5rKmJ75afCgXt79/aBQvs+PCf49baxj3FYLVAYZHKajC1RjHSTezYCg/77yXm5CkmxgwWRuaIneU
fc5RB4xJjy1KbwSB7hpgjo+1KJuQmoV0BHL4dTbIMWkml7Nti7IELDLDg/5u9tdW4m2juQgE3dSm
IjNXAHeSq2ytmq86NeawfV0JBLEdY2Rr1HTfvwja6/j7IPP3QAsoYut6AzyDmeSzxARv8qu7Z+ky
/CKfZC5r+pKmhpLxcgqkfCrSPN4943HQm2hxCDdEFqBFOlIHmwgbmIlGMXXstq320R50GBYU7G/T
E4m7OpgWfFbKqcWiJMJ+eca06zfixWeiUAS3qKFm4Ih/3t1jIFuk8Q4CguMmvaDhcZBGy5kVa1GP
AJo7X6z02lHCKUw+ET4fF7T/eqJbwUaNACyxupFAomIuSDHYo7+T7dM95zDXpbqYlcmvY8GGuePy
dE+02oNkqmXez1w45vGrgS/GBAuJTCts1QsfZoLXB32WkmVnp1cSuzX798YkDZvweRPW3UmtipiN
2s9miFWG23InyIvDnKdKTUwl/S5fK990qqzfpUgAi2Wo4fJwabAZJZjhJF7xr1Os3oQ7d66tGDiy
nStJdn40uh5IOr0QuqjrecdtD6bWMlfTHJ78Ae+LSDjZ+zNhpZTtU4kmAbpkJ1g8I7YE8tGrpuvN
nl2xLMG8bHjOXPFVMfrSQa4ypLljuIk94aAtEwwsFpV4tICVUBvyszA5XYUNBOCbSba0GucHFAZ8
sAwryMeIW83XCamTgrLD83D6TtsRtudC3CZGHuO1GBXB2GNQL2qFUYCImGxttJUY6ebbytc6sJ6O
yl7K/knA4vSgWffecWy8oQ1b+ntqQEPdkr8J3HoXZhEzSRBBL588WNrDlogYzimugUPRnlOG46Q9
rPlveMEVPaG+LE9TQUOLolFbJai3TIWvv28MRGbTuGXSgEu2h8+4UmcdOMq70nzZXaEOlvZG1ohO
UMoDcybqgKetCK3ilVKh+ZY5pQkVjUGCfLjSNKg1EO79oRlxhw/cHJkRC2x0/jwgBKWq6VMTNTL3
LWUuaxCrklta8ySro6H23t9GN1wr46HtHiVDDUmcNR5CivLnghKfwSrNZTIPRwE2+6tm/Vwxnix/
X+JavWl0IQTs9jjmIp/IoJsKWA+L7RqdRW4o0DugsflMP+bnW+iiJMqEy5zd6R6+c1YLZZJvZcze
X1fbqJk9ZX80OQaM6SjNAjFAS5IOa2ophvVBmekpTFA2fZhNZ1ZGUS/kisC2Lxu+4ytz53e5eC1Q
50Qk1xuaz3G4ypKd8n+GkBKAru8QC700BWOmwfCtuWr1s7Mgg//65GWQpPZthAa70HtvO67Vg87x
yV8JRjN1eJv6dP0TJeIThiHH/A15BzIik3TIYR2bbzQLELuBMtPbcIUzjn+8aE+YlF6oqP5S93sU
mCyuWLYk3P/6u0IublzmcSCrrnV6VM+RBfY3onhMi4UEQGpCDMEev1maBywlIY8neWlQuHjW3Xg1
606yXv/M4ds1iBa01lvfkm2gJ+P09d9/an09nMnyOr/wyPCATMbpZVJbJNBfvzk5mBCUagy6scMm
TkrnJHh4IX8ittDU+WFH33ujdC2r7qCjg3cvFHOJXreJa0ALe1DDcGJOUsQELRmhXv+NqZmufqJ5
KDo5dYvW2syR/G0PbPTM3eZnrFpaPhwzcrA5TcOkS0tIDdKtTRKgDuv80dU88OGkCOkbt0UPwwjZ
oq/F0tSLHw4hY7Eb9wgcVhZ27O5FaJCHUf5KS+4JiB3zmJOMs2PDRQPqlk/6Mzzhq8N+cNXO8AGd
QLqHkvyCfEi1WNWL3N3AhI0Ni0QopSYGd8VbmpvSOLBrIQfczt+yb/X07oc/WmWnI2xWJWteJ1JE
1Id9BuYSKUgCx4fZWWAtzP8zVS4g6EGbJEa+qrmcYdiVpa2FLQC/9Z1RS/XjD3KtrbbQFZbZ09mc
9OhXhjbbMONoEraY6OkyYV6qBr1l1ALiEp+4BcG3fhnqCWInQlOaLHItT5eidIlc6OOIEq3og+z5
f+755n9oVGRJ3fD2ImG+7pVpJ+NS4hHBifurFkaZi40cL6D6TOkNO87xCgH9gAQ1RKqOZ+EOjzs3
Nmy6pckGOGgiigbRuz5Z6m9iBqqTzuhCmKKGQu3vupM50PGmhaMYpzhp58JeHeB4XqdVto+psw07
CQp9ts5MCvX6gxlSXS41/zqsLXxTDp/a6/4Q0CIraMGPGyU6U+jLyF/z0XRfTv4s3Rwh8ctfJmcs
xZkgDsMhtV1AcclsB3Fpjga6DGFAo3jJQ2y6Oi4Vxk7szdaYsTobI10JcgxnEVcPPr3SFxBi0fMM
YqSQP/YjW3Sv89dXxcFcR7nJwZuBGP7NbGDuPS2WFdOxfglhxMfVwLllysi8YVAnxjuKCc6imuyN
xE1XeaDO59lZry/bKmrADCXvxj3TlbeVhDfy1ACvlln2Qfi+ykCMk0AZpbLRMBc/MY0rbaMU0UV1
p52j2ZWCTxDdbSOVnJqK+OUB+zXvGBC8QcaUVzPdB1qvxJi/QG8gE6thxqtDZ8J3/3xjodp0qgVI
bhAfutxU2VkJ5X/ubXUARtUYRaMwdigwKX6nJs1mKmKJDmXPhrdn0saPgrWqGNh6e7mtYUilJZH8
w10yZO6JFdwvObNAskWX0SWNPrTP3hMR8W4Inud2GeFDyxVooxN0AtTur/FvkIVGYVMYDVRp0oQt
bojjEbxEwH2voYtJtdxdkNOPFiB4pUruH/tLgYHTolaMD3+9mn976Hyiah/WE/cK9FiLZSxRdYQc
b2l6ek/CXeLOf/pCAb1XKSRM7QHx1e1uTDxR9Ko7Uxs39RQ/Oalo6qXnRHvYPN/AUnjRfaZq75M0
GXOFd7iViby58Gub6TwJdtKB0jnbVRlQnDegafgEE0NxzOJdpPbxE6fQ+HzEpUTjf+gYx/40oDNN
aFhXIpY8kg9trGNxLq/777w0VQcssbwhU8jrozvcDItsrFquyHjWE8KPpbb5PtofqSxzhvwZGKLP
Zfh0PyIzVzINrypHkxA4dPxlvO+36sMksM0At0YC4rdUfJQ+kL73aVCkEv20xeCgS0HQv0pM/qgJ
a7t7TopAxf4hU+kAvDccCqd0ApPKP0MvK/SqizmjsXh3Eu4FQC5Vsj7RoKDtlsnBcOuO4o2G07ZW
31OYJAMaEEKpwmK691p69PBHyR9W95Lu0RGdTs/WAtgjIAQRCzrk+UTey/W73JTyUGMEtcvo7EJN
UHogkDsO5V+V2la0PNazOuJWx3ebtyAfeNtBTx8X8UKFL1yfkaRhntTvxhMTcamfF2RgOB9w46Oz
sHqvyAGdrEf8MmEFlg3Lq4ZgWgwPqJlzBOGF6bDmEg8LpV+LiwRS3deOp5q1sG9BuQHOl2zkg03V
8o/4NDu0MRpyHYN+1yIDceblWA94IOCle+r6mX3cTrcTaRjDjhhGjMp8zA3Rq9iPUlHxU7oUU8P4
ZitJrih5yHjronS938lismMAxiRKf+lW4HIkSCSsx6TJdwxcdnNOljtpedKN85GWyxt53j8KgRP8
7XSOuAgmSnrfglQKD0IcfLpR01wKb0gNQD7VSV1o1DO3X6o8kYUFqU7OTxCbuc0NLemWQ06CN/5L
2cLrsN6WCjfpX18aTWy851P7gih5gwV0kX/rjBEG2S+tf8/hnRdA31MssYOau7RC5vn4Y8WVYtw6
1fR/d53qEpR4J1bggivGmVuXJP9PYWppaU88zoClvmuLI9csA+Jr48/aJh8bMnqgxBUD2dH/g/FN
ysiM1WlUFALKaCofN5PVmd7ChepensBmZagppTPFO5KIVlM8wkJu6iE1dLGx4J1k5RPXitGYFcB5
xUyN+1/klCdG5IM82cytUnEGlOBTvMyN/9bj9TwkqbZj3tJit33OeQYUxOCLhSnE2/Bj6mhoGUIE
CEXod4T/GRoDOO1JiIpoZTjdPUn6/cEeE+8R7ySXwry1JF8ml+eE1EETOggVkB1JK8f/xtqpQuUi
B3fiSfc4hMyoUZ/lZ2n8WCHzimkTEtkiRCCw8ikaJ8qBFvolSHLpmI9vZfTmcQdA9srN+dDFRYIK
UF+ylFqfb33Fsy+Whp5Qcf6HVPTXkZzWGr6pPyzZim2RBJHeauXR0mfBPT+f9K9XHwFXVn1bSeQi
FgKNFUD6a3CkPrYxJMDcbm+Mi2+GJlPPVS8Td755FCjiCsyuKTtksboJ3u+2InW/ReC9Rbn5bM8c
w3Bk419kEQEzK4god7DgsGhZFvZ5vUZMamPebEIzczxBeWOJ/54TyscR4J3UrVXH/0Aq00ocB2Jr
G7x6jsYKpS8myoZo9G2LZG3IrCYnLmEhVwgORq2aB0/nytEJRk+chKNB7xb9KeAAtci/jNQCnEBd
4H/SRnA9jDJv5cg0YrJoNl/NEwEFi9TJm2zH+svUEQZedBzkdNdkx77z+c9n3AP1gj/+0Vqc+6XJ
MOpshOfJ+Jv9eFsuKQ6pL3xKtsDQK9/SyDDj1RBladFDljsnEZvwYPzn+tyMGqw6IXCoby6kRQwg
TGIk1zDFj1PXx3CIjpHQJEMTT3Br6ERdFF3tP8CVA960Alhv9A5usFCMP0NCz4Vkzm/9gfR0uAjV
J7u5ODwmXSzlUIZPYH2GrbOSg1xGQwi3eMDjsuBVjwLXOwVgFCeQYtJbx2LT6Euy8aO+CCCHbrpv
nEBwff0beAaO++OuSEweyYb5NBqyu8mxg9nT/xXN3U2MUwd/TXxM0Z0hupklQns0fHTHs+XwHyhX
M7McOU7WkdjHfEs/xXxEFN9DuwAmxanIhVXLgMHtNiarabCWA2D20uD0rpLJ4FiYJrW5XL2syukD
Ung4JaCfVL9JEMSwFMx5fCBwilhv4YVR93tJvKM9fbF/j3iZ6x/tP2f+kHaGRVUqUKUQU6hdXQ/i
m0GdibGcHBy1h24TX6WhPRqWNFjKRPCPxeBz2YH54+sh1kZYtBCmuZiUYYwj8aUhUgTTpbYL744A
70coW4XAxKW7UfY1Rcn8IXRNAK7+5IUYhJxp1g8BPqNSDPbZ9fKrXQeZlNUi/FtKto+DB5W9b2qR
ILBWB4tGjO73wt50UZ1kSV8yzNNN9wHaJi8dWX3nzRyR/SFaGH/V3h8oXjlc5i/et3N0HyOFCqD2
ZEYQJaVD8kGqKmqEabjIaJw5p0TUJfc3F2ArvNAETkrtQ13tLaLf9qU1frQRa7AYVur+wdTzvryO
DkSxmjsgrydMnLRquRgpFg5eBVABtDH+hhtkUFCKFudh2mvEJZqlnHFE7Phufp4x2Er9bo9a/BSf
oCXtSIbqdVdFL8d/4aqwqXfhPdurfLDSM78G9LgCTOSAADb9eKXLBzs3BEscrj+tWqwzn2gFqLST
nBUO2Uf93fAFQYzMovbQfHSAgjD/pou9meb2nJt1mduo7kCzNqs0cESPpGsUgqCNUg3tC02Z89g7
5Vh20V9IaLIiyc9diZMxaUHk3vnvEoYdfpP5Tgk+5BCpZEonQ+ni0Sr8T0+STURsvnRNug8U19LQ
LoFsPoP5TAljjrfy8odmpu3y92mvZSoNzBzzIdnoo+nzCYDoUiFiYavTafL844YJ3WRo7IqG+mKa
db46kIf/HO5fUusqwJQ11xPtYINJaLimLH94Bm0Dtul3M9Kv/nitstDISUxcnwBT90kSnzj53IKk
QMWEHPAHBQ2X8NhQIpFL5AKTcO0aNgZTT3mlIM3tZkqYYXgEKVwsmvcqiNWft8v+4a3MNMVOyMqF
0cZWf+KASpdLPEW+gRsW/DxUmVccHGZaz8DaacXy0J+pEhhLIHMo9KUI/aRWsmMaxwYHnr3zicjM
PJnIHVuPwMUWnvvINNAmzeDhZZtlw3na5HnSlGHPQzhmKp65dA4OzM+fbibIigUsEllPl4FIVqLB
2XZq+FFOGMDckikqkZujit00+5dN8GgrsroPpy7v0QbVqgwAQpUpXBW3DwqJJOTaGc333fxgJ3dC
BioGOZQxzoxIZQfy5xe60IK8fWBa7qryzvnoD2xg2nUTg2KnF16xyA92Y0ZHmPA3BRwIM5bc6/Q3
uVXNRI1ThhOg3dESggy1+0TGvznaBMK41T6/NHAoIF4YI9jF/xT1/+V0pI2OE+b5Fs3Pw1oX59t0
x447JTF1cQ7UDUBlB2dSZ3zUwsskxHD3YnTu0L7GHWZOTYz86qsr75PYNtVOL6dQog4o2xCQ51Bb
EVDA/FcXcPMIyoLPJkmLrDZ/JEnU3gjOKm9m3r9IIl4txSZCcVlv3UFlPbTfAsgA8Npj+Eqk94J9
MikWyahbDUIk+qoPk950GIw0KsfDfKrkUfPZrf4dwePipYXHdYKF3feTXm1EbBLftciqAy7/4XWW
t6UKxJvnOF46adTKsUyEEFQaLI/4P3agTv4Epgga4qV7OJijRIy6BPP6AnRk2IV7VxfHNZNAb4UT
AhiqWESRQtesPMLoAWBlNUXljn1DechP4T8BL+GoqysdJ/6qHU1LC821DT4hf8+gDwkHW0wqIqjX
bS1C3M91v7Gg/cL1fRF8spUTzlJZgspejK2a+wriQZgaUXRYKkNV8bKRSvK/GPlwkF0J7F6Qab+o
9lFr9apjyZ23RqEHjOd4clladORs2rvbu7xmrHQLW9fNfv3ZzXyW5Y2tN0z7wGI6WlEZCR18tPqV
qRocyakEUmbWt8fQ0gyL2fXJ/WdWDP4MiYbKdWWCTEho01PQVviyRgfgYIPL7eWAnv+dM6fhs2hi
ct0vVl3Fx7hxYi29jMenxxz6PtUzp37ZDZ82UEoWghhRsJaryC2bMhO8+WBhwEbIjhHo2ZVW0X9F
HVpvMUwlrOq+orSHK3n0y9LtEMFS6LSPHYn2xCsspqsoU/I625TFiz4G6fbKm4CBHdMZqxfmsE4M
fvT/iJ7j2/DsdaNo7JlczQY4J5AmQ2iCzcxfNlmnH79e+wwG08yWfGJUwtv6sFCLxNbLOdUN1rii
iOCbC6KxaRZFsUCVt0h710SLgBrbg4f1FXjdskeNBgpYX0fwtjgzNclP7dgIFRtznvdRsu9uQQ4L
3INTdiry/u4CdkhrOGjbssqNerXrV2a9YqReJmxg5E8+qTppWmdEkANXCDMMngN5howCfwnxAdSy
0jwA/07kUKpalegbcY+PTnctby1j6by2ce/PdE/Q2MjPuJt7EglXGwqRpBN+OngDZ1oQe9ZHZI95
Sc29AtmX6Fv3kqZP1ThvZv4rA3UZi/Bg7eXv1TKv++tmjoFGrgzi/PYbVvb47jtzg6uPabReujXb
SbPj81c6TrektvRYSXjkZjbY0P3i9R+ZAu/KRvpZd/1Uw81inOLt+9gyeQebIWEjuxDLrfwjplHL
ZMQfE+Dz822uUuCTSArGMR+kGYMazljR4eIIKlxaMnaZfuQYlMulNz2nb/SMo1M3eBn+mSC7T9Rt
5KoNeDbKPBWzpHPQ2iXTSlKxiw+m1mVUcQcKUWgLBKvLmK2ycTjwLGrGxG4FXdPxBa4pkML6gbK+
qCu+9neXpNhE9FRDIk0cZO+EDFylAgAgcMx9/a7dQzhDqx0jnWUx/XmaOWdMotX9G4/KMYnoJJvr
hmVQyF5o25E6PRvq36Zdn8kG0gQNSiXS/7wp85QrC5bSjegwGjqA4r8fR7VQaC0qSg/0wGC1lvrT
aUf2Sf/IKYmQ1sjrGFnAVqedX3nSCodRgBvuv+2qdRrHNIjsCyQy5saD052g6/RIKjQdu9giv63Y
v/UBDr62aiGwVaIiMl5O3u1E91ngq5vPMQjD2eW4tVQatFnF2Lg7NzZMMy2TyCp9FynH93lJB+Qh
/2Ict2DoDSlioHKgPvdXjwMUXXR86d1twekBBljHq7D/mG2ibMGMSUuzUGW526JMOt3FV+JJAab0
PfRYT5j2wZ0J/0NrMQbcKoPoRo1+TRiOe3ihkDswjIIM+4D/QME234hIsWvPVjkTlfgiP4e+6Faj
SO9jkf1qcGxpsWT2TZIImIfVKHRohUO0Z+w6qX5S0D7VEdAySw+ATNroXlAPSSl8Psfuborx6Icu
KeD5Ye2ql0o5AOW5DzoFjXQjrajvWQj8xeVNVlv/TjzfqK5vz66wNaT/umwtD1s9YNRhCLrTbv6s
lOEU/XeANlLfGUBxhV3VHZ8MGpWqrqk9I1Zbuy5UMPCDSYsKc/dKi5wPpj3hd9luHCCr7ZbHIxBB
Zh8VskgXRDCLop8m+zS2bR1l+rNZA+61QgdhPGXGd/+0WbdMz/fQC+0Cz4XN0k6LVori3ayGWTQP
Ue39t53INCj2lKh/aPLQpdI3nTvBr8xZPk2/lh+y9jfWeXvYPD9ICDyJsRFeQq82GbdueB2iv7ju
SrvJYBMMaKnKs7N0kdRH9Amf4cPELMZLLljjw7a68v/f+II+w3xkatwLz24HgwF9ZVMUjIRoxMhG
l2ikNN2L9aowMK0hoDaa9SfgT8IE0hT8PHqo+XwCH0fuW1q9iqgHFN5P51w9wrJ81d4B7FAgZ7ah
x7udZ4PoWqqNRgqi3sKdP2d5c/FaiB4mbgH/tGTsSiBjGxtgpN5RUsrn8srB9VlEh2+b8eUi9zpz
U+4UAavRBTMw74WDBG5YkvH1BIwaufpoVIhDK7QmH/hsaUSxtT+wnJJZBTSrWZss4pc+QOq6FR41
1UdrNMPiAQte2jRBlSvU2YM+XA4UHREzmOMQwv/eOe/fKaOhdgFyCqrl52FvDMEfa9nOdtTt/DzX
JrSMyk/4d8caOM/I96VY5pxd5qqts16kWbLjlzqzUTJf/+BrpOLPzaKeqPZvxV5cntfRmwJTXMzA
ZwOpEi1ZmB1CGR3TG/66MNH8BtXEmA242qK0npHGiXT1YbCijgqAIzJB5zVZKFwn3DQyudl7Pp2z
BxrS/mo0hizhvSBqSWUaUSsdykBcA3SwVgPAn+a+YVHcHXP8OK3bxQBNfswKqxFvelQEwzqCiji6
zui44vvaZpBVESOR9Y3Xq14OWihGMTz75gX4fZHbcBpDFO0taChVN6o0uBDpYOSoOBvNM6d/Y+8v
iwDVQq+eS9hwkCvdcGtdWUqX1owBPyxpG0eXpP4a26km7Onxbowm/uf+XfFervyjyd1lME165Kl5
zqAn9EP0mUQom7Q70hNRERwJ65zZBlD7UxE+lKxVcl9HQizXDPTVwzmM0JuGUlDdJy48VM5ywnCE
NtUAcBsaRdt5x/yD1QaYj36vrgfXVNc77v59HDtYrEzccrHJXk5hv3Ydn+NrOUrfV024xZ+eS532
Etw5Ubhkl6I2bkX0IW+0ejpNK6Q5BOSQNtffCv2zBLYuRb1SBmT4J0G8Th1XGyPbj6UDaiWri50z
tG44uaXFntqwwwesrVYsFtTEvcG7YT6tfbWQsiALzd2MfGk1oq5gqhvnMRStrUAaxuWPLq7uwuIZ
JAfOrtHKTxsYghh5rWFHgPxSI+7s2swWENceTuDXMttSyim6UrHsZ5/nPUjmHqjOU6rzgmmsfzpd
XE6Va37ERN+Gr7HHt4roWzhAX9ZbQT+80P6mgUEtEshOhKw4zjDqFoDX1KJrUtmzWleXzWkq7bJ7
lP6sf3y6cyUtDe1rDkEJ39VsyGC4YNVOQOG2uwSAbY7CKzlSFT/hE4yob9atoFpSOsah5gVq8gB7
+5ZU/pO4c9asBsPuX4Bwz2UOcTYMPNbcSvVRUGGmGuGGuZsvpcscPqqunkUvV9ppfoPeqHviMJJ3
NNJb+7CR5aXNHVp1pOwtWVXBdQpVa0eTG54Vjx/rcbzXDndA+B7EEuflni0QUpx5knG0GwX6+Moy
qEuxik/r3u85Rp4Pth6zNWIAwaGsNnNTPlWuadtOCoVqV1tmddZVgkpZQqeAKVGaHGzKw89ihq3C
oKfZ1TC/jipSJowPpbdoP3JXxQtP7AEMbFmDpbBkT47wGkvABxtvIiL9BjrHwQmbdqG4rs2Os8Qe
9jp1E+lNnMEQB3kJsxIe4V0gqmvCIN2giUq9G9FY4OJtH9l4iX0xqiFEMLNezUO9bMwG/MRa98FM
MT5ZdJK9SjVI5KjeobJChiL/NRkpL9IMqexYulZ/mtunbKP1X2c3tC2dxe177Fzd8xwp77xFM6uw
tzxHbLOU4b0XmorLYIswPH5LBzKbYrKJ7JdU5fGF63jdDfnH8JLiVT2AnaorKBTFvu7xKZ6gSU00
sq2+cRKgX1q8Qfu8dXDo2/zB/lfxeZFLkOZLxdl+xkna53mNhnsxZSNiiUxFMXZgJv3CH8MS8sM/
HzNTNAlGrKEP0I03a9Sqvf/+lNa3rmkm18wkLulsWLvbzbvOoyKC2WmVkA0vhXkWmvv/6f1s98mi
DetcftTN2xwqGVYlLzd7NKXTSBzCj8PdYm+GaHjmTXkdj1alInQUj9vQWHs5Gd9fyb36FGDA38jx
vkul9X1kergHOof4vb/kBmSE8ZfsqqGHewuutxxl5Kp3lXZvRau8iC8BQHuC/YWXRvvRABOdCHFE
vo9kclGR5MaNWfXiIqipIEgtjloiZjaWyQZGR0HAv5ZrieNhIFlDf4u62f5bpMJDhDW6DsM7AKNC
TD9/f/Q/rG+dGn2Vl/ZyssBN2ZiuQR59yOg2nPeiMeyJf8YcXmAqCo5NVcv2wDBLINyBqdwnIoD+
xwXZdQ/zd7t65S3R/t2lf1Lv+UemBfJR9jxnHhaHsZ2zcp1Q3hyN8HVxEGBfu6ZgWnSVauIxX3qD
2jrc7jtD5ObEulw1OrfI890n9JsuDgdRcM3oQm+Kp7vZFC4Cb7dieFAJDATC3I67uWdnhzcGgTrJ
tmFOoFfUHAd5rgVq06DafUPAc6va8paMMneqBQPGsp+FJYTHEr6W6cPcjHV6IRq9ZLns2oDw6KnW
avQVhK4AsMWg0MVmgLvRySbwkx2a6iFWHhesWUE73rJxCmOGKQaX/o2cBCHcFlrn5+21tecdj1jK
lhLvihUIsgLNekrbFmcAJGx+RlKTeObSRXXDvm4ccZdbRbfpFIADz24O1I03X/AxXH/AEml2xIOi
mL5MAwD7kO4/fSSvmOG2mR9QncP4NfRVC8fqLdQeFC4oILn1sh+vKjfE0PWUkjUu9iDBYrWWoP2B
vWIo16305cb/Mi01jOaZ7j0PXlmjkfKYB5BtBJXFednd0w6iwcTAh22EHWrW2XzyDrJxBQ35uS/I
d6BRDLhOYd5e/RCwtG5RQsLZxtY+VLsTuvLO+eQoje27nOyILabjnDJO2uIp+Yt389KDOQ5RqkMR
Rh95y9ytM185YetHBWgPM9h8cDo03Gq8a4dtCRr2hcFaNQRMzmF8RP37IMFmDj46hvKcY1EBLB4U
OKt/OSboU9Ze9vrLlGB2UlViJn2mHgHUDmdlJYNNodxvqlW0TumfAte+fm8Dd6GSSu6z8Ms+2pX0
ruUoqNuNH5ez0fW7Hr0Lx/l6WoozMqDSu6qp1T8G39nxy88Zo7W5ZYBs4S9ShiGC0n5Xnciuwyhe
clWl+HozaHtAGGv1Y8pSy46aJv0VeawT8a2IdUhRzLV6plQ/tjCGauW/yPlTBcTe3Lkm6uJNHhBV
dq0P7kkjUwvm3Z0l/b/Wotu2t24ge0FbDXIKsu6zCYpcl8RylSm/vUr6gYVaaHRCOxDim3cTmwwm
zMgx14Xe8gwtR+ARkrT06VC/N7XOk6ym9giBTflO6JjDxrsE8ZH+fUycM/U+EVJZSu5+lsVYQaXl
y+cMsQHNdxvpInmLpaitO4Bx8vTV3IQUN9yM6FPdPw5zQPZPOiS0lhTYws9ldRVKDIyYPg+Z40s0
LWI9CBYotOvPtt3Zm7ZGLDWW7OJAY0F4+PHpnH1Z/q2FvdUYxk7rKg+4pt1yM/15Z7rGiFiWomZn
NqlPjOAFBfCwyL9I5ZfXom9GSoyn+Wvb3IFfSfuUP2LJTLSyBgXK6OXqyiT7op2D/vY7gl+Scv5M
7OBCRvpT5EyXvaODNnG93mkytTnjAW46EhiRGrOcRZnFopSSckQQZsnxAJw3eQQ8hPBH7oh+GV8w
NFd+6r6bi8k5yvLkAqeJ2exYM0K5P+5tXL/Q8EHDYBwwxxSU8fn6ijW+pU4frh8pY+UU2Fybihuv
7FF35SK/L8HgGoFJnG+KVDGUTE6vunSO0OHupq9LCoeF852FoZ/jRMdC8G03KOcaHj5RtQBXjOkV
3iyk7LC970DYroUxduOJHa1d7i1G/QJi4hQ73YZjT0ZfTHjoj54XO4uydTpQc6mhRZB60zO5/KOu
CQmS0FClB5bWZCJkUbpmk9aG3932F6BtV/xgL13b2M0IrnkfV5uTSlZ6UNMGRqE4DoIz7uBOtE4E
D8ngUK0OoS93lTSEI56YmUi889iGbgpdbjLv3OUgnRJu9iPZnQy4pXrm9KsgzJEnf8xsSKCoDE8o
tXjLSIwsQTzknaowflCvRvPdiVTSiotwt20Z6GhOcuzns7I5ylcI8sLQ54kPiATO2UmDSY3Fah0z
2jvlZ3G/skARxpZS1O50hObYCTzVGkeuDHYZkZFDpz7313Kyh8jnPhgd8aUJTYwBYC9MEAOor9Yw
MZPprWK9B2eDUx97dN9Kki7gv/5phSdhfK8zdBZpBZSdeamWXJWjH57Jcp4y4DjSicsFeAWVAPBr
mms328BxUm7BsDaJu47OZFVG5sR/YQGyPpzaYhLj+YJpxW5ODLkPHbDbr6e76BZw3G4RLGMwt4PT
9GyOSftesmwHZd+fRlaUBIeAlWz4jUay4d6hL7R59ssS0xX6xYVK4BD6R1KWYElpyfIZIMw03Oty
N3n2CM1o/J8eiCZMlvaOC3niR4GFb195fggL4agVskmcT+sRyRmmTHIvZ35ByJ974FUdNUl/GH/E
bZWQ6njVTXowKPsDQuWbFu2pWfBYE+F0og09xLX5EJ2nuZPIIBTaTaTBXFe9gsVsE6N+RdoA/hGJ
4h0O7kSrplP/VxrFT4f2VCmwBRJciKn72wBcYebvpq1PqWeRQnhpdMyDOKU2YS5NEe9vT95j48wS
Nb/VqEHTyXNS52x35vblKm4u2NaF7JSrVRwGaZESjBnQwsjI0YIV4jzsgrcdZQDDAuMqwFImc7BS
XtMu65RoIb0crbSa39ng3EdNNiP7QLFFKn1P1kIJPagT3Np1Ph3yV4yfGwPwgmpJBxUyMGSCQBFo
IVcJEGquUipWRj7Aqh5zRhFHK+c/xjIhTmWxmnLuqYFkH+gFPCkTRMLELsjoO+i/i3kTZa7m7VHv
rEgCFuqdBXWYLZCXe9SQLLb+ndMolZpXlwQ4UofWPSlnQUFio2HmwSESdxbAGkWl/pD3otuYh/VQ
MZfLWlJyJyiuu9KhQasqetVcdCAVOOO4RXc/43tKOV2L8BkdqskUICJrCZCrObZyaYehLxn8spmr
N72Vfe+K/+ZOdHJqB7XU+bSdi53yUqZpv7ExYjXvKxJaZ6bigQnmUDDLCE6pq12aJD3GqLTz+Fw+
uKsbAWFaxdITGbxQRPOjMFV0JKvOoNGvrJGwIpWPr8Gawb4dpDhS9vFeAkbq6gbK9n5Qk+vphTiq
CKOfq43oCzDHVfwLopPlzUBLpnyJb847oJV6ROveUdSF0HCarKzO5fAQydeqFRdITZ+jCULQIJMr
KkuDHuZgF/2TOthGDRyBQX2ewQbPHbE2ZW7K4Z5ZAsNzfFufUs6fhblmoDAfh6tfW/u4rm3TNj2F
lDf+cut8m+n52n8lmz21tQvLkUa/kEqIlUu6gPE8MxeyVWHzOPkX2dA1HItGwN2bkErpdSr5ocP0
CaJTeb0scVjl0YZ7UPbzyLMvr8jAMueK+hTO2VoNVKAKBKpNyqKwYloyF1JDAs0T+rFOylfl/UM1
fJfiqtdwBrs7QLFHJFUTy/UrkR+DfTaD/yCR1Jie+Msyht19rTBbe870bb1x03v0X5o1/1frYhx5
NSBJ82bJxLG+oG3HaKJqUMRGIWdy3DEXXnUgF9lb+LU/1CyfXOdaB3gZT7jmmKfT9czGXkKDrjSu
35OW0OWnwE5D9MWc7RqVpnz3aHS7a8gEJz5qIKyc0EQXDPnuMG/mjeoGe0urKcs+l9q4K3VJqwYO
DJaAqrw0lsne7BBbFaJ4CbPefjcNjYn6HpRqkejtUU3HtCDXBrkQWwBxPwqPetw/tdR/ShT/VVed
jUlHEVX2fd5S4GDBoMoRhgW8j1KonjTzmQIAb6wHFptp2f/6U3ykzYz+GPjnoTN3NvxUu3Z8PueQ
0Z4h0yxx30iUeX10XnUghDNSqUoU8oRST2g197x2dEzPUEi3CHg9lvyoYT3GkOKSbqAIjMTV8zWu
6/wBD37L73tIOJnvc8XlaLE+AaHdlv2qgK9ovwr6usOdtmbxII2bZ1uS2A0FUttTdzfdcmEKzoEh
QkVwvaylPZ1wHErhYkDmVHIxHMtli2NizbPDf/A+SbllouNSC3lduL5vWr/F5uRxaZHatNbNKB8T
rF3gO7g5Pq9p69u294Eyg9ZFp08w78R5aZTmAg4yH+PFlGqhAfL+uEaVxPFYVSAXrlWqowOCZQ11
VMhTMZB2z0EaFJWSOkKCZz6uDzmpVUsdMolCgeMrtM4PuU2K2KS7mpg+jwq6neUVC1BKUBPwqSzy
h/a6nD0U2CjzhBdOUzggugd+R/U+Wf4dSgKkR8GBfK9iVUSYhPX5MSsRZ/vb634/C8MCz/3hcePI
Vk11U9lOLDPehdc5ISwpGnw5COvL8CzsKcvSaFAc9j1YnCswmjEeH7S5vLB9PJFz81HVd2bjTsUa
roNhcCrG0t3odUBrL/1gQbXs6apIo+RomGhSIgq00KHd9yVNdOtIHLXkt+sH/VgJdmxhbcOAnP3z
psLJjXqm1iFEp75kqiWO9mceyy5tIJ0BLLsw/YYzQHFJDwT1x62/t1C/sPLYETTufz/hrJAOXJAu
+HYJcWFHaSsZNTlcYV/wvw5sg4ZWMjeBzKHAfAhG5Bep1yjNVDLbYM/MbP+lOqBdZtAnuRAVxFmd
W6+SbN9smMVpqXEBwaXrRSfc/q8eie3chijNusKeXQnxoMejk8ufC3GT2n/ZfXkkTmWoXqtOcHxP
G32/ifSPo4/xsnHascmyHKS0WQzQXz4GxMn9vkiFSx1D+KGeVF19ER/dlcasqSmN10t7P/s5aw2+
2GcVH9NanzwOiScRV4/KFwDUBCtYkbZQMoN1rX4BBLAgVdck9WZ8jklnykpE8pxYaBPMpBcaknzj
k09kATQb2BeZPESDb1A1uFfPYvdp5dgZqdoQo7kdh/QMdmMAltrjKh5gf4JAeMMfFG/RrBMLCqU6
ZEee4a9Eqnz2nDINxD4AId6aiGWr2rNWJfR+yDuEDvRWZj6OixMh/d0ugI0kJZaDMLL2j7jMbohr
BeUBd5JwMAgaPacd/pfLgsjCjrkn0xQ1E6tygmSh4MB+T7iVjUkFLePIlpANxjt7cbmYH8v/Xdy8
Da9IOYnTp/0lRFYPo7DzrZW9pCIzlm3mbJGtds3xu5gKe8EB1TOgtattvHGOnvNcgpILZqANtDaR
7m9mzfpRq/AxNXqnYoe06HRWkSCO5qkg3j4FOmV3yGcG4Q9735YVD5J+3ofC9b7AHVBG+etEq4ba
OPrNrPEL+3CAzf6FPwcHfdZ15jW41ZiPoCOVxZ8hiWztIEJVhdwI6NMeKLf3ACCcnkKQT5zNYda2
dNDFVdcQZM+t4+e43a1cn+HardnaHiAvU5s4xuQHz6auQRDrD/v+dX8k2KiqgrbsbFo13pdhO9o2
po/Y6O2LrRbrKdHQkxWrApa9nXol//cEMltUDQEpvoNTopwQnwj3DlXVaXcLPJ4K1BtAPILIDldK
nn1/M4BXkOixSYYPsmBG+NqXdtd3RyI20bww3rXBxJ8TDc73Y3FSZEg7lfFaI2fzb/DBYNeUXH4P
wFCUqxn7T+iiem9GIff5qWF8vkCySAyaIvv/g+zQP4EmHOPcjNts/eXfk3Gb9Mq2KlXE0v7A9j7I
z8TNBof9m/7q9y417tg4S0b0gTf9825rfUlhBZ+baMhLSqrVzoLfUDz9iZaqEx7WV+5KM0qdDQjg
rz7Y1TFl6TmGSDboPl5WD3gnm1NarXwxIpbcSj0EFT6+v8JIqZXAgLMIBMUGX5l7uVK5hPiDrsBG
cy7h+QM4UcvPjnZGlgkQjOb4nGakmcqCtxyUP82bB3GQAdHV1dEiGN5m07fCne8XSJVND/XVRLun
F9I+wsCYrhi9ZuptIbRPrGDODCm3OyxQAPnKdshjR+qtu5WPwVWTVfKASFXHkGliKdQxY0H3N4JF
BSCCGyt4cvbL7z/EOnL6x9OsVGEkmzhXQwucM3fT9hDIWUTO7BJ9SBu3yuVNsmCRbhs1SHKNgnSu
KuObvKvSfHfmEkZFrubnWVLxNKrvzEJ1oJXydJauFigvujBh6MFYxCgp17ozOH7U9b4rClVJD257
AeETzMPYTdpzbJjyitlTUlP/YQBK766/kJpS8qs+iNlPqAgUi704E4m4Xb8MHcg5Vv/pWokdZ6Tx
t9VsoWijaUfOReRndZhl5dllr82gAbCg5rGcJgtNQJ+57j3fZ2lhbCqlgWXQvfzUhG0xOX2rxOSz
KVC5d3XkYWA8pSeDVmdWcfcpaQE0ne/NLpKwIo1OAf0jsDBdnkx3RUpB9pk4xA02XObdtmNaTxrV
NFHIQ7Q4Twm6L3NuO/q5YGJdfkMPQnH8MvhRBK4GQfby92tZ7dG7wEflgwu7eJZQGnTxD+ja7/qc
lXp21ejCw4KBW9Wb08b+iYuuM7cUuzNdxUVFd/U68/mqQwxUgsubseRxvot2bfGuqqPbVUF57y/2
q2bD9NExR6Z77C5VBLRk4AGeD98T0CO6xmbjsSv/xK3pnbktuYsWcRkJAG4ZWhg9j2sU3lq02YWq
gxrZ7tbygtwrQbM9klx1oXCbPlvU8E3DpbKqsmjAam2i6U7mUNb1xT7q1IvDClenNy66MclB/+gr
UtlKuILMrRJkaN5mbdeh91ttun6yWLJLP80cBVfxtmSDFrta8F8vDGBYIn2qmHHq3sZOmPW4/XPE
G7JKSU+Xe1O6wGyo06a27qfwmkKrg5kPvIer9ZK1Zf4MfbZOFU4Uh+IK9vf9l5fj00AchdY97Frv
/oN3bkmFJ07YHtG2iSZIvsWLmda8xngVW9x2+KsuTmdxCzwdUKMCHs3Nk6GVnkYkpfOaFXblH/fx
heGIFCiF9st2tALRQXGwSlRTUo+J6fz/OWQv57gqxhVt7p784CWXV38sq8P+EzVSEafDbQrMSOmJ
JRsHrQt9/c0ThX2iVhqrqqli6NpI0R48MK/lG/ya6rv+3ang2TuOm/HV1+1dHemU4FE4WsYAygN1
k5A4tbe7ce8V2r5cx/hqFTP5k0JM0B91V+Rj3AxQzFmO62voYOeK6j09nyq+2dg5Y72qk3ln5Nz1
MWRUUwtJGPmHr4X70mrzS1uNE02kYe1Ywn2k9jDyabPvT2eekzKiz+IMLkmciRALedx7dba397KN
VOwVZnv6JZ/Pg3zsHILs3BhFe2lOH/K22gJ7ZzHostIdaLbsNbU3t0bFxoMkVynT5GK4BYTK9AzI
YlSy0OsVOSWhThrg0m6yZMuwJZRBixi+OhUvAraSv9si+0NK6Ih+6e1vXVW8WYEhcbq1wdQGe4rZ
fwAXRr+JbdCDAaPpdujDrHkot++r45t5MadyeZgSIL4dXv7ki0SVVYzvEozckSucftQnC1WORWJC
/YapRtAQx5xUKCtfGPOrAlY5tC/cEmFkQbu9M+vUVnUMn2T9kJVRWFhJMcje+sq+tNfDW+2/JNpk
rApWRlSndB/Nui+HXOV4RLebMnJCj8iZzCosGpAYy534UiNMcY3LNrPoa6iyhDwDffuGiPppJG0q
pUmj6fRGE7UCgyIw0h0jGDjtmf7w9CD3VGiQPqH4DEG7oQednQTSKVGTcVQGp3dzrtHarNLVraEO
5kp1Jcd5hx8RX/Of2oEFlcBUCq73VNCWMePuiEnmIq7tKLI3qHEM5TqMepP8UZvC3JyMtccCwPoi
qpjTzPgbxDCMJet4u4Zjd+v3Vr3Nh3F3mfpMYwRxVOSYLBoSeelNYTlW8gPfJFV/f1XSgWoAl++1
jqWIPscKU8faMiuEYEeqdjsjqJCqNhFd85IvdaIKYP7EsSBDybiGOs92W8SO4Oin+LVxVADc4sNW
zpaDpiFicq719UmBaMTehvqRIvGu5lGW/wf5EnlqkIMftwD46IN+b9gS2j4H3zo1gTl67IA3XEde
0/yM8RDXgZMc4Mml27xckL6GlIurQqFf129MIKKTDifPLWV3E0ktZo06XKyKJpJXCyMeirDbQKZr
V6sDx6Px4f6sqTwt1Vsz4DtpNJ/aGHcnLDmU//KR5xr/jGYDuB0IpH9Ofy4wGI8IQ3bv+HDk94ex
GhXWmaaK+SNni7G2+Es+r4UqHFjYmBus7CA47Hga7JmVyXdPyPmQ4ohOUsmL+py0gnfS2KomMN1y
kl6EuhGAbidraQR4U8mFYQbHWDV/2Tlyq7Df4sY77hQ5h0stdYK4yEoQNth2Gl1zY76jH2TS7brm
YroJ/Zyn1dqioMHSkWpBhKmZAjrCctUFs6JIcrBPkHVm233j1gLGQOdScC17MJJrkoeUEo+sigw7
vsWrxqIFhzve1lV8ICtvunYLiuyLe/HIiS6d9XFURddGLs33O+KQ/0NbSkNt3sc7zbH2E5T9C4gV
bydWi00iMEHO/cKz4j+82XWTTgb9nFx09sBZexOl69HJuKRF4XUlEEXASUMBLNGP50QX4DgFfcs8
wMtHNCLyEzmXQOqUXSX199xgLJatJX3rY/kY3u53BcuKKsVJDI5YP1Lvj62qUHlybHR81qGbWVM/
lxEAUlarG1nqKiJaXPb62mgIEsQ4XwlMe18vOg6R//QbEZER3oh3UtnVP9xns+TsiVu+ZmixZmVp
212154DbZTY6QtuOkfbTS89jDQSVAHYrtIhVE0zwhdpb5bxODllT1homWxi8Vz7dG4JZETHgaVm2
vFWRg/xMGqz06ymm7RHAzqNVR7GY9+fQvuGcJ02NnIpvGufHJfjeCgftG4XXWb6UtaQSx67cwOZR
kQc8J0JZ7Yhl7JCsDJK8XvZiJ0k842879hGJZuWrNacsl1wea1fUzf6vj6Iqif58i5j50n4zPAE3
S+SazewQsTZ5+CdpxDc77KgpOWGbKpmAtcj19n9n+327FAqJ2mRufVCgZVfGAnQLF0N8OSi172Rk
VFHv6OG/CEuYs7/B5pJQN5V7kqMsc6GAetNNKdW0V+0iLS399M3SvFWtEPHZNClgSbmfTH8x7DJF
isXXISyHFzigvj54ePhBEGei5TKx/FGBBkEpBX4abM2ef3DDPVSrYPBbTv0ugbSNzV9rrZBRHdUA
iIvJPSrxcofWMabxnK/MdpDrWbAMQSli5DsLffLx8g9OFY34UnLfluDcCQg/Lg+I1jLsMjrHCAc0
U4+4r5UME2zO1RMRnNwJSl5D9BH4eydvY4lEeyO58JnR+rUCYdckKtA09v21UfkZu4cX7NaIR243
BlrLODDrwji4aDcG2Ms64i8m1B3dEXWWJjPNcivaqIP0g1x6oR8f6krAUZ7OKYeXUT6eVxK1hGPv
D0Zko/EF3D5Gpnm857itMQZzdP0QxrAd7HlSNU56dwEaOjjrqClZIsK4cFv9IBhV52Ji9Mi1svI7
URgaZO8/Oa9SirFkm0IpLWxlK12U5w6geSfCkZ5vsWH9q59+jE+GVQpd4I9m9u1iRaOvbmoLWH6+
+sEgWsaxPqSm3s9sYFjfVOc3BVRB07lj2tlIWGg+QpwqeF4+2jVWP19Z2q6cAUGnf0aS/kDlgpbS
Hiu/why2AqAu11ZYNha0MI1wP2s3u1lzCmsI7Y7vVHdGkxHt8L2y5+HHn12LdnE6m8v6qf8vpDli
wXa8ALlstlmOMty8RnStkUnXaIS6u+sdG1yRXxEVWL8yrbLLO850QONQhvQuy1vZH++bXbzrs1xf
cg6R9SyesNh+O5jpTMB6l3g+NZhhy/Ugz1Yrp06diCeygIL+ehoQZXyfXMzUbDADJE7d6hWmdGuK
ILGzUcI2muvlslp0n76HrhE4+D5AHo1AewGjB2Oim67RrDXdkpwDgzX90iZbzhrY1xnMiozC07ie
4ii09YUqt01XyQusmMSTUVoSjvSal1PAT+GjRN/1k4KuMquNMUMlj+414gmKpWPevFvXpdE92Fv3
8zM3X2tdsFqrdTJsCdrcJ3rDW3C8o6XIVYHNCWEXIUpKQIMaVwxkw0TGgj95eYHN/TBrCgROMa6j
lcxPnz286UR8/oTzE8wzutaXc73GOwEOrEleGUOOEjFtrFk6cO1h4ib4ZIanSdBPn2qNzbBDTLUX
qhioYlhYhGPnq9YOJNPCb+PgSAxeFNMxK7ieW7usTuE+eB7HvffusUWWZqiD1fLNm5FFrxH+lvJm
BKQbQjXhIxNVdc3JiuYu8FyBK71mJjv2vjZXmCXNW9OwRurHT79D8QfrqZPc8AaTXjfUzml2H9qi
SBebDlB5f3WVUz8XtBULLtLs4f67o9BNEz2z/qy99V8OKr4qkwFjHC04gNE6UcoBYrPrFX53GfEv
D0RdYPMGenr/fDMtbbrWPzyCOBtXRq/wro7LRWcMstiPAB5GzS5cdgY6Qi/IqmWyl/14is7wNfel
a45R6SdqNUVZ63TQVUx/iIjYLyeM9YGDiXVzRsH2hL1OTb7UVB11GciJFAhF3azHFbxcxr8FaZKv
8f/l+uZJ2Je5c1Yb2LcAaR51actj8fYg13h9Dok2Poj1vahlHT61hnZw74yyt9AkQH32/JTD0olX
1V7CaUS3PVjr3HMmdDdj6bOoEmrKoVfskjCFv/NrrDAD4hZZFIhkh191uX48RSRli6gi67FOoVfI
pKautfKhL2t8e6R6cgbcf36r0gg+pH5urUQOjRt+s2o+INu/SyDdtEXEXV0tIevTUocQOOGZAxch
LMnCkpANdNAAW4nB78VdqDOHrkclNnHDP8v71m9Jr7OtdsjRR8JttMqdt/fLprhiVGCGw3JYQEck
kR3wnE024/YkOslfwoqfSivnFEaPk9mipomH14dDysOp4c7K/cUJAhTxxhbxP8OFqjcjFlLq9h3t
g13dYJn600wZyDVsdqN5Q7pIcv89cM9CWFfDRuBJoDrjcCd1hCtUGwWLhm+u2q0lu9fhLCKhADkY
oN/U0fg65ItZJ/o5E9m99z13EaGs/wr6OjcX/B9cHrV8Lyr6XwHPBx40+52WGW+1npGPPqncpQB0
IxseBOAv221fULERLH0I9OSelgx0rWWilutidUT6mbWkOe4eh5VIiEdxdARQeQgK8zBWxnT6cg1m
WRiRjV0J3vcGby+3cMQl1+KfhwIhJ5kMrmbwZPKcNQ37a08x+Vl4wcBjjvMIcy5xZDR/jBRm1q7D
7kTtt/ddEHnBFC+wdPrhEx05nE91sMc05OrFtmSgEXj/KeFIA+n/ADc7/SGOo/xyl0S9HF5Xkv3W
0DFChprAKKpnhHEoOVSb9hQoaHOxeMstTGC+kNZo/4Ljq7ktoWlW9u64Fvy25LwocrmHq4yNIudE
FqBmpzS1uScGFFnjLpMXGGDoN4XrWEm+DSlGVg9Wwxd6TrnPWjvrgrYQrA6b1WFu9O2Qq5XqAYUo
KTTa5BdmQn3y/aIrJJVZYmzq2xY6Wxx/jX7+0Q32D2xLNxDz0eGLZ5xXm53moFZmsezF9Kahysjb
ezuoh3wwY+z/nP4hruDgAE8KxMU2/7rt10mXeDeVnTMDLW+4Al00eUNxiqLkxKDFS/KAcB6JQyri
Lhbyq3npaDX5di5LF0u3qoytA0EtT01e6U1je3Z0EbuW30FQfIrtfFM5C1Ty/MrLX9NPIUIUf0XF
yLqAxPoCVymyXVskhPjxtwp+x9KnRrVh8+2goKwrhlX1WO8LwPMq3GCuRxwrfKynvAxCbgd71wGW
KY9EDwGVM/T5YSy6j0J64qa5j1ULE6VnpJqtx7Yp6hAjE0l4ir0LOKXEZYWsNaq0xaax1Os0Hyi5
gt2KmDiHloX/W8TvQ3uToRAvgHi1xDDedNAQXtpnmsbB2GWrgNE5LEnWVT6pbbpdLxkF+2RNQ/6G
N38n452LVtFGRba1bZbgApBGPUMjt+rkBHMGjYzugnaMrogzjFUK9/j5IFKSGn+WN2JELbooj7qU
QnPIZqrupf/IexVXiu6mEtQcd+kqidSHSklDkYX12pgQ3INxDR7rDtG+ALohXGEBCeOX/H/LCtwZ
IEWuNORum+196oN0GNw8KcCpmqchkvLXvoLbI9rmQNkrrOmrLlMOPXcxbql4Qjt+8r1k90ivbIyr
jKI/mQEJKcpUdnZ8HhbtIYpvZH0/sQVSE3co63W6fWqLPWPzXsUL82b9ZqJ2ha3PnYvkkioiUTDz
D4ow6CgM89W64Hpt6GyVg4P7EhSUEFlhV2PvoUUNUviIjeu4zZgWes9/TQTFMGlZbTrwSPBdSGqH
7dXsIVzcZ6w4fcqkVsvlf3sT5oFmOIPwXhAlxoq1BX3k1NAe7dX6cEqzwzq4z//zluROrhZRF/Q6
0CS3/BVclEc6KUCY20cx91//fjYUm7xhAczObswohI7f/C+MgE62S1Q1S6Z0ct5MtSFcLpk9ICB+
eyDl3Binv/95xUKTiBD2U6VW4Qr+54Nsm1q1n+iDILTb8RTuYRQ5WbALK4qwM8IVEfVHarXLYdH2
eITccmEGYnHZlbC9BVfV50ONAT8M5HtVpm0Ffi17kGSJtGfhJzC5fncLNmAISPmGNI51m0hArHL5
FsrKVoiswgAxyo6gVt75H+bAuvwjUSPODyXqirC8+DqYo54+35M+P41wa0tUkbQ6xFwWto8Gg0Dy
x7M1VDH5JA/xol/lglEhcGOxehRWDI5N5j3cGqYvHYhlG+o9RDMCnDGZRK/3VAu2y5mr3TQU27z+
skP0ROsEqzTqDMBu5TLhoTTZWGt1nWWLX5A3ODivI573Rr5uHRO/r/0b3Fg4c8mcC+HBVPZ3zQ2x
tkXSsY1MoEztHJ9l9i4Yy6tMM8qJIkR9lSLNFqmd9cFrA+3j7nj4OtrWmz1ofgh/ibu0LNzCO3yw
Q548tg89FPWqdA1hsdD5P24lZcrhQgFVnBxhr6U6hAFym7hakcp0C72WZmnxxXb1b6nI52E/4fHw
x9TDI1SjlgfJVaF/HKHro7TItsPoGARRXxtedh5w5Cj+SAjxnFUCNPTsE0x2CAU43a9MTSGn1zB8
J6f0bb49qGFA05rADQc6L+bQsag3uOUq1Y/b51Qh+2h88VIz6wO45dS8dU8er3NVHkRx7FFvc2t3
IT3aNkMi1e1d8SoDwS1M41MpV4y4UwkMKqAS+dtL1jVJi6QnBOuh09V+Y4/1B+PqO1TwevpwLHmD
Y4BJz7Hr1C+ypwYmp72YHvgs+Y6XFcjj4VuKe3me13XUpDybbZ+bxQWrzw/arVvo9ed44qtJMdbj
5wmHuIVEAojz2kY3Iv4OGk763ZIuPsZj8ldZKCwbZiw3xsL8lZ3WJzIOvNrPciGps02uLv56fPkU
em0ITKVp0yp/zB4am+N0FmBYJZjo6WjMSIoF6lQ6ueL9H8kdCgCBMPbbvSLipJ8XIIvKAh2qBvBq
5/3VipUU7xL+UiYjk7FaRWgJR0+LitVE9A6Qc/6otwo2waK3TLN46W9DrM3shLKRbh8yBewP5LZY
V8lDu+INc2S3htOCiCr1XGUZhE8uRUNLr/w14FkyyCFi8QxJM6w52XTX+N6Ddc4WWIf3HuuBXvHL
bNomCewvuLyhkucRfjFFYN41oFkFJoxyEBHsRgzQTqgmpASHEAUgDgRGcB3PDxrcRSHYEsWq3Slw
sn2T+JH/nbEsicd+Lu8aul+ALLx1l7SsniGfG1WTcTZaKip2NngcpANxDQrXsE0hnGrDh1ZyCgnl
n4/Q+WyAXzZhfua2XqB5tBFHZpNme8lzj7tcB81VQWzm5xAi06Bm1FHJXdMAiqfz2TmDLDjk/ru1
tw05YapKkwgdTkfd1tpbd/szxBr8j7reNfp6+lOioPTtTP3hJ+hMEsT2B0d3JxVoyh4Npu/CkV6E
RAD+S3WTxcsnFccUz2RiNa+bwSmoOEdU9a7h5Q7WIH8qOdL41jO9NpTlt8xkc84rz1PcSJFPniuI
+4TSkjqyNMOXJ+Qsa5kH4YOCNt5ydEztCOT6jDaOsf6wAV/GeOA3gOwJkUK8kAwjhWhzjH3eGhdA
yVOKwWsYwN84vgcbiQtV0ss0lkxQfREcwTNbpW221P6eW33hLIlNCXs8P+8BZh8jflYxSF7OsoQX
wQrUhUoQBXbBwv+eg8v3wg6AlDc5K1tzNEQCBSEsJMb452Bj/ogN/6seansSj4Qp9tNyjcWxD3i4
fLLXjI6W53EmZ5a49G+ReC4fm74kmGtaHG9jkjN6yXoZV0N0xdO1Hs7EtDenYnIPMU/5GPIIJlmS
NK2Utc/+IT7AwsmHLVLEkrPj0hMkJifzz+me0NkAilcLARfQLRKTF1Q+fKNQp3XukCsmhBkeuOKJ
WyIAxsd0DLBOT3MkrpUdNrlOPMfvD5NghbYNCY4aRm37Js+0eAwRvX1bO92JkLza0s+SwlHrKgPt
aBuHof6DgTTEJXBLhUM801L6WsEnSujiAHyZy3e2YAxjngcV+Q1AaiLUwH1E7QjqfuFftKGQXI8h
0OkefM9rrztsXLyqr19xo70Dcxtg2JOjWb95TsoO3Fod+PLzS3o1xQx+G+vxpSV9/7PATiBOnAUA
GgMjjdsTa1iv4AB2ModaK2lh48lNkYFWUNIE1lHpdhzO25R/sQAPwgfEWZidXXLIbxLeuV+wknWu
s5xe8MlIYKzPII2KVyRZKBLdgZJG0aWyBu/YV5+F5yC7YDNumc9V6hcuZe+GmXEmPr79aSsDbu9F
vKiPmHuQDSHEP0EDqXypJuR2hbkHpGwzSKv4d4pEbbaT0bUmMcEeWbf1aNo271DG+kThBx48L4q0
ZnfCxkGw8Wo3BgKadcJb07xaRL2Q/BKYdP+a8cu/HMxSFU95UYJC6KXCJHjv74w7S74L3hFXM78+
Kbo2Kg99EAGDjuJ0cmTUla3qNS23aa3Oy2eWtLY9Knwn+9l84fLgntKm1Yt1fIWSsSp/4+Tin9QK
MUZ6p2NNHvyVVz3eDCjjo1Vw1bDL3X7i8WE1LDD9Z1QDVu3DN+YDgGDW/if7dv4uYEf79KG2uYMU
GA2xlztloztciXgEErN852rIml/Abey7sfL9C/fuDFK66C/uSfV2x/tz++vHSKYmRSGmYaYyawMQ
XtV7qjYS4rSZfdzoahAdljpryPKVzEECJrIQ7cUg0GhzNZZVsOSwfHyS3mr4gA0dZGHzP4oRM88D
1ErSOsdZwEM0IZL+8LurEqVpSSFdw3HkmKd62UPex0m1jF2XEkJxvQZYZYGxafYaAvVOYwbQ32kE
FNWyRacWz5/9mKAVpP0whineMxbHJG7xUrqSOBkMLFo5C5yxcVTyNVCnGKbDEc/v4Gy2s/dwyBvX
D8DjhULi7ZQ5f3ngdU8LxCXAOQsrlsy9ybt6tXoqILEQa8FBixMN2dUV/VeMv3yPfNjB5UdlZb+w
ErWD7kjBQWHRwIfTAqUVVJCPP+X0vUSvyGo8naikSj2R6XsU+v01ceaRThz232q0+4zCw/bOGnQN
nAN+oduSnXaYkB8sF9Kiv5OGDK99MpVoAtndRHOb9pfm8cFjJObkrvzIYr7CPq/yHdr0ISt+No+e
upiB0gSNrPUzoRGMo1TKSrIMXh9HWoHAbxQPlTzmEqMxA9aJRXIw6XgV+dNCuVcDH+/1d6ISS1Q2
GEbnUJqCouXmJznnx2qRzxfZ/Vkd3QJtFCLA1/1pcXeKcQ3TjP44AMTBuLGlIATeSGUhMSChZ57Y
4lEqBWXpSN2/DvuYkQhP22DbBItdzM1pcf20Shv+5qi+wW0+nWovcd3g9dLkSJsaN3yodfoQrXUD
vFSJjy2NuPwp0lPMPb0xub6hcK6W8a2K2MgVNNCrLDQcVDnO0V/GQiUywiQ/BCoXROy5WJhRWz3z
MvV+PYjzHlAKloNO+FA6qTPz4Z19xelL/KLmgIyjpq5MThn3swBTIpKGdkFOqFppcGUY1ZB3U3Be
lXbdctBVC1OTj8YfnlRhyVRouOBs3hWJMlG1eHF6AmmPGOk0O4ZT9DfJLDC4tqGijSPW3eMcV1VQ
fJRtEzMPVTKUju5BZjOYKwjMQrXdNLjkSDLxPRxIaEvu/nvQZgoTwNOCFeSnRfKu9h8U/vD/UxI/
KUBJ37eDsgZ+Ya1ZYzDA/CLAY4iXJ0rU/peLuMeCSRzKcQp/KSy87mSFsdctGzJOu5Piv/U8GDXI
N+cABbeaxIKfjNCNHlnOq0Ak4/NiBJ7vVvGy2XzV6vUOmGUnzer3mis8H2LCQFk12lmIX6frdLir
G3c5f8DLr2cuu7rTYIZo8931CLu5CeOeCqwrmvduLXaOzMot0q/tyEV2MPNWohXrTR9hJCP1SpkK
uaueZC0QtNdnjXJq3OSjrpNOSgpycVmFUJyFVwIUOdEX6n//DyLTrcATNMlQySEfx/75Hn7xqRER
Nb5Abjz1PnHGXQPHeHhz0zrmPYIYHlT0kp1ExJDHHoRYAFB5TMzYr4Fek5GlWZvf1fsv9ZcedNQp
hm89jIsfQ9gdEboxyzcB/fQ3AS9ziFraqniuXMbKAydoCTlDlTvXLXK7SB0Ol7FhlxU0YIDHZRKP
iIQr6DZzXAdxWsfsRwSBnngHMeFfd/zP6jBsGgSp5VrIy0ilNHMY9/zvu614ayDJ0xB9+gUVuvEd
CBYnXI3Z/lrVIyGz8VvfFjEAFW3v/4Yv61IZv3UebabaaaZUXUb07zKAJpdpp8sA7arjWQhYsJWP
zwfhu8ELDIjcZb8P3K/6LZdy9od/ijdjWVqaPDDL0EIwrzs8RvcWuafw/oQhrfxFAkRw8t6Vd40g
JHsE88qaNobbkUnfc3nW6D9/uGNOjYxNejv71oB5rOYIw5IZa6rT1AxUYhUJS+UeOOgHVXSVBrsv
5CN60rd1lM+Gj0sD/0iljiPVx/Ce67jZBfIdAeHoprEgMdxLSxLkk98mfOc5+k75naFRAaLOROYf
+uHY+qfT0c+3fDAXUKo176JOWbet0oYuzrIpdee1IKEQaavpC/sQbXdZ+DLOkmW9pW7My/bXZOZ+
JVWxrmG4zB4/0pRMOevA3pr3aK0gv/O7kQjyNKyN+9Dt6swR5QcRHaeELCLrD7SAMpU3xFZgpfHh
Yk+lxZvrtk3DzxV46G5nejGu2CHmPYHTzMgthss1ENPTvMNAw5Y59wFiRfKB9AVVLbN3F1s0+SER
h37jE/pCJu3bBuk2G3WqPlsgI5EdQBJNF1icyOXXcjt1jyHLXKMABZjEUWmmGi6Qk3Ngvg0GBMke
VXRr4B/NONljc6ltes8jVkPD7uveJ8JE1x+75ySEpt26XnHHj/0850ildcwe81k0Lc1jfHR1uS7g
JNeFkBhdkODxdW27nKkpjHEqr/bZPrsJ0YXW1OYXC4KESmE+wIQI13FXT0/mmRxT/5fT55Au1Bve
VqJ6E+ioo8ZxidDWRt1fYPtyKVgFWcDEo98E64PPgnCei8O2qQRQy5ZGIAp7tbWWw4Y4ZoPETFWT
83c1O4oCcSrL/TPDWUhWvbVz63MaZfU+6NztajaBJLDWWBrrj1eE8W34mGqLImq1/ZuoNIREihq+
wRmihvKNiNltqlxWAzTybLZYWQsEgi7v5JjpkjwCb5neR5is1LNGG7gbcDJ6i2xV9Zg26nO2JDp3
cc6g2+3BFmX0gxugfBl1x1Kjq/sUWsn/GqaIo2fxEMp6cp4h2qHNWudUbdCEmeweIVJyklQldZlB
XgQyUeN2i4GxGfQVHxr016L2Z2oHG65YfMiDNUiyOSeeYgmZ6bx8YTdpICakqvcNONSs5VhW/eSh
37KM0eT5BbI/OXhxLSkyI0pQsgtOWOJXKqQZp3hjxVAckX6DEYjygTePhJyhJUEmSCNPsQRwZbkH
Z0VmKz6ULrP6wmMUyiFnMMwxIA1d34dyVv+/40fNwrP+uM+6ubv6Jj2+3pCp249TutmD2Wk+dFIQ
o0J9XXcwq3G3QEe0NzlVc0EGyaVZ9RLfdXtQ3nQeUcaDcJiB6f55+iJt72+Me4IbBwANEuj/tvBM
V9Lzq4kgyxZ3Pd6ZX3ZfwNwVakfoptGjS+v7yZOvawFBp2wKa9KRPCxOZVYVCw+VWj4vBp3vzsgl
4MiXX3/3I64KDrSyIZ/ilxiFnzJeoBZ8oyJIEYABpGwxSaM/HVuvbKJNAHF/ZNVtmp4rcQqvpvoH
NPTka/mmvnHm0PskZ8zlMIoQDs7wO/x6pstCHKTCLQTGAqIbPbCqwSYZsJnHEAhUnNixbhmn7uly
fa/fJPTzCZ+WU9JxF5j2N3etvKFFC0GBiANLFh1Izh+dmUVtwgyFjzrD3kxOszB3fmiDTKzbouQc
SHEqEBCxumfsDgTAJvS4OQ4Q/MghwQg4+ClkF1pTXATR5rFvkHENfQYMoGlLqcHEK8l3EKAOXgU0
2e/zG8U8UU6BspikPqqoOYl0ef8ZZYV5PjP/UgdbygJ1MqHUudmAONVG6IsSgvWLKgkR5SD2Pd1U
ImNS3mUX4c0zSeWNIl4uL7xHMMJkIafrPFWAdqHz4FDZCQWbwjsT76jd8xxs8iT7gEdOMjIHeirp
u+fgFRGyR5ZzfY4YomzjMOb46OFyBcTXchHz2uWKy4ZK+jichp5GWlmzFG9SdhRUCAkRfj3rHeEW
/PYomjYIGXIm8ZUbPXoTPmdEcSAOiaFgT56sV4qtamtvMPsGK0kzsFz+VxX4iKSNkzMxEB4VHayJ
/dxgAQ4Rpeh1KqpqQ0SvttmXHlux77zGUWBrucYCPGbnhrEkGxRLLXy6et9wwB9BjcZ9+mShDAz1
AWW8YxH1nMTNWAlT+YnDPM0K6YAlZR9FaNbZoZ36UbdPUzd8A4xyw/v1E8UWVSvokFXchtkdvVQB
71rIGVIBSiSuXyNtPjjQdEORFiflrxgo2+E6sYPXS3RiHlbSpdARV03HpISx9CqFSjVTno/O0uDk
j4kpUXxk88drCKLV5jVQkeGPorJiqXUD7h3h+z7SXUrKf0Vsfb5r+M2BrfK9ZUnmWGCTFNM8sfB/
CdQt99OhV/xG3fkx7QVmLYw+dqoPEPQNalzdfehfhvChH4kb3kr+cudJOHsLeTucBB56ujFx7+/+
HbzvODWGAnQIvk4kBZ8WcAaByc7UCFf8umlMrkMHSHi6OOwF0qbOgyJnuuop8qKhUPne2dgx1jg6
TnZTX4Rh2OkgvZQ683emnv524ZkWpSiy3oWyIGQ+xgdpnMCFVz22JRex/FpX3gxkrEg0nU0yXT/I
Kz9Al+yFd4aOyV0AJHvlcfKX0RCY7Cy5mHI9LC+D5mABLi8KhgKgpf7WwpE7mE2SWuD6VWrPKU3V
ZUW2OzbiRhDZ9fVtZjr3CTNHjq/Im/PfmzVGbdIeSALAJlkeyGbr5a9KlCHiSe+ReXUZiyfIFZEZ
DcK0DYT4j/U7C/U4S17LaILpCwMhum8DWVtwSxXz6xih+7gaAeQq6/1SAl8KvlsVdo62MAGUpklK
2H6zYchoJeEB8ogD6Qc2AWGs41bRoZeEPL34g1nII6vebG1Ge3KNPl8x/7ZRmOz2S2kGWmQSgIV/
0MQM8luD0Zn+lTPLY3c+5GanCl2gcgk56SXE3hob2Rvtzw3xLWyW+L3p8yBVfKOCJJ8yEvGtKWKo
eK7A0eFtNkuxBSJ+uJD3mow7GZI61N12KHyu+IuqeiQZexxp7L7i7qJrMBG+kbrriON3AzrwfSHX
d1m8L3dmUbz6JtLwpyOV8yGax9kgOtO7wSmZQX1lheyGq5dpHrbUWgvAmVFF8pfIJiP2Z2JGDzbQ
TbQWTaZpPIFknD0AObBYpRYvc8VI5aOdPxeLYqEGbGFNwM+ITUE+fgutWs38+sgzJT1CKKEMcNam
N5LKtlnOLaqjHhMztJLINOlBN1LocW1dohva5Kdk4vbeo0+QoXreWhcUPtm192AZ9z/7YNZr4fx4
XwCQwbWZvT16702j2ETWquA41lTWwheMRcihw64drwPmQUDq7P7rLVptiL5IZxxrlt89k7CoBFmI
MFnH5AxbJxres7UXR0uiuKJcBk1oyMoC71OUX8Dk4KpDc+bCaSAXhgozJDtr7M9EoVeQ4jH04/yY
B0iz4r38EAWAi98bZUlaJuqkSoIXtxWtIfU2ICZ2WflLHkDUhvL/AXrHIfRYD9UWFOfECJT+eu4t
vcIidl3Lq3YGj12lUucYAD25w6MefyBW3YYdkCTwDUdbQ8spId3IhdH4VW6kqkW2acF6e76oTfOq
IEYDkEXX0L2hbLF0RYuH0l2WQnjUr7rPELDiHqL7r8TZx2B75i4qgOynuUOUfruQDlrw0QytYokI
nyOIQWOS4oqmnPesQ+uTcOkzwQ0VC+qZ24+rlw2hiQI/iKQEqbljZA15IXbzd0K/6vV1piCyCObc
OKMJ/FrEJueYF0/wxZCfItg3bGnWBNxVWUWQ8EOEwIz9cCATdpkhlcIVcog1PvqZTRh/aZR3SGtR
u6iRHHgiWVDNIE/4+BaGmw3ObdzB0FMifcNcwW/5NZLpZxwK49MSulJW6dHxhRm/H6PmpqM5fSI9
OZW3S0unHtbDFCun7FzSXNjTWeXKU4tGJjM5xcQhmtlcm9eAwP0ZZSOKGg5tKGOrXTLLEmut6fne
D+mwEYlZeaKwdBYXxx+7UmrBE6KuMt+89eHbXEza/Ms7dWGzmQzmd5l8nKeDM0dL2ByB6mOaoTsd
j81voS9iueieZw3Bb1aAvG+nr/Q4cWmskQd1SLsD6isUxSDahyFSUtQjC2YTOXNifzbiVnFT5pQD
8dHVmyq+z9NYd1UZG5+PHgdVm/eK90ogwe2LTHOklW7VlyENfBXk1en+i9/hqcRqlz54eBMpcBAR
oHFtLvTt7Xy3Au+CpNgnoiiJRPRi1oEKOH5P+X5oNrGCrvAbMauJ78aHD0q9G5EkUBA63bAiMnqY
U6qMi5S0NOHNdqh1zkAd0TQIVHkmgki5qjP3AI2IuzfGjlnoYQ2Fg5YXVOBR8T02LV49pb6/hLRG
IJrZsewlyzj+d8tnEWZ21MPbVODTXHhyA4Iw1MIqtnxeWHkHnlYw1sPlkZGeDNeYAxRbbBj857nE
6XSW6c5z44vXyovEvIYeCUhLmiV+udmSAyls8pgSzutoSvnyOluSP/LNaAC0FnJxV1eOXssws1j0
L+OzdpEB5O6yoa16DAr5CKlwS0vCV1I9F8kAkkeW5lR/DX4EGFx4CwNO64FSJ3tSAJRtrwHBgsDs
rfr3XShbAPUQuccF5uR5GvJknxHHwgEg0EnDMVdpuNhRXU0W+xZGBlicXZlwNvytJY+AJ6QuLnoT
hujRXu8mgAGCZa+daYjywKaKsjgMHGQaK5Phv3vKUycRBhQAg+P9Na9rRmt2xjdQpQUS/pAhsuPj
gRXrjzgUgWNN4z8qhjn0Y/cbmIIxtPu26uVar0omqOes1i7VTPgmIPSktJLNU6Xf47MadVFAM7Gx
fzuUAta2S7G9HfJmfycOAPuJa7thND6KltoH1QYlI6JzanNZhBQhSPYv0c4/OWtxYNg3Lvq1z1QK
ehHaeWPZzLcmeBFgyh8IqRJKwNmU71Fe08PJM1qFernKKQlaQe0/Qs3D11ljASB9byGpRkI0E39L
C32rVdcFbCsoNZB0sZa20CWhh4gndTXbg7dGRdgOuAGBbpqi0kp2RZNSJENmgz71QpVnS62EbFo0
weOPfO0eQQ4DrvWVzf3xQXqCU9WH5wulc1ROahYlcLZ0Mp9AbImujz0pxByEqDvVtSiSz7UWD7HC
cn5X+PvjVX7ZFWBGcMtsYyG1sbLQCthw89SC0dOW/3wKANPO7hV/2xvshhjKJEmEaLlHCSZuTG6m
5F7Vy5TS0rYdUaiUrBn6+GjDaO6Df21wz17QgXQnL3/dPghH+vSmrkfk3VJ/0PuXD0rk83DrvKQv
7I7qpOoCcoLX11b6Iw7D+VbNxUilEuJGnbG2BK5ZhohK4DTpHaXUd/x30irx3uj8/k/s+0xxAAdk
9quNkAwt2ytu2HkUX/S2tW+sIg4rJ5AZjrutfvnA7dH4FwqEMA9DvZscj3COWuZ9DifBuVr16eaD
WdKuUG/O84jSn9OSQolONkC8r50Z1BWUs1VB6btK0c6CaQo7DZWzYiOP5oec8Z5Pf+vhqEM4P3YB
Hk5DHi2rb/JMPwTxQCmc2qvN9CmzhNk+5P+Xs4DYHphL5gFw9Mkl7VPoSVXCXHiIdb4DSnwzX7Kg
IvCsXJYrGgHa1dZoA318/gsP1QoniMvRQZIdqotCzDgC5geJsAee+AcGK/cqdacVEkmxFgekcrRq
mYo2XDeHBDq0e5vqHwvGY1Dm3xQc5K3RQxx8F6mRXE/aiMfWhzGAtFKOlB4BSOHaBNhFNd204yfI
0fRUUQyRJ9jBxLcN9rD9yIDOSHJ8m7vAq3smeJUmp0JJsHVd3hKpH8ZAU3kxjo8MdoJuF99VCCOa
NN5aMnmVuNMTZzSl2ZTt9HIBqYNLJs89Y6qFfzZPs9wDovhXrDDfuELFHepS0k4QRAc0O1y7eSjc
X+pP8npFvPsIOyVxHx2u7o/gm1N5BcKSPFoK1s/FWDpKK4aDLr8ruH5+0QQd4qvFsgE3HcrCdmY1
Kbkc3Nf1KoDdmiP+HXJwIQ7GR9nLkOsFZjYkNtXJgcw4IBoKZOrS2a2ZMhJ/Ree/qQZirouKPHDD
bL14QtJJ7DGPq7n98sOOlrqDpDdiHl5cyc4C07WDl1nDaAIqIRbr6VRgADym9NSsP/QzgJhFYng7
1VAImiHm+xZieibGLhICl9EsMbpuvgdpXNxmhu4hfTDhXNiELFUX43bKcGXxFPBU3LGdEiEBaQ5Y
VkDBR8ARvDBhjmJn7kRrzCpqxkJ97o949d1rcLLSY0LDZNn2UuRLVRyT0jQWh/r/TI2DYTXY8OHo
G2NWfsq74qWH1JpgsSDxJ7RWeV6TOi25DwivTFzi2yErlU01mMwM/XcFXFEtaukn8LocbYR8Ia0/
bhZ68bsdYJAH/5wTjDQSyGU8O1hYTcREfDL4unhHB+srZ/F+1PgrC6INZnQ8SiBW3ZRpgWaCV1md
mrhVyilZ/SAji6cDIULdbvww/adXBLXq4wwS2gqp7hdbV/JbfZIooJAbi4mYix4q6fEmWas1h0nU
KIMOrh581/q7GWvDeG2AIcDf0U+1ngrmyLYMt4R2VoAL0z3GUQTF1DEUywDkT16G0p7Y43jGTjXz
/WpNYmL3Xk78uzAoFBqRrYAhur1M8Ofdt1kPtQ/0BGOguoii55VIv98m9bLKQ7w9KMxLZxyrDmY9
tO6Fx9rKsnlWRaduCxCfIt1krJhr1go8MU67w7KvoSUlS50qmQ6Sq+A5reDqwrmS4oGVxt7dCG4v
fIKclv/4N+L/5+y0LNdD6XQY6d8NmBLBoZxUIt5qUI6WkQLwmhBwoDgHClCirQzdYwdEQNu+1Jki
3tBT6V8UvkNbb5m+Tpy38EhK2eKlpwmFhZ3i6hWc05CdOhZgIqfoqgvxlUkp6jhR6vyl4CjIWUwK
+B76eVqw/MKw5+U08ozzA5VdVg4hKp423rz03A/j3B5s0MGBqJl5zIr/HDvuaa5yZCinaquE2c4D
wNWAF56/VPXjgcKkuohmkzHQlgvuHFQEB+JkbZrakT8j24wmcWLgV24oePdEdZ2ZickDU1QAOp/O
1dKlKF44mM072LVgKZtkHhOS7U+CBY++zFLpk8bk+i47ixwUMlqL1APy1AmBkDeW6N2EmbbwqAI7
YuCI+vlI057mPhOmd4k2cyKes8ZSB9OrgqYQk0eoAjmhV29FiM/t7U2g4uhHA+xDeFMv9ELEnO1V
4iws6ddeTb8T2pgUVOG5W0zVdwE7W1qXl5zQEUK5xv4y6rnShXSTOstE3N04mawLuN0zrgMT3493
fhuoOhFzc2v3QybpnRXL5VDlDApEfLuBXOhy1awZ0XF/qu00IN3e349a/Anh1h9SGGnZElRIIMBE
Bz2zW4QugKSDvq0PhjuDhnuDkHVN4kdE/2kmNKkqavzVYCNV4kk94hVAvWxQ12PRbDierjsZO/hQ
Grbdc9h3CgqotBMC8GmCE/ESpwxhxomsHHVQ8lZOv8GvIVZBU79I7r+v/aRFFMliz1/3Ur+8zO+t
UEgb1D/YyORqhBlMcSo6hRwRrYzxmSYG0I7sR/rgCNT9YjG7UqqcWTAmeNjFfjNjNfpgn9sLpZ8R
GiF2ZoKu7YSiQItYGCyNbCDDcvAkILulXrHhH3vWYRvcZKg4EaXikzApgBYnWXFdJ42vdRRKMdik
f66t0GJ6WyDSfrv3PKuF5mc/5nM5W9toMlPZMBaPyau1nE8Ns1EaV5rt8LT8rPPacpFs5KJIzCbe
sc5SC9XtGBFeB4Ugyia4lg8dALyb761Tpi3P0baze+cjPq3RP9o+6iRzIaUoQs9/rfjHn8hFIihU
zHN0qJ3bw6HgbsTUdTZHtC4+G/1kajp6SChaGhpTN7liFA44+Ovb9YRhVKf6nZG4nMv7fhBUricW
g/npByDv9yCYsqShkRAlRLtIZcijKJZoHhuuut09HsiRj4XRiIf03OH7+0MuwABBXPhc4AzJiQBo
UR9W9tI/8uT8bNKRyVvGF77CfGmLGBfgrcs6iX9tMGPoc+3Vfj9l3lSpqiewauvheAup14zGQOiy
U56I0CAgsY9vqicMkSsb/hOE7yrp5C0PIzuJRDwarQS6DMedTAT7uGuiQRC2m+Hbx9t5UEOBd20s
RS+zIMUEscUG2r+1izRqK4Z615g0XiBN/4ks8xG7qvnX+w2hody53o9/0Q1n9sBiR0ZqE4MDN/iY
HSYZmypw92M1fLpbIgdcnHBI+aPdnvEZhhKW2Ft8tdObtgNnsyyxm51WVb9xYyRXtMwlBQpFJrMu
CiI079/jQkWZX50JbAXpe5ZS/tof2tgoA15Ali2nm7nKK4F5GipuF2WeeKJNXfTennuoKw9mSJvB
I4scE/HRRyI3IgM7kHC7pdgl7KRgRmFE8IskKSlbQLhVP3ySqtqsdIpyMKHHDEvd7lv469RltJTz
hdubGXKBCSO442bhZXW/lKlnE7mFY/SQyZFjh48yEL6ezmiZ/gIf5KktHgLrZ80RIKk8JqtIjv3F
HlsiB0FmXUr0JUhBB3l2qRoOezG2vxLpxqgwUepAkaib6/O1mBOvkfqRfxDn6+fTtp+0shxdpNbI
n0u+YBaK+hk/zaQHLGaNdgcZn/fvWfIWig5Jl5RKTUQQMERSes7SyedCInBzGqfbVjfxONH7FbfA
GisxcgJfUIKTzoUwovT3G7Zcbn8lfFqM/Np9cs7P4xjqPgrFRhaEU5ogdYtzmFoKNdPllUBrOuPk
r9JA8K02cymne32CQxw6hvCANGUnqwO/YcrRDOcHfWAztbgumwUoIH4ZVOIdzoaOTlFsn0DgXz8o
s1cD0HEp8G/7b7e2yX9UQTCkFzpQQzfqudm8Oyplp8LUtCwDF6G/JF8cLZeiTsfmnAyJZewkC1Ao
nFgZo+lHLm2pctQ/Uf/b3A0eb6/fnd/BK9b3rIIxEE8naf9PUG1XJyVhTegOYxgxx1F/Sf3+OjoR
mkn47TWd6FIvMCh0DUKHIRP/TYIoqIM7QO+3H5xqtl8XRVpNsMUNJUqcoKLtMCdzPF3Llp/vlQO6
uPpSRT3Nh6vGmClkdoh8FEdmw+3BJ7Z9OWvRw/kYJxy2ZmYTgKLdKVX6uNnLlGbTCeiqVgNPSIGS
zEpdRRQsFll88YEYU1bYuv1yW6v7GVcdtDCA4NDhXB/P0/XYQNf3yvtRBJDbmt3RKN1etlo45Vsj
Cll2W8nQJ4dKWdoMjZ6+CYKgi4pXLzxzZrkXbDKVksEHAqLn5WD7ZrGy2/tvHAHPzPEbLGsf/I6g
POKiG/ATjpG0Fm0sfCLP7YK3QU97giZzGFVm1Fqes2vIXjBDVY0bbl40hE1HEc1YbxYD3VS1+8pJ
r8BloNYxtjESMB7gRaNgACuySYWSfIqr91Cm0eZCUY4yHzponncL8HkJmypCMfwxgW6O6O3lE0Xp
V5/IlqOcGBz1b3UowZdsplkAj+Q1gIv9PUa7XGg95voH868fXJDQxfgfemE5mNxN3HqysZh2Bf2T
u4jZ5PkuqXd8vV77HfZ9eYbbTOZNNaNAA+XI5Wa403L0nx2rA6wVcFwKL6YzZ/Zp5gAkz8o7XHi1
b1eFE+wPUUhVD/owHdVT539wDsqXf42OnTVtZbi8SwfDwLg0e5cwFyrdx8HC556+QTF9cNkwOAud
qlOkP6SIPprHAOkfGnibB8MF2GGiy+LKmw6L7DlHbCysdnoueUWU1Dbd7WYPDg+RKz1nC6NG5YoI
IRKWdia1PtpWOtiaAv/o2kwZp+kQJkRAoZNRtJ2a7cVx9lMsihtGQvYMViGvwiQETXZ/uFIVFX+F
+9hzN2LT886J+K2E+6KH69j9K8SFkNAbKIhStcsJoXGgNiAIXMQoetBU+zjJMG+sDjsytjgUuAd0
DYcM4EM81nk7Bk4rjS6vJgnDHlRCsnEGzuQ3lGdLXzolcoe731KpezYKo30jcjwGs177FtbO3Pxd
BHimBYZBIifrMduRFTstDbnCjl0g262mzUeHLaR/hf/Y1c9P5OFTxeWXoihsLHbWd2rKW5sXouuR
yVzYbGhBbxDgCPulVUqMLxoujindQUkR3Ph4C+scryX7cn5GsXwXvQ/zUPmUiGIrM2kp0m5e4xlV
jsUGF+zkJUuNLcyvwvK7m/PaY1quS0/SIe9b061t1XZU0gwCewqlPvhYEf5q2ziue2JUmysHKJLw
yl9NbN4dGwOfa6CTpYJiqkSVm+8CVzU+Kc9prWSQGZ0ubGjARGYgl2o1BDuIjJpF6pXduJiZNQwd
V+LY13fqSIgzgr7OwxoUQ5It0dUz0Mq37P4Jlm8+TKf5bYw+lQQQISJDMfNcIy8O5rQiLJX20A1I
gRea1/qpoksWTYA8ZEofglDqUIdNs8gTSK8IzFrU1TF0eQrzMN8V8TizLcQwaS29N2H/LYYh5QnR
1DwM5G+7YoeU2iNAM9hAANntXPbbHbwq3kfu8sLBAsu0sp/2V4W9ex23lAvRXTrhMr9cW7hDHlxy
MzlqOe1+enZbv0GPImr+FlItp1OW2dy5XB++y89NP/cax8gZ8myup81mI/q/8kihRXw5iJ1z9kXt
Kx8xtPVrwWDUnhF9vYoSXex+wg2ikZlulrMm/AMc1xJEdHH6FhPn2XjgaHG+ELwzYOyEJXyGxuJ2
nTWwVBEuJ9O5stUH7JgBUGnUJFaI9DNyCBsGjGA6sVAv0wZesFDsJYWIXtHKVk9AxUaGSTLNPn0+
q7i6ZuqDtts7II0rgDiMSBGTPVkTwcP06QUfwTxBRvGJD/brPgKHE6yv6/lvfmftBku46sB2Y2/U
xeANAz4mzgK9Bykbomo9dXv2/sZAx1/ANvsnn1jQk1hJb++EAKJ82U9DJiyFpzWeVaWXkZfiR4T8
6BINr50duVDVFyZHOQzoDx+pu7Ra8zPBqCI7z7wFO8S9+NBrc5wVtv4Cyn2n98JCZ/AoRSN3f/pa
8jIYa+R0Cgqlo3ZXLiBBqfmJJyUPV2znngf5+/J4/m23JjeHXY6KFiwK/4q8fIIfitfmBHWxmivs
LZrbkD+LcXLEeuGVQtir0JU76DfhUmhkzurKaFfRRLAa+2WyfaGbft95ZfYL8s5/s6Dyb0zpHf0y
GmGODGpALJqvW53nQbHbnYkJCWSF+ZR7ekO5aHUJlfueDCO7DWuDZfOKdtSkDQAZD8PuPOmIcqZU
1mzSQv7T3kSBX07mKML3snzKQcqLCRTDNwTRYPlgusTfl232ebi7lEvTCn1feqz1J1GAj0eilZMa
vEStVL0JEz6wm3Y7kDk7+08U7t0ff2XNeVNQ7NxvnM2B6B/G9pY8Bu5cjdveBEIdD3B0jBS6W7gY
XYwtw0TvmyjrdKU+nghqHRBtFgAvs44BatyYFNnJI35P/DxkkZ1+dhm9ud/7I7skEmCPqjnqETDh
RNPL+Ks2roF8jMtURJLFzZsO8ecMIlnRQnMCNsTnWD7QlKSJTnqzyyslMWMSsca7gIo8bbcJ7SZf
2IU9tzKXvv8ZMHD7TB6I5HNfORJI8G2BXFVrYf81c2OaaFg8Tn2efP+LYFtHg7ZMYugp7Qo9zFEE
pP1Z12NZQ3LNpgERzXzskWvSXDx1/7EXOJVNVyioYkmJ48Y7Bsic/Pr5wllfMW31LLy6A/76vbg4
dvWaNFTrS/ao2h77MgorGHk+1I1b3McDQqcqOb54IUG7XnklxykDRusGSRw4XKNL9DlXyrKy4Qln
ZHkCjmuF0rjJrlKMJBLsdjITdKbFDdOZE+EokVVbsM5n4MsMeKdhfuqcILZZ6ZddLGd1iT9guIP9
mVQxTnmRh8TM/ugAQj7i9moXoaBfRsjks/h+xiOIF1N6uKEj8Ons8koLK+s0bMLMI6L4+sbQya0k
EdbO+kFgkwQohzqpmLUaKsGCQp887Ghz12aKOMQmFcsCkHSVkzCnnr4rN6eqaQ3BtXIavwe0yHaP
Qu4fVyv27QYVqfJec+GcX9j+9Hu9jHngqDckHrgayk/iFBgv5BvnNLhcsD6uPw+kz5StTmsQMqBP
kO67SGO8ULsGdQisjsQ579msu7hYYB4/opiC9hfszFQqQaZN0uzp7f4sRAVTiJVJFN3VOPF3jKhq
XlwtPniOCBWv2W146QZa3Lcw3VRHGDXpEX1BygvFXx8+O55THTwKgkvZo/OduUeWENn7cVEs1HAW
ILtw5WoDz17DYVQ3zm4rXfSRhu9qttEo3qH9f7uXmUUig/z+IgJo9bzCjVFB8oD7ALlDdyvzoCAa
AnLBTDYXJv6IB2NaC6nbwoe9HovfmQO1X++VK8L7SpafAz8qXhXFrvIqgdPfdFkX1ptv3O0Mrv6y
BeEObiqo4APDNrQrcVcuTqfERCBfHL3Fk/k8tFgt8MQuP074hwroCvUvZnnGWF+yvlLGFwWG9bUo
Tw61IvQKPTdrx+fHCwwNZvNp2ZhC3+I9/m+AsTTiTBFrKr8VA+WdiyBgGQMNZ/woE+y9pFRj9I9a
1uFxObr56DFhS170Gh2ZZsazy0tmVf25zF7djfAwHCSByVMt9kfdwcA7PAxT+Cpu8ZHxd/bTXD7u
hkP5Hdl/L8FQM/rS2crVmVC19vK8ZqjxffQfVpaM9b3itliph790cFuAwIuIVJM4PJgPCWVhsPCO
v5xk9zCTpR78fQJlQJiXpVQ9d3xL/E7nlfWmPCWnCDhxkMbp3fnBUkTbTHm9VMJGKVwkAkV7fTP2
+6U4x1OjAYYN/Iirx08QqEpp18NNO+6jFNjPnLVeBk2VEd9KUA3LW+4SqDKUCM/vbUth/CoDXmY0
kBN5X9bydDzTL45GtYQaGEyWx5FwyPl6rZ2JK4XcMZ0LkxP2eWYps0CZP91yNFdrpoBePH48ZOrv
+NFVMlbTZNPFZAdKFPfwm44b45fNugEVHlHVKsgR0HLtCf5tBiQRDMYEJTO26Z9xLc1SFTY97tMr
iB7unzLQei0owxKjuMfZ7cTjrBvn2o1CbmUCvn1Pm2t6pAnsj8wa9IL6AOpUrsmcQWElrc6JdLId
Gv4h2VVTG+iCx9B0CriC9X7GTiOdr6rl+9vzqpVETS3wO7YQmJP6bGEsMkJfDijKdqc/dM5iaxa3
LVp/JIsjXuD5YjsDZBn4Ni9ZlIRVEuletERb3xNbgcYDAblPiFRo5iqoEbiKku/81cTo0KPAqOn3
HmsJYJqq7RlAxzk8C5vAEas05UkDQUs17PabEZTsaOCCULkxFaFydE6QIdrTSgVYLCbwI+/L8Zzm
OLR/L3qAV04azsciXgp8jvE3JTKa8TiT1TO1X9I2qsjzYS4tLEaitnRxxo/LAiujrwBHxNTMjbUx
tjaiykj2ze1MVF6eixbcqUn0yIvd+bo7klSftHsBpUvC4XWm4IIm7ZCnUKwVExOnIp7aiYMx6Kbb
K1op5JxNdhiRjvu5m8KrV2rHnvbpJc5fQFM6YLKmvnevdobcUC6/nMEG6xrAghxSD3C5secNq01D
Cy2HQ8lr5/CqReNmDwk0A+RKo7G0aim6y+0n940k9JtueIcErv4BmviV7Lf0zkyBOfjj3VD7y82h
pE4YvVXaF0RNlT7rg8cVXAP9vtkW3KmXaG0hZQD1ANtU5ZwCcjxKxp8iBikuuvidqKzj4mqj95a4
RVgTxTJe4bcyj/GY9LuDiZO4JKABpo+/c+Auj4e2CGCwS4yGf+K+PQjU3c+fr4PDjNCfEaDr3Rs/
rckv0GDjbgbpzLsv/pXqgl2MebO7O75Ap0WVEafwh4KTwiPTYK8ytmbhshHtbHnXbWZbMHyWt9eA
Tj3axqDFg/WtJaXAiXtrmbFzD5gFBS5zBj7PacKPO08g0IanA6SMShA2/p+vWolGLGRCQ+UAzv3j
cYi+02yUR1wb3v9WJ7BK4BQFcuXTjCxgy1oAL8YKr1AC1BWvOiKuKLTlNA7EaHTzCNugDhl3MfW5
c+RNs54Pc9CeVw6SbrqGn8IEz0j5NlgXU79yWNVOtLiEU3NHSWdgBQazpNrFTBMcC8L+dxX73twi
oICcjuTgefr7GgU2vD21N1+3puZI8QPPL819x+iNA9nFIWJ4yg4MiHiC6qAg7kRE+mg3mEgKKbK7
cKtqqkwN6Q8vCKH3Q/Z9xmbpft8JL1h/qMQbhEzlEk0StEJYXmdruBqt8FadxsO1prHx7GfgcTPN
rNkDdoT7hSLMR+Fql8NbgAED35FDnLGxzddyolxVdLIou6+MUvCVrbiEytEgvui0l6h4dADhlNU6
BXssi1ik8pcn8CGu9Z5UdKd5UtVLDnbGchpn/sg7w/v3wuPDn27e3yon/zeWql8foUo76QcBFrPf
hzaBZu91WZdI67Ie5+a8qIuH2rA4s2lKo9jsck+OOwiYK9yT92QVmj1leiIuhKFOTjgumRfG8WE+
6KDTgynRMLtLN8aUnOA+Up69iIKAL7/pb0dgmBmpwxxzDr99WB+TW8k1+o30EXV7REstcundZw0B
r++ag1M5JHRu9zBkCfl35PZdb3Uf0EGzHqrUrK8JddP20Y4FladgJvNMWJhQSyfIXpJC3E4Pzp2d
Ok6f9HHQykDbnRUu0a3iPUMEWMI1FJW7aQ3AeBTUbysTtu30h9HwpvoqC8IsWMaWzyHhHHV933AV
phK14Dg6oHYPCt1A1J6Gy/b4NRJ6G93IZfoeexBxh21mKNTFabrsA/c74tkpFUpJibj6BLU50hfs
XjVQCKWfkMsjig8pu4UhF5fIvFzFmF1J9rLeJoyZVqdjlWYcW5kn9CRB/k784b7R+sJfMxeseWv5
M0//x9YUjsoVxBO8WFt4VI+hr+dVI2M0M2qrlrpsv/o6pWHsgnVZ972cEwADuyKClJy++Xg3HQII
pcaCoST9frAIRpvKzPOhWd+SVOnbo8VVHqlPKXa8ED8saUdnJoyFnUQdSE+VsOP0ShrdHfLd2YUt
YjH88sr0/49WGr1jNcnPwgu6DTOgqUlSFVADuKkLqgwOTa1uH11VCcVJS8TEKjOxcTAHpqMZqblR
nN57UPVEEhQbkGDTdLTTxMfho6rvFXoYH07fiJATTN848/KFtw272YBqw3M2k23nv1yk7i+3WBIU
62WN2FtvgsDgMzUD7pQ0OIEgPB6xi1pTzk1wW63/Gx7ChpkFHYWD7GV09fL1s2OtyCYXZVc+vyt3
FtF7ABtlq0fjyXFhvnf9xHqos33NhnwmZyHSZsfEc008/RELmAzCwijiav6B8TG2EPLrknQ8PIRO
PFfbqBVUL1aMy1WqXg5hkHtz8+uoByRgBZdAcZbSfFi0dV4ufhULb+UQcPzqNSIlEsFJyZA8GnHo
SPGCR5demMlXM24/IIPkJhoiK6vq4a5bDY2IG8qzAJitXGkDK97RbI+BfF7YmXmRoaCQuchEz34f
VKmZN1OSQEecFGr6ckgnWEckcjjPTJGOJhRE9ALr/Y18sxI0pqEReRZwUSQrEvm+I0U7k1VAB2Bz
OFjdptKatny09ZvM6K1TUCfMHiSdg8Ae91pkCpP/U8hEOAlIh6qhFaxalP2x0V8zxwyj1f5W683l
3wVgjGThvg517iaPXt/u4WK6UxQ8cNNrkDjjk0jm7UYSjFjeJ3uRx/pXriae9jxeAt7B2wMiEf/n
HUxBAIbpOXRf0yETD52YQspufym84OKrBzd+oU4BdUHJ6kkOp3PrB+U0K7I/m0E3D+CNzlA1hXET
hWSSFFpw4netF1VRjwEOeooz6oTOd6t8xvN245jnLWr4xZja5mh5Mv+ll3hakOmYSJa3u6maeDcf
F1uC2h0/rKlkEeM0t/dhLB4rOtmwF8xFgrN6/WNGZFHTuPDYoBDHA7wD1BoHglxN6cxaRKQeQ+7g
M3X+X8fmEpdM2whNHeeEo2dBiRYB/VHr8cPB2aJa5Bpt7FqRo+/TF0nbSnlVaKFU7FEYLQvYcPjc
8grdLjGD+Th0mN5vuoz5OMbpEqKMxzVAqPXgl4Aj4PWauOuEnc6hVyhznpZwSuqKp7ip+p6696Cx
jA33c0cmSP4dbzIO6Yi7szFlaW+2TXyb1Xk+Kg0P8ATqLIw58XQj/faoJs+7cAYLxOZBcgGiyEpl
GG7U/Yb7ox8yL9lZ1Y89/re6kKitXgEP3VJlOJU44fRMjbxiIkmduHzMNi9VxYhzQhcr/RbNmHTT
07EjnOOIbMUb/uXo/WJvCZwb/aP1HHq6P5EkZgEvDnSYhY1KqwmFJ/+Qu3EgsgIJsHvD8JhLqCUq
kqHzOgB2ljsZ7MI3PumewzMa4Gn+DwSeJ8rL1ZNkGymDOuv7NHuIMlAMqGLZqlMA+bRBUtzSNnJt
2h7y8Zy5Op2s/aATJm34ukg2EnKQwpMSRaBJ6P+vFtiWUEjTLvVTYKQJcSuUgXgIjuvfqM7LzFP7
En1RpSy4R4mcOFa7R+lh5QgX1RWN9lct70/Dy7dPLf2QqLbycxlS2IjXlYeCtSR9gJX8FPro2YV0
9bqxC0bhWxADhNU6IdpxZZLLXJggFsNKveKvpKvnDprrN84SVVhdEgQyNEfUkapSs/tNm5WQxqNJ
J6Yz73dENWjAsMeW2jVSj0hLgkFQEfRUJY2xW8LOtx18EXlpR0k8ZPEfsckSlOjNJy/jY8TaeR0U
Gu6zMaocEmfMhD82Ov/hzLXD6vxNy6wSuAq+jauGjP4KDJ7RdBR/3K4+keDXizoJVVR14cY5gUIJ
waehrIH1fc0ipcRypEKJ0+1daYNbj3mV3KkISFkMSBUePwXsDzLiIWALkA+P0CowE7wd89SHI6RL
l20Y89b/riPI16M6zy+SJxOJyLhafzHHcr4fHRr8tTwtvzAsyokhr09EaensEG9rypYt6LMW6XDQ
gI+TlkDBQleHlKsxgs17svh3Vkt9EUuAa8mwqI0LqZsxxKOBt8aHEvDM9nCLt5s6SPTMSaXrvMEA
9XTFY/oi0/I70vTvX5+7IphWVyG/B0c8gD1ClniYT0YsfGLHr0fjrH5eqjo5EjQqOX1DJnWHVJHr
1uENfhdu1ckwksG/hjJeR7EnlMggZMSg9aibQOO7NA/TBIE2VKh6SCD3BvTzPzX1MYlyHJJ27rB9
Co6rRu1nloSsGyGlrfwILE5JgI8cTM1Ux6JTnWMCUFP7Bm6MEimt8J/ZKKsxV5E2jLtufbcl+mJa
IWrO2z0xMLNM3x0ykxHJnGBv7706VfY7onrNIUeyrMURani42C/gBFnKYeQVzGqiiT5CynLDod3y
H7a6SBnHmPu/HMQnszXHf8z3op4bWti9WmcftJfH8sFegfG00tWX4rhs5w1NB5OdITcdyOH4ibXt
uF+SHcvlx57ZnFBUsec7t+K4esAIg/qP9zQaJd7VB7fOHzeRSVUDxTQqOblp5yBrotoLocObTikW
uLqaJm5ccJz346xSucxv21bWYDoeU5tcGfpNWtKqKl2CRanv+w6Fa1nrT6SiiACF9zlvHhKGpzFp
0hvNU6+y5H16uTmz2RtZ+AKPZbWOEJOzG1P/QWRpmHphyajv3DJ6fo78Zw/07c2YFeJosDihKMhK
lJmGl1TBN+W+Tn/d91ub0XcqrBU51ajw4/MKqFYrHeOOT0Xjg8kqoCdEZZ5D/RJCF5d4PRkc61Jm
HspaI2D+8hasSW9dOsvPzM2nTnROXZwQGu/HGxsUzNdOni29sFMUsJlgx0SxDE66RjK2RKKliAt+
6ABuxrvVlT7uLc49MzYVvJd58x87dhZSWNR51lWZnTlUIrBEkktpS+ipLDw6br4xBNYscOMCy7xA
YslNPZszZwe7vMeob2G6ihw32iCV4fWLNaGNRUjjOajkLaJ3X2MpR8qfnny1FmYiIaVTnwBd67wj
WmLaR36AdXc+w/4GHTjQ9VmxLeiBVvoVOGEzw1p+IWjfr3bSjqDq6tMKXo2/huBbOmlhMj/lLlLK
w7vwH3F4F+wm3dMgm8H0Z3ErXk++TVmO8YjfQRoD5SNpdEnvYihkqwqdC0WnDKSo+WhfFtSErf90
pdL75CsQP6Rk6MSWcl7e9Vnn9CreFu388m8HZGYk7oOXAtc5zKGUdvMv3xk/ntY0Hmr+71I/QeJH
5pVcQZbR9fvihFowbz5xVmYYiB7F8i7t9mspfr0P8SRmVrHl8F4tgUoV0uppt9sEDBHjCBv76QNM
zOINDhdiRxyOpjMNVkHHrL4e8ExXif08s9k/dx5aRZdqANHEL6MqbhDiLuCg5+j+tdMGvgBZtlnT
aStI6/272bOaD8npR2VzA4cktxetjoyyiUTbeWeOp0joOdCnEuXymI97ZbdWrx8MFxPIk8lIeFcS
YLBIh/9zn99oYG4QhSq1pAepk2uVxxz2grzC2TOKHLLqtmZeVCg6A0a+LNU2n2eonoddadIyXfs0
J9aMd2cBedMVHuHa/HPvNLMRPFLEEsCAGcyiwPdN+D5ccRLrChmDBcKVpJxH6CrZ7r9rtdm7ifPa
78U4ZmywvSOsVtQzPK0ust1MubaESsC881TWxww+j0T8MkY/n1zoquXT6Hwj+ROS0SiUrFNJAz0+
7FsyXYWgqdVFrc5LOSXy1gA04z0Bi7OIzH/3lf3GPozR2LZhqdsbXbUiq1V4adtj0OJyr2+qohrq
S5fTTeEKHZ0P3Azx6pAro348JZwsc8E2cM76jB0nlsnH4p+cdubKhYyTDCuRjkB6WsIqbVWfvaSf
NrUCzTkaYT3LHEqIccTlZbsnIE1KUaFVcq0z+BfhOC+2FG6lZKfHXsc8vo3lbppb5Ke5aqAbHBFf
7h2agEhA+4bFFg6fr8XsNHfM+pOJmsAXeZa+DIuJMzwJwhgTEvAsKxyrjvGhZ5mggJzeTYkOFXCO
8m0I6LCSzjxi51pneZb8WNuVhM0OM4eZqNd+bN2IzRJIaarKXlJIs+Ay0olDJ9wHh3EfWQHw6tsa
NC8pcZT9vMC8KB5SOYuxEy9bNkBO/NSkE9VMKXmxvRCWvXzPzvmJuJM8Y0i5rXjruIBjO47isPGk
O4UQfLhHysr87A9HFlCEo/VAK5KnUyOUDkxjcbSA+Xr7ncerdtmPsMGV2Z1TZI1vCjhWreYXYB4V
z31SEYE+sF+G6aQWz+By4PaR4Ov7FZg1Lad6HWehH0oVOAxoFQoB27Go1Z/GTVz/FpG9xGCO5JgH
CI6jXFUxHd9bWKwzg5kYSNZvO/xCB/Vq82S/lpx1aiM6j83+LznYulzhVFA+O0sTzoN0dxoT3KrP
V7LwYX1rKzE3N43f8OdUisr7VQ0XH5sXrghXqmlPKyIo3Oqp4+L0XZM7zs8yed96biztHkO6Wm4x
aVV7cyfDAGBF5oB86gipgxWt8uu849M4wdTDPQv5Z8UxjHjrop3rMF0KgyoAmLaUS5tNaF7Uhwjm
o9JYzITTLCA/ZwYjZpJLaLIiiJjH7J2grBUAuqIBJ6aQ3eMNhtRZ5j5cX3puC+e8chZ8/PQskLwA
m/GNPALIUOYRqd264vrhBvUiyMqnrHGFGoHDcR5kIJUXljILJOU4HeVvW6N3h8Z1u+tlfRQjxKn+
88oc6BmOWIaHPPkh8YbWUb+YcyIKtFNjsDCQyfJ5bzkK+5J7D330VYaJEtj/4T7Una72QrlzMGoO
rS5/m7ISzW+7dpKmKINrK2n46VFrp4PIyDjfosTSI1a4X6fqRqDe0vkOWXyt5E22ko98hXcT8ckW
sU4/NcfrmkSEgkN17jM9DbNuTK+3dr8EuXFDyFKDUSgt+yJDHDkabFMDKh/Jo7qfoN7hVnkBLQ0n
YEIpLbWKxbO/5Zl120mjZ7mG/r1wgh30TDPJ1ZyLfwSaDvVeCJPDUJHUKy/R+LA/snMM4E254IPT
60fxffFZwdrA4HokRT8vRtiHoqO+S+QgPyTVrIM3V/vuVBAC9Bd9AN2xA7oHMPk8aqX2xLVnoHu7
0XZd7VeFxQ7OLqRtVhYP9ulIl+sbYy1+ZANUs7ICQ8BUvOabQn0gTzjHHQK6yWreeaBgyPIM3/9r
+zGg7p3/bNHdWf6KwDRInGrEcNmtoPFocVFmB10zFfFM9X8u4j2zRysD/jVB0bZ/PIsgJT6uv0Hs
4VO4Wsiu2ZbgFwF/5Yl6B5AT+VZFXStdtbUdMnIhha0EMx4SIQ/ygGz3IISe/hM6XLk5HgawLTAx
s1K+NYWs5U+4KcleEn3UOqZEswMeY/xVuuQcL/gKoSvlejXShnSKKHNRYDJ8oyN8DaZt6KDjagvz
adOQYK/SpYxQ8Y3mAf0r4YioE2KTDNEecAdgNX1cCYtUIwsR3/54HjC6NQkvcyrCr/WwNF1miNpk
2rvcOyqmqDuVhIepsrccBlhUz/c7NhAZClFwVmu6rtOzm1YKv4oTQr8qk10TDAgwG6QhD+I4gZ2I
MP67s6vxsIzYdJdxj6yOAjQpA/Tpswa8urxCK7VLyfoJBpA5w4UDw3s90bnNBwC3F0oOR8hhvIYJ
cQJR+dpn0mjeSYdJ/sboydAGhmGyQm2ohspRPfJmZVl2q2FQ/swTp5vAvMEI4lU0rTQjQFMYjLDK
1T8+7C+JfGfY3H8v+xe8YguuIVhXM8Hqp0EqkcEwQHzoAsGSM2g6aNqVXxvELRs1xaA/OJ0gAJNn
+ZO+ulkQ/1straEXdhCYTjjlbxYpcStdWbDXYoMtn2up1moxqXebIqooJmWS7kXhg9HroSMb4ip0
JVXrjMkEWh/eAA7aUlH0I8GHny8lebtXBjleVFbTmrlahErUPUO407mqcTmhLGmX5mrWWvrtPnAc
igLtVsM4X8N/HkSdDQ/SkeexvBgKHD5aM2rpSWlbFXlYLpVLqUDJggKglDaZVXeX/1ZvkJ3GVIoS
1Y00VUNf6L4g4oMljC7KKzHsfokGTnZ4twBk14puDSLU3Bd2DVUdDkY/VJ5ZyRWA0ZyaIAzyM0Z5
8jZNKPijum1dZYkiJVL4LK0VZ2KHDO+OSKGPpCimPFLMK91g+NnPFENY359VZKyNHQac/PhGzcai
LlW0ULqtpjptMo7CbqaaKqFSMLCWEW/cg0qP2VSt3EHUr4RN/UGrwXx+OaIVATAtM/jQwXMTfigq
B2Cl3LBVcPEoU+wMs7xN3bQCxquouw4Tz25QSM2EnfKA9V+p2YBveEvUS1JTAcf6WpTa7z6Gybh5
AE58P82ODScz/OSfiB33PcoqRJZgqbJVKeHMUFTsnJ7ieTIzMovmlujDwv8KRSp3Uk+LU3bn2UWG
DGRkUMRPlFCSUbdng5gQS+iscDcJgCFZlhAvLEUmH/rQreaCkbcdfw9eRSyc1uIJf9gCZs3M+JHJ
8WmDZOYG0+3kXtxopPRpBaMwxmheNpuMScSrW4mQZOlFP3Na92ixxCJQeeiNzfqof1H3+a4+cC9p
ERA4Yt5ZbPAPoZv89QJQQbq3YomPV0t2gahJkH6t02ORnvsDKKInlvhxnf7A/iLg4s02PBgaHhtD
9eLh8k96M/gFvXyB2j+eaiXB8JTXcgC+3jujaZ+yWkV2GZxL++rBUVT18QT1S1omz+ycsrQlvVMA
6c2+NbTTVn6pzWSLQPV/yC4j1oTYe7wAUxjWVrxSzHbtzSzziWhWqhAtFAa0T/SBfJXGkZ/3TThS
4epE9Ti6t4wIjEHxhoTaH0l57vTXsayB1WBZu7ydQx1gAaazK9bXWrSTrYAgoeZMk+hSfeqjwnz6
T/u+1WEp2FrgU/pVZzt7l2Yz/8qJWbZiCy8bxVGnFLiy/iHVisLZVaCWGGlE5vTBC0s3+zbx3sOt
KRpGl92at2czbqkJBDa7AWf4mTb7FIRRYOy3fu2R+O7Q8mat7sLZhKX7MBQdlnSjlZykYrRmkAdt
gtlDBVds/CfnAAd93sgSVb3LLP3SVC0YjS1qXXy8hkbfEL7QyYViwWvWfSALVcBG1gSMICGKMCKj
R5KJGKJCsmAPKW7+JKY8JNAjpJ4ZvlckZsyVqXMDnfxBPibBBR2DuUImW5G8LLhw+vigEz47bC+b
BPJq6Qwik0urynG0Ykg98iYokqqp5EpbmbSgxhsfjcTme42vRfElKw9AqKMOrobxxlFWi161r06X
Uf+GfDnsIYgPG8DTHA44eEcTTkmSI/c6u//cHJdMp6TpZAuK6RS5p7/Hgu6XrckrAQT5TuhXvcEm
Ta3W1DHZy4HtYbxb5XRzEh3+XLCKJ/xkSJkZoObXKWWbBH5P4YR/bQEpLgt6B0pHh1eS97Yvz3AM
6iqLc4+VmWMQ9/3ncZgx+1lSP6ZdGXq5HY1osc7gk42tlC2mCSk2bMYeUBcO+rqHdF/97TQ+8B/l
I32bv2Cbj7UoLmT38PZAdPhN5ddHzk90DfAWwohInN9Qmou8mTpmpq+OURw/DGLx9VpnhxlhJuZ3
l56j/LubrwnHvUIeN6AdK30coXha29piBE+GqECICnymmhjPbdALKbHdJCz5buRfJ0oXjP0y7RFu
yp9NuLn6jCt5HtN4usESKjrYDna23YwedXbz+v4ePaIo0Ya4ADaFx4mMEjDhWYAJe1f5VrvBXbUd
kVFqrgctCcPDUtjd6DFKV/zkGQxIhn9hQuG5yKetibEy4YsA6yC1TZjOUwk7gPNcZ+RJyfXKqMh3
DiatoOOTK521MD8OBCJg65GURO3Iazarg8Gq3zUWVJf7jy93J+LdAqgTr3tnmPA6Frgw6h6dFfv7
1TGsWEuzbWF1prQAqtgNc89VIPACKo8mvb+v7YzN7PdgYeD6F1XlwcBBbbAAT0PsGTbwKrDXDkpJ
FyNU4RzZJ/uOFy8JenFqNxa9NH2HckVy3+TE+66x+WHmQlz3HeRQWnw21Kl2Flqu+0qd/t/Nttsf
PnTzJGnjPTGT4A3dKD2FpREHVBFmT5H05MQCoGQ6Je1Vr9wXySFFOZ3jiFW6hvTtZqZ33PP34Da7
vBFE2dii/nmOqeltc9e9iUkzvaxc90A9cQ5QGNO/au4rp8pzfe+QsY8N9pidlE8Y3JxNdyl8GFiD
51Tjo/QdwxcJxa2Iwb1Elaw8DQjT1I2/bZUMo7wC4wZTaCbgg0vVpD+KNNZjvxkwcAAa3XnQyXL9
NWqw4NYLZ5ljXmbNW7QR/mLvAS1NcX308DkeqXpHjbKlgFC6vi3VDSk9WtNDJpMRY0SoH/svRxXg
qnb/K5hGjtxBjJcwERWc6EbL1q/Nxoxm5s97bjHhpmSvU8Ay4LEXxSRH5IAlDbR+LagPezy9bWtp
qHn+ExXTDPYHrCxI8gNjFdONsSR0Z4r9YtHt3Ix2g0H3kkj1fjJpLOxDoegAAS2AXBDWvgkXKn59
rHJRN5WhgsOzx6fgipf/vg1i7Eg3d+NdEsZmC2f1KcHzXk4xT/mq9H3zyvtdylGGofFFO76mET6v
Bc7V/oJosT5iDhioZtywhy/yAON3duytVL9u91lHHp9wp723YuprvRacCw5xL0ZbIVzj9KwOjXVC
tgJALXvIeRuNOb1JCDNW955WwiahvSga+8a45IZVSAzdIHEOb36BI1jcDelxn+YciEk4z6yHu3B/
UvbP0Gc5YrJdQl+FnilBbYP2ozPvgpaxDcrsImlZdE3YTwxcS4ZlazmtqIH7dDJ2XCYIfaqDN1XI
/5MSd88CuPjHUYWvRmM2R81jMkeCPtFKyYtkbotCT1AChMU+BVzbzqxf/Z00Hsb8bPE3H6J+/E4m
UgFvCAMV7MwbEI8F+IVVFQkNnKbaIo8dRRVG9U5b9/XBpAp9LBCBuo9Gmnn6kUXh6viFgFOP0Vt5
JC1pQTNbgS6EoI/evb5f9GqaDgxBklTrShGDmU+t4KHSWnky/HX4jz/PT6RucW4wrE3S6JGv3RlV
XC6qL7O2jWg6w02+5jsLPvyQF7E1h0aPZLKInNaRqObC6ETXxPaLWvYczPrhRXtP4zevVx73rnzb
eu1Bl7M6aD7s8llHIUgVMUJi0fscfmb8jOuu1K2Yh4GRfPesdpHEc69LgqQbiQdlsuAuykytMVs7
HtEwWp8BCmJmLpFsKUDCpspEKdPqEMODz3/5694M4K8Qeq8V5OpOSGc3pd+JCqmhB2X9rmXqsyEH
bGKKR7ue+gy+NBV15jTMTf213SmJVb/3Ez3OPIsw1IG6MfG1e7sz4CUXZwJd6SvaXXfMn7Y8GLab
E79ccRhAjotfeFPE/VXv82LYIwIUGYlII79/esAVQWuhaPq1aBw4PZYkffkkRVdMlO1ipbNnf7ZW
tK7z49K27+SJlqhJ0fAnQL4edsLoOEVLfP1ifS9tB6cLgyim8nJKlkyr+m95aDDY40UUQhBWNfgK
A8W5eiz3AV7Fp5cS0YJyVbuqLWHUfbzBH1CE4Co5F8SbnWayJ2Z+FDFxQ5phZxOXK625Kyjk0aFj
ILYXdtGESCIijNPshOT25WaRBXARLTr9YnQTY+x47975kUSZ+Ofa0caqCYCBQiJDqzQ8u6UqS3OP
sOh+cgUj+ltuGejHMAZKmW8OpDUeL/RNrujkRFQ3XjO7uA0HYeEHcsFMFMCBiGzDKlqBWqnXanFk
5J/9HD5LC/kvWfSdNYpB5bExKYaODFc1a+TLACQeyG+4qsuz8va1SoqebIhGpraeZnf9iLRdS2Bh
KkUUXaGWXSxEZjk3yzOaSLKS9W6RWJ5iwuxHiwZbBMMUkD1gxOA72CUaSv8KJ8hyzdhzVDfp4gBW
65PbKr0eXtYnUAgRnJBAdkP6Cgk4U38EkuWW7GMH+H011zwnUHYM0geMcSZAyXwxYlqwzaapBbm/
22GnK5VmnrKT93oxBToB/FVkgEw77xSwW9uwt+s9OwTWtsanaEghy7ZZdj70+9oDZfJdPxwLb1K1
lG2r8lwFU3cABPlbK8ZZoHDaipVLXjWjMp5W4ikp68SpO+2HhWwd5Xp6dxsq9xpMEwpL21HTwmhL
z6UChbO1yDaeBRXu+NBna902kpMEyxokTSask/RFeRF5FZo8stGGTQ5TMe89Z3sY/PH7dfvOBwav
X0lBmfCOjSduM/EslCDYhKkxQDYFCqn6K1ak+mRclllqgjxtStxtTtg1Gkxhd+7V1VSD/FQYf5sC
IbV8qb4KF2DdCzHxkLZgAQlJ/KuyS4kyjzfOREZ9sGdRzgoNGFgnRQFiuilzZvQmZz8iKX6E4ETe
2iD7oLxo7eCZ9WInLC78g7KzIINiGkxCZSaylLI6yHmXw3lBZeagfrlH4kj6FvnQG6IYzbzB+8+b
U6e2i/Jik5WEsTJL+9Px4Tkt4uKg8ALg1xf8VOLC+nQLLVnzZ7EpFZ0COK8cKqOoyW9l3O3w/Jt9
LEcdF9xXlUO5323IUJa+worPo5PxgeryZt7ZnHf9qDDg5Z3fZVUARcz82JfpIQ2ffcROmvEQOG4o
Ive0OPcXWjNoESkodfsOkGMWW9bpNGKDfHWQS4rt4efCKq3JJPsn77UgL1YAts5XLQWdeqcNNbE4
245GHBX+KH47wHdy/cN4YFVLnsoGhLOuydAhcIDpegS3PQkFzQyLwbQBnWU6UvTIsUJSlJpGgx+i
Pl8yEd//Gc7PqXmzlBBJ5LdfHOMavyeOXrQ91LHgyIvgfTLlCa8rBevpE0YmxGNK/kHUpDhBv8Jx
F29LRNOIQUqWILSnWSL4SG07IGNekguCKjFZuhXZx4MLC4o+uS3wJg2/1kjjqhnRyXTT8Uf6vj7r
vY+Wa53pkaRv4J1n/VSaB6avNtnSPl4xD6Bwbpca7O83Ifajbq5Cjhoopv++bB9ZLqrJLKITDxq1
yHb/ks3QU9x50ug9qw5QNa3TVwlqIq5dwRBNrsRQ90XxUdfNNy8y3VJ/NMfZ5sT8q7QECArG6COI
mzRLYXXJYduVqzHArSv/Zgfm8wv2GU0Zyw8IS3eVnRmmbGs5PYzh7l242yXq0XzlEJIdVgQk5Hr2
sYpWcyfi4+0YSx/KlofXNlcO5QYfzGaUcTzJbV6RL+RagWTpuFtcsLU1jeYVBrRujvnAbMyROI5s
8iwHYryEwNoVyBXqew3KTTSZRxIMP9dGlmDB/DLl2jWdUmjbfvjtwDH6ClOcuh8O2DcOov1Cg63o
/ROlecij2K8+rb8mmD9j+ZBJLjj1ZURhufiFfqx7Ik0RhlaYfMU1mx5w34WE0zByYTWbi6KhL+Oj
RwQ5d6ONCJoA5cVfUlSY+mGueTIXThZ8OLVFGoAucrdNid7lR8GcDXtgisB/joLGDiNgyoEEaY9l
/juta9hQaBtiubdfieR5sD48SM7OZbiYQEV1u3s2GbcUJzcfXSWPZ/voUMaw1V4l6pzYFD3xP7wb
9VkekCIVBw+zJjJklZKSxzXJ9d9tIcdXlud59qXWdpe05HIt3Dw5EKnBqOVhk9zHqcUEIt6ETT5l
rCNhCxgZ4n1OwIUBVNmhhwZXLMSnpYoP6FlUP6bayj8n56NBmMRAuiQpKfGXkbolFnNrWijg9sFf
xd9e7L0Dwoi3Jw+3U6xiX9y+cEsg3xm1ju5DhqTvzya50d+0vKJSyfkPUJ33rePWIVlPLXhZN0IF
w30sObl2F2B89heIqiNq1iULoZ5Kzbw0GLU0EFpYLTBU18SvPTiG1+ox5Gk9rGT1yTS7Km5S2FaA
fW3zvMf9AwDGCCXnG6QTOgJfJXnvRtOR3+5PywwuT9ycmEwnuLi6c6uF7mD+fIJYks+3sDwcprlk
njGtbaWVFOLcfBj0Z7Q7pof3GaMddkqUPFxuTK+zThX6drq5G9lR71kjcQ3xAd07Dx3tuwFQqlWX
KGdc5cQKym3TxF8Bm2R3u7a0an4m2YHK3EwrgCFq04AP3qP/+zw3VZQoMxOWLWBta4r/e7YNlxJ0
s0zA4tVMdYOYG3vQOcb5igz077pRRjqmsEBzB1S1pFSyg8z4/qq4emEUp8gKyL+lowJfaIZsTUIM
sg5jJ4Rdj83CybkZFED3pMeMuu/aMS63MO8BPaZoaZTpBjjalm7OFedzEifJQUolb88SwC10ZvJE
lrFhdpgEJ85lQ3fuRxH2L/tLMHvs51bxJd2ejBdfPFcVkp9yqGYFTbbLYLg+IX7xcDUn87D7tAwO
3Cu1STUsj/Lcpsix5npk199pHkPno824Q6QWMNUy7wLYS17VW+nqPxzfA3lyJQSbNrO9T/mkhS5z
P7uojVxcp5BBdQBJ0zPO8FVpGMhDFuEUZt4OLqzgsnDpFxds96NJ2oy0DlrAMkjaW3EOfvTr+e2D
xtZHxjpikGEpBunPXtv2TZ5LUgH/1iqhIi6+1MN16rEPnmBWSbbT9dW8HKJa2PfsA9+59ZOU8y9Z
kKglXGo9g9I2RibPKa0OfZdAwjMDsNSFM6TWxhyi27FyD7EwiI+RJvFKbyqpsbiEp3Q1AFTpQJie
VJT/obnPIDPGBqhKOAhpkB071Y15Xba2j6yGGGLzHb5e0355xNEGzSJIyoBAR3Kj2TKq3GxhkNkf
pGUMIsPTZ9b/fbPldY5t8++q4hvRzRHjyg4nwcUR+yIzal6CR1mYpiA8q2akOSVRBLlwPsOYD8Gc
cSPXbwXUeONDmtda06OtXZxTcgXUYO5BQftZyfcc2RWsy/mZ9F9K1PZ8Pt2EOJS9HUdbMf5suYqM
Qv5Zs9uCrlpJ7/Md6CHXAn6Gbe7/0OPAJKn/qmXBbWt0z6iX1tJYahbk8oDS+RIuhJjJV3HuyoHw
6mRiXmAVdzIbNHSB4fKkIQ5F3uTWhUcggMVCOPO+uCKdHKPXPK6zHtfp6jUjObSbxK2j0l+TRXRu
8zGPBJdKDUZci9Hix5ha8YPF3xCjwz+YcGKt3Tx7UF6CcobIA2cZpo1+yUxXUakyDqBGJLvuyViP
rNvudoX8vxqENFeczGPv2b/IbtSkrcj8jl8e0TiDADsXYM/m1U18mS+Uz6sbL4HOo1xwS1kHmAL4
SVzupqF6VGQuvCJz9A2QyJvNcfgwJqR24FcVCUpg3XguSkyrTkFgAuTNDW2ACMGLtWdHGTQVYiq8
ZJIq/eNnIxzafKjsNDi5ZgygtjbbosgzkKRWMVsWYuboVW74pYZwgCq1rU8TWCkbxtVKQEwFJUj2
EOEI0Z4Qnub1I+BhuBfJLTY5azhEiIetTMr0h7memjmRTvrImmFaZJg4tqqIwzW9RmHou988wyv2
O9tqd4/x8TydVjiWzKjEwTYjGSvfTKiKUMOiN4hXu6EKg0KJm3nC7vQBMZ1wkT9EwFTSAsk16EAB
EDHKSu0+sXEKw5j9QMAgFtXYVdX7zORk+Oj8WAvVZV/2dBL1v4P7/9hpM5jgE7bSblb9ow8Uel1i
bpJ8KKeJfWofVZ+gryNjsjJL+3iRp/HrttCZQyC3DS7gA0R28dRyA9U2Fz3S1SE+Jx52yXsQ6cVU
a9AxdhbzogVSDVY9B49mkvgJLpEbJtCRniISPtNdrzNef1z5kD200x/N0HBj94PVo0wL+JuAHX3l
pCmLXo1pZZ5QKwpGmlCMvOIRyVEXSib2D72yeJ33x4FGkIh6G83amCW6MBDgA1gATxw4H8luRQhk
quVrChHnzksB+wCb7CFWbDhO7gciRSAYZxWD2JCzvgRjXng+nYkgRX9ubYV//9W09aEFS7qma+HM
Y/GvCgcYSOpZVBOjrmI2HAi/Vtjs3lIFRal5mfKgN6BBTVQ8mC1iuj6QF9RyC83mDoiu2FPSbo51
Zly5Cy4aPQL3tzpg8NofItZ8LmIbFRkBn4Y2Wh2FBXnkQns+U1VT5SjbnLm9vlZpJfCa8ApOAE8+
lcGEP3ehzoinsGZuanCH1vZFzN9io3/Pmcrk0wwfGrFSZBKZydIDZM9ZlbHxSFC0xuROplYWkZLr
I38B2hA7W17lPa7jNtcsXc5Qd0JBiF+1BzHRDk7N1RAicVeKJu/nPEbzyafZLikT9CMeWEldHnUN
wVhSrArfdkv95VY4zD/sqMHoL7dJvoC+lkptVnOJeLEk2chcGj5wJSWRB8RqVP4wUy9GuT1kh8xj
pAEgv4sUDYtfA7JfZMJ/Uf0Zrh7aesVmYinn6kxjaF2XQsTWnXFbjnQghDXSVSILDKI6mJRXjTmZ
3LDvlNWGlZvEzatdiGi0ZqI8XLZpd9ZBCWCQrTVinpkofl6pwODijUL363v22qLRgzvWomZ7T6jZ
cXHGDLxgoeKyTXOj2vsp+j6ISAqPkc4ARjrU+/zJQhNtezyjstDyG+gIhPdI0Z++3eJodA/nQ7fC
EFseqpqKDPIuAwUSR6DRKIK+KkktURjxkNsq+dD0w/Q+2PlEwA0G2QnbDzNA+BWsonXi4nHceslT
YU3uvR05A1k9/w/txfTOkYb82xSN0B+iLCZyFcvoPbY1MlW2VfVi8TfSnU/AOTuyaytSFm0FwovW
BYK4x3am6EmsZ4AKmf4eq4YLQCs7ekZdoL3soWYZMVgB4McXXPTd7mf9xn2p+o4mDqqAtahwFuKW
c/zQTDUDmZfSpyteG5MMHSjAwRO9F9EAxio4TKDV2OcoyMVn+hYzLnGHbt2+gLVU8Gi1iSYkjDdF
l2a+70IpFl60hU487t9ewdBRd0C3p8ymd2r9jJ2OmWrl8R8ghfcizHi3SGUOYMhCSElXflJL3ts+
4wicDyPh0kToEBdY7N57tXzC6B9CFOHyO90HqR3HEXkBglTPNt5QII4IJMwkS4fYWsIGxq4hukm6
rj3+FblEXwbybCrMzjfqCySojzZS4QMSCo3CN6xYSh5z5bV7vQaEExi06XzX+hwesBVFOV6JsUDy
k2mVqlTWMIRr9SgUbpGocEj7yR7Qt7RwNNEfO3ynWj//IyQuwEV1XN9FML1HxT77895FM8KpMEiZ
6UvxRyII/AI5dM2Qs8ykdxy/gryuILJZNeOFIr8rP27CDd+rNYXeqEudyeG5iy42qTYmgJaMEvFk
SXgSyRXsX1u/rJmG0BHAUTNUGEFDm6h++m5MdyCJuUyKt60TaMl2IoJI1Y1imK1Ym7fN9XDSDhiX
bsu1cbrg0/2yva7TJFlEndzLTY9r3ZkA/wQ5OXBkMYz6EOR9FaYRemBkcFhyPfqSMRDru8JRDbfN
30sHbYi3HpfUo2wql5WDfBoKSuy20OWmIgRaS+ooKVBx8p1gLxqKJ2abeIJ0tMONCeYl6HdEpS1p
b6I24XCkdb2Jot0atLOxttY1OSUnrNbXn0mrl7c1BE0rBkNUznMt40m5HMdlcll2ilGc5fjQoVHg
L8KkKOSHn/JUjXfy0SK30fT4xLlXuhyIS2E27As6GZ0U3Wlj19JUX5ttxx/lZ2l/SdOP0RJVV8jf
IvCPBB2BQpOgUP6N2dDipwb3PPTdFlVU84gBysgL+E6B0TmI2509Ld1y33c+XmE6K+cNTgQ1Kf0V
q5UUduMLO8C2kpM5md5sLvSufl357eFAuB72n281lkZL4VZIq0+Ah56EHvXb7gonKcN2rdw6KFaa
ngEbMBSYXawK0ILXw3HwYlmjxJUKXyTxbyxhnZxYcEuTwjJJOhngOzZ651hr3tIfZKC36iwfQR51
sOA4Vnw9bqvUqlz/hxR4feiqTZCjYSwFI/clPqGMRSsqBUDs2I24MCJXquDBWTN6CExJ+IAxokdh
R2jBIwlaU2afnXT5P5xlodoKFmmhsWRwC0FW7UoGGHEfWxwk1ZdWwISjY/4RvMxd3vdtt5jXPtYX
Pg46I/6oltma3RU7B7oRCqHBZnjAFtrjqf7OU5ygteLna1H7ftJFgFfa6ofIhZ7M+BWey0lBqIVx
+RMW3W0IGe7BOpVRm7p6HmmLG74tJaF6vCGwvFeV6LujW+lYME7F4uFs3OfmVcZFkUkJE6m/tPxd
QtIkcDFX/rIC6KiHDYeahOVGgr5Fa3mYG7Hp2Y8pPi8DfJFv19g5eF6nUeHMD3QmhiYSVarz3R28
gjJs6e56I1Wbt2O1PVFsNpmXyNS6haKcMjwesgdy01nuApbnYOtpfgvVXzjDbc6EFghyYq/yHN47
1su/rsatvC0hZ/kooz59eJA450BMtoNSDc4T1hWqJ0Ixgcyv+NX6QslvpM6AWBFBohFi0zC8anWi
sVbCFsmgIS75FjGyNiDwCrdPpw12PWYwB6PgBjo7T5LXM2GGegrlh5Q95JJmtCsYzDrdpilCfQkH
uNoJvRdW19qB//Aucoqu8IXP7L2ni5T9ukjwe4ZTVAz85evM8j/OUtqeblOiU6SI5Q29vZSfhp+9
LwXnnjX/ChTKo9R0AN1vRPGi1e9FedZw3DGNIJuuiyaRZmWFRhOspuxQXQVD+9mgKjMTeHlMJxZq
6O206NeNGKrUeNyxgGP/cVc8JoAElIghIzduSY7jLEBuap4Goh81+HqmuQYuufFdyhPjWHqVm7xc
3EBvVzQhSRtOKWLhpinHNYNzektlIi/f85EbvJMtmi4VXjBUHzkaMj7ZcluCB8vLJ8NZnY0S/C4E
GdLrI6MjgQnE0tz3LuFpsFgNDoPaC5CyS1vUXjFcJSce6tDPMpxg+860UebMm6gbU/do8VGqa7Qq
CGVkpRbDHz3p3NegHxR4iwcLFv2QZnL5z9Sn7ez7w3EYTmLg57CpR98k1zqTq1xzILnKI80NGHjs
p87tKncbLQgCjih53+rg/T69rHgfsXYvPAcCXPrpcuycqbg0s0xiluKNHfXOfz0eHSA9BuccfjCC
zIqRQ4uhL1Yuww/SF6820WBTNZdgg0f0O64xdpjjKmKRhMEiKbsWqeb5XcRT1dPFasZbeVpETb5i
Dx+i6QgoTs6iUEKbeKEDGifzBNiQ7wvs132kVpUDUtciUS1Ht3DwZoKT44YA07UPFP6c0pwna5Qt
ow1p0esXe9wJnKnZMEvzdF4q5X6AJb5iK+OdbV9RX6HSlKm7WIL3IA02bxAzZtVs9Rq4Hv94WL3+
6g/YWaQR0Z/BWOPC2GMLtH6NiQ+dSskVq+BbyAyjKIVKqlO8xlGONZoqE6E/hJ1TcFsq3sUGSPWA
ZBq46uDDKSchLDryRtpy8lTJ9CaSzr0p5DUKELGx7g7NgtRi6UhxJll1uNQmhWT0ebYbJJtSp3Lf
tFf9Sg9KcTsP/OojnKNbnd/Y4vjATXtrdR8uH+cXr70fdmMTNfhhkoipFkq+lsWudbgKlr9YoGGc
hVuiwuSIweY4nNwSW28ABG4iGVxDDHnyi0XljQKbq5EIhNYCEUDOoZUFY9DxBTE20QSEKsV1IbRY
dlkbwNEfBHLGP6fNaBKI9nSDmNh6N8r7C5//3eI5Q3U7SZ/Kao/mK2r+bYkGHKe5aag2UsRyYrBe
1OnC/G0trYZcXhkF84+2PKyyElih5StqVU7P3dsTwQQ9DVG0KxR6hmaYIlBabMf9GRIcHVf+l/nU
jEg+XLSWVfevyAVdqaKpjiXci4Tb7fB5mn7uYhn81mW0jD9fjy9HFK+cciRBtaeJfBW3K1t8gyMw
mvGWRiquTvZQ49QkRumC4+Fap7IFD2rS2Ovs3UNyu1fgwmULjQw4iuJ3kLwvUV9KC2qtrpLBxP1+
qz3Im3PQQ1A3WLo38QZHY40Q/89VfDvFW6F0Ia9utv5MXm7pk6sQNqv3WT0yGDECIJfz9KxjXVN9
5rqoXs2lJV1m4jBlpHVga7omv/48Ek5L7yhV7N3Sc462BmwP58U08yvjUlSbo7chD8CmJdo0AR2n
PRgtXxK5SGNrbSDbfr/4hW010O8vqeergFVKEoHxU6oiUg93e4RaxQWb3nx26/S8KKgN3rRzwGQi
O79WcTGjLWkwlqMiBPGEu3paIiEVyloqwuyQfibg+YvNm7ogzciRz/FNCOAYw08Q8tAmjGtvihXy
qZVNNtnTzxN/zj3vqVCMI/B+kfa4Kus4+hG8eMwsAJcFuLecNEDB7dc2dfXqm1VfumTBpaAnJX6O
Pt42ECQfWHRacr3XUE7dBha3/jt7jg8P9rfB+s462EzRlBpxBvG0NKn+0QgIJcMhLAalsbGPTo5i
9Rr8cnAb8hJaikfeGDFd9wdAZi32SI9KwT0h9e/TRc479ZrUggPOixulAfjTse/JR5LkvKYz9WYo
s4x/G+se5iVLS34xdLUgoWDUwGPMUYtqoMUNxpgBh24dHsRbllprBJYHNeAGIPl9dQsHXATRvtrC
J1CD5RjyXtsaGI/zgO7qdPl2EQVHJTimtHGejtQB5G515I3excYkOFLxCkGlvYv+YeRPOdbNac9d
YuAemj8RM6bqbPPX4gLEPVOvULUjNERRL86Be48AsIsp7+ToW0A+3haAYAdf3hAsEVyzvkILG29J
i/qV+0NC0zejfoQ6eBBdYVr1cXnmx7/esLvlNgYxB1ftDViPjT/qyWIsqz2vWkHY9Mvim9QuIj2G
oP4v+lXu7HByBHuv231DGueD67ob7/ardJihnVMIfaPVAEGlM002/DT0Yk4RkZBuxdNCNR4l7ekO
4SUdH4wxL/BP+VEep8NBatEtN15vJ/+ToI6b/Rjvw1tXZWPh5Fu2a0IhdV2OAhS6ZKzo4v9DtwZm
M/59tsWwUUYneMIOPJ87s8fSdnGIKPAEuyhuueANfxtRuygnbKGUgYrQ4qNtGJrM3HZBSOQN2YbM
vqsXvb0nnqwcnV3GG+YEeUYqXezTTcdC9twod7+YmPSnythIvmQ05Qcw6qxRxSO7niQRwFrtUqce
kd9hUMa5pROFowKuL1yZptCl70IQzCuUEYprgeEW9m1sQZ6TMxDWM9KPGtmSMuaWBd8eaHUH9uII
xgo257TdfY5EFA7c6hAATrP4AML88Qr2nzb9M4HNWQ2HtThQa9ALH37PGOh1k3+hbbBPlzAnGqb+
MWSLJKJbApqkm17BXnDb5mqN3s2pTN63aDtMbv1NlY/EjPFKQJ4BMTJupfgifSkiZjM2w3cO2t5d
XCEfIsnG3hap58FhVV+rCy2UT6NgWLliLJCzM/bczKhjv2lsW203eem3zPY/TGnx2crAk/xikpQ+
ZbVCpd1ykZCMNA3fv4B7TPxk0o7WRBg6k6lP+OwTzSQI3bhPfVnaPqKkJcA+3KiAIKYlpjwoTkZo
O22Pesw2EB9102CaiUdcqbiykdESgtiK4PwmhkfyU8Zx00GnG7mcUbrdYf5ZR8qz+W3996RhTyOW
1wFcbFseouz0TSythgIq5vFkvgBKD5Gr9OzGWfsWS4QS5MIrXBZPOW0MXxoZEqTm+ecOgI8Fv5m0
yH/TiU+ZmGwT1Txic2ZBugQgwHsKbS4Q1I4wkqWXLgH8BLuAEmBwu/ZBhrhIHO6eIE+GU/rTubGP
D4Vz7tAeE6q8suio4uon1HC04EbmulYpwmgwPCKEWwBHkAfJGwGxczxdBXXJkLs5Vb/Ga01mfPGD
I2kqpD0uQBvHsZ/0m/5//vC+u/+hDuqUcI85pONaYw6xtWhqmSM4H12lAbTq8Y+DMLIQxXThE4eP
0am5Je7NMhOW2crFs3Xk0BTSsqb2hzT5S830LdomgmN2LFacDS5/AtHKVXCxOHPYaW2llIKTspnj
PaEigO443IFVBgkPYkEXm488lFJnLf+nMYPM2zrisTu62rEg7ENE3MgxUBW3bU7Vx/DUzdl/24JB
ZzqHdJhstNW9b7BeJC0F7LZu++H45XBoolq+yg09digmBi0y9GhQtTFQo9eluKjyWGJlTwDNwc7D
rjpz6EK/u6PA6OerWXYNwAN+OoHTFq1anG7MI4myc3SV4dO6hoPswdygKPn1Fi6F6f9jUKV9xNpB
PTl3FtzJN3nw7h5IcS/4c0RlmZ3cbqQdfdJtXRYwEMtd1SRcTJ9KcA1sybvLMfMM/gFjyfojGnXY
eSgkbx3NZQboGuGcfR2TzR745bzqJ7HJd7qb6SWC5MTc8av0L40BdBdorZVV+ESYHubDeM4dg+TB
g4Q6eFl5DGwTVbzzBfbsH9K+0SZrlYgY68OLfx8BlsDiqB3tnZHBWYbEpSSoM6RG8zQkY/jm/P74
YPfYVMAi+CdyGtpl4Po0OF+rk6nWdPouo6qm5b8dfv1+VoO49l86+2nsoHwCdxwGrw1ZsReoObsM
OSjOyVPvKZCc6kdrCjTtW4vUAzVb43tUur+xyp9wuIT0VB5h3bPz5MzNJlDbimIpgSKoFLMKyFAZ
FSp/z2jwbQgSZ9WmcTukiNypHfsVNZ3xp3dM4CldbFc2JvF10qVXhSQOrA7uorzEnfz3MMUHXokp
LjRvIhkAXE+2rG6/8pFVpA+7RtH053w21lcLEflH4zdDCMoCmF1mWyyMhlMKAObXeL3mlnv5jonk
WvGcMA0Yfp0mR9QqMUOZp0fOSnYBZNBGGJr/Jy1toaHHhHxhFe7rYVkNPhcXfUHoWNJlzNOz4/XV
oZ4F6CB+tpyrdGv/QOBktnG/p95+6aaxHrSlUhpNXjpSGcGwrRYp31kPO2dZQokF3YAp5XJSmZGw
/I7rv5S/ZxguU1LF0K3ZOw5kDPJgBIqOdIzZH89G1Lhu5AQ/b4TK1C3yDZQfIPPKFiaDPqbUxrqE
o2pHzEaBFoXSP9VN/OYQvWdzYsfUFa7lzvKfzBWx27JJpiJZZVzNYUm8ibkGzO86q5H7LKuIYccO
6yXeSbgLlx3SjnajaVdL8VnrrAOqZtX5W+mF0fBBwVmwkhpb98WBsg/PNBZpjksF09UEneQs6iMf
10wYt0xHj3EppJfqokVkwDmiawhB45uj8eFqOu0rOoQiJ5qBlUHQDddH76CgbxVGLJSl6hRc6edO
4NNh3eK3sPZj46I1wf/DeWukyRR6M9TO5p7oukD/pN2UQhFJmc0yRds+B9IUMkS8VDzr5li/6ItO
w31ulOR4HSfGfkACqlYWOhDD4bHX0flImPiBGoJKnmFoU4aNF/1a9NOJN40vBNoU514FzYimKm2D
yvfVOFgixnB2DMJC/A/Rqfnp5NhdflrX4E5pH5qzW2DoVMiEYc/BQNsakdK/xRX9YP1owO1ldIHI
ems0+4DSz0jnRma+/u2afyKgQOUhJeyGtOZtcDQL4iS98Z25EjWMyMm+ZvJ8MZZAS2xHXjsiwpEx
/FKr5md5HiGLdwvo0/utiiTteW4qnd6keP5rAubDWcj3qrI0vNadSihLSuJ61dgESn29SJEKkLHa
vTxC1z9XdFyAuX3DP9vLrTO86C0v2zFZd2blIKAC0VOSeOACumGMK25Zrcik/LpD9P8xKKQOq77w
rSw8SxQkw2PS/mIs+rAVWsoqDPusm44zm8QgDmgvu5PDyBRxasttZT1/5Bu0FugXRXWZ+5eRiTD/
eKyPtkP0vjcruOfdzZL6/TbVuEVueb776vtPlLeNFP1UIYP6cHhxXofNZYJIPY5fwbRbjCHQxDRO
n+0klkAwEnWfcYsqOppLEWxHKaLLsA+ZCiofwN3f/lRBr6E35h0K2aTMxd+ljZg2Cg68t/OV44ZY
vCtORiXQivxOYbgyJyICQYsc+roeB3TBqwDkh/Kn143Ol10cJtBaV/7RBOX8n0KlkfKlPg8XpOYM
HS3CbPVGCIjW1ALJRWSUXADjDKcTFEEGd2Vz9XYWIOzDaW4P85MHK0iu+H7t6lOT2BsQJ3i5sC7p
45vQRC+3eQcN8n7QFMjE91Ef6wiS+Y2xVzE1A3uSyjUMLA55acv13xmOgrXQi3TiOB7WjuYcxOVC
evD+pBwuK37EHSZcWlmoogxHpEunIa/BbV67+glbRL8rR9hp+tmrb2UFO8bQL9a9LbC+bksl/Kor
TNr3PlBMOPJCnwQcufYRlcAGhqF5OERQcdHMnti+k3Hw+qXX7YV2OGQ2GlJWH+xZMIQY/BZscIHp
VkAI2sla/WKCESMK4cnlHcCovpQLpdrVnM9C9ii+KfYrNJlFM7yuMx4m0T0jLg5Zo0GEHg6tBn2d
AITIfHFoq02OUObQiC7O9qGiq7OU7tQREtlRVC3Akkq+mlB5rZRJ+uYJ6EwPicDdT7dWwH2hAmbc
cnT6cpdkExH93K57uWIIwMo3mwGvyZu4zHw9/5JvjSqN+Wyt1SmhW4C+T8sGetvUH/7D0AXiztE3
ZrBUzUyCfW7DHHah5Ac1FOS5/UW8wCOTLMpdpIyzrDfkrYo8w/n/ME8Opyjdqsx7T7ldTZswX/5j
GPKOaYgTzG864tIdT7sALUPJLuG96OEeUV+vq607S0LSgCcFV7u91stuCGXzodYYeuesmm1B1TD9
Aa6iaYKgnCoUvhBHAueJRXiIZi0E2WGQKH2M2we2y2OqSo/WEK8bqtmu7Lf0RezhgHMPl5lnuydD
RyBRj17etI+Gk6qfgjIKg48C7XnKbxOxo+lDfj2oFMUfypDySiBdM9huWGaLYHvE5yrHnhVjDIzu
VfXopZ3qlj4idulm43xd9qchZcJcU9cGKdeM8mqhXZGFZpP+n/ztu2o2OwXZxK3u+G+eayhAUIP6
KoxFjgDtd9tCzyrCmyj/HdpRwlQN3cMPbYdyCTso8bnr2Ua+TiJ7U7OyXR+cqB/5ut5ViKHplA6b
+DkLG09KooEdO3qycb5vSbH7DP+HeceSHCWiG6WI1R8E+nMGKrER8tyt7Ndn1wcdmLGMqro/+Wbr
tPDC8oWIWv4gmldZyxpbebsg9JtFRggUBdVcJ7rzHVIfu81vABeHxf1xlyrfpIpemNb3U7Pe5f77
ni+vaS4hGeeOvcO7CJOsVZkWLJBtgPZrrdDPkIvuj3wUz8gf5vD1OCribuHthXvjixDLZg+yvMRg
KeI+1FGDefI1NiplPBrFq7tmSJV9GKBTiBDY4mdgD/fdkGi3boOJatyEb9nVVOHrazWvEgV05f9u
cG+O/Ns2f5qocwPuTrfC2Bwa3dyDbqGFVnjkLVjCA55Cmh+K4+Vj5jOqOiWv91QFLEp7GX2WKzoa
BW6elnL8cg9w5NOxW/Ed+8Ir6s+XzdcuDOO9CftF0TbSXSKOmYtIedRR7rY3Q/TiIWZfklo8fXss
lTLXJtPo4+iz8ykx4RmcasAVuRjK1Tdo0ypozD8wgjFsDwfTm3t5lQUJ4wYw94CecKDp8b30donk
JlqLrJ3GuDXtrEAlkm3K/0czhXeXxoUVug/veON12QOpUh7OoLg2VYznTdiiMsyesnE30eeP6R9X
IbtOxVGj3wykGRD+z/2omEUfLrE2g8Zj+jC/8Jx/Kgz589DvWBBB8JPh9wmzL+cAo1HbxeaAo82Y
op52RHh/gsgHTNmpMMDsZIjpVPwj9lzDsPbkjlNLMwz37GvGq1+oipbF8MIRNgGI/9mmC3rJlEf6
1cOROKpTqisxIPBDn0YZ84w3Nth1wZsYaUY8ZYAHAPP3Xyg3Ca38YksW2zFpiq0ip4JWJFdF90xP
qzcGb4U66QiEUINbk0aBOrHEaNnzuKLTEcPbLA83F+cjrtd4Pd5YwHsOqmJO1VbpXcasD50QzOjX
k+VUIn8+bklP0c5yEch8A9iICvuHtLI8dX6teJwwbjVAKhYJWk3UccQ5s4Yf1At73Hz3SWAkmNpD
zQdbHflgertoi7Ra3evb+zpE/8A/nStwKOCNKtwvgKz0c2tBtZvA4PJUqyDSH2gRKZxSiioUAO36
LOk+IrBoq8iyAEVSNaaNBEr60+zKxGQdSC7aL0tgKxYnwwVjjEnYae4p9z5GzkVZG2s+zWpYGYBZ
XUTeDIxYnKcMQ9KMVMlS4v707ZYTxUGOUjOD2UGFhGp5s4LRqnJQs9dMqu8hAtamnN+TJIvul86U
MppFdafMFRDPrnXbARfi7ak+LjLWIHuKgfPQiFOnHqfMj/8Q/M6QFSOKGG/5vVBTDL4/+cpaCLZU
oT7yBn7uiQceAwOkGg8+TZNBB7/RzNEPFYJ/hx0bigg+tpb9TykIL7Hq66vbVEkahtjfd9EHB6Dp
zx9c/7q4yvXR7QQHePWTCW1riaTBFbq9bsm66hkDUKCzCiouGgNXxqpd1xqG606CdqA5E5sb8+zN
AjPh6qO+3+sqf6XFSujnnHt8Am1FK1cvCpICGcu5P+sUsOMwW8+jAxY4+awoIWodTFIDHeGWEAR5
Z5/ZpfS6Bv3TsvjW/Rp/WFi8C4HV4d+TRfxjQg/FiWIBl9q18/0bC7iS/dDcgqMmYnSoNPmFnOIV
AK0U5vfKMqPpUSm/jh9S32LmyjsyOcn4nJj7FH0mLV4LKmCVSBjeh3QujrFsHtjTyadlIgyvUvj2
WhZImYDWEegMkYmAIXyUuFIMabu7Wj98WRq2a7Mgn7TpkbFrufkf4/hc4V82wq1z3QUUOYiMFLTQ
Pj9F0wolX9gfI6H9Zv9+b4y3wPo74LeNgdZhZrh+dy2lkZM3h+65QoJ7L9SF3D+zNGeBZ6hTQdG6
HgYL3kfSK2Nm5qhgQOwPTSzrXLoQc1Kpp2bROOxT09isb4Pv9JwNlZ/CBKXZg6TO517veGuA6Hjm
XcRz5ml7x5Yeqle3hYF5c28nx30iXOZUXU06EffPukQ0blLXH2DrDb7JnuyF5x6FuJauVzOh5FMX
PMMtB57wtpokRH4u9tz89enKZV+GaNYD1gFebrBF5ktTKpllP0NA/vtBf0wAvL89r1KnZg7aKq1y
amNdCS0BL0/ztX/sHuOxEGkA9ZGVp2lo0HMe5P0SVFyfFq0Mxy47nvQ/pKhcrKOfQlH+B3+b68q4
rtNnwVuzK3s1J4mDrXeI8+U95a+t2QvUKjBSRaW8lMfXHXkNghahe2sfQZLXdLpQ0Ze2L+e4ENOv
ekq5TqROzFlIW+CfbOMNyLpIHCPggdu1nKTwBDU3ACp15EiV3o0goqFGLgwQLmRp3+7LXVwZ5Efl
QQGEoY4slbDemR4wmt41ynXTdhj8zrzkwiXRSZqAXgzodzBKqHqHYg4i00cPJDIfvZXc7SqSsrpz
It986JAE4TtMuXDvu0lSi0n9HHsBufGsOYCbzOv7Q5RvZDEJXrZe16yqvLJtiAKzZibtkzPn1YUY
gC5CDNUVlQkKvmIbiwdXArn/U7Bmor9TpZCj5r1g55xv8YDHltAJCsakSyBrTzHuhjeOF5ENXcxW
F3hvVQkcj4lNtowXdROXeEMZSoYixM9GRoBU6wA+OQoURDo0T8KdkWWr6TXqSFm9i+acnV42pPKb
XiaoshHa6+vNt/V7iqVLUfhAZZ64HHRvmXBqOHn9nDKBL8HylBpbplHbKYI5paZdOPZsiisqz4GD
m2MxUBQtGcOky8QwstmuTZ0WD1Ewb8vTIdZjMPMK4RYxmH3cZUrW9HhLlRd0LYonU1Of4T9gfSTF
e4GlRAAaBunyHjaSWUv81xO8uJpMMsB7cTVzN3fRbrDmEfbBayyFvDOSKW01cedXiA3pdFe2ZkUM
bb1FVhw9WzBovllInryY2khV/ts57fQoIOGNqof9FANwn/mZ8UBmiyWvSawJ/PemRqvGQYC2B76Z
QI/DA31vBWRiXNK7MfKwTD8wxEI/wzyFlmZnsElXR7jvJ13qPCGBezKOXGd/UCbIZTRuyIKfamHm
Hsd0GrEo3ZPvam9Nqj2TjzD4jlp/FbixqZHccqiXqgxmleBQGoYbH5S36A2z43OoPGKHA3YHkYlG
PagNQGxskTnyj53xuB2Btw1dSJlyiM/07VtI6TvMaa1iknToM7/CH5VYO3A3/9/iXaqqAgln++el
oL/AvzstgdOQYLq9OXUK90I39ygpmj5nvhJLiruO9aIQ9FfDz7EB5mg5I3UK0kVu6G5NhPZifagA
voOrR1tRo7qMHl/2xlPibwHGiAhadH8TBZi1J8rwQGM+qcny8AL9chFogtwYRFkKT6BidP2RBpgt
M1Mlm2TDdkq9N04EvlICRNbSUVHvHNMGA7B9j82pHDB2lwjLwbrWn38lDHu1SkJoRZ9XQpCFoR5K
WvWaWlvkSPmvVqnDOVTUr09H0MDzB+VUlXH64gDWYNXPWoK6P3OKKU46uTsUweuyC0rWTYNT6gFY
mjyKC5KRLj4PCID0NgrsKqQCm+R8CknnmeYbJydtXPODlRX24UqkZctTrgyl251uRlRMd/vUXNAn
yIWTur3iqn2TAXhHYAvoVheE4McBTaYrLm2y8bPjQ95Y3D7kUS+4xh/NrLTyQPvB4ulccJmZutUx
Vo6wjcAh1amscNIbhwkhIySqY3nS1E6u4ZWSN1oKlripnFvdrQp3rwheqMcH4VrNFd2SPrWIFaqM
O1sAuBaYWxgWhThliIVXVTlYb8ars2I1c74lhqm6M5b9PuS9DssVp61l+pu80b1HxENo4JYWazeQ
4FxjgACWGOE85eJwEmoIIP7eqGJUIWa4UJIf0udjf5FlrRu/qOZcuwxbiiHVRbBfOW69oWnooIxm
llfjxNXOW2EiIk4zWnCbQ4X7nMBx63BSqtEj8zSMBjlCqpIIjnhaEeUBaO31ElcLeHn5NH09pSpt
SwJBQqzd5TsWoQmwVbYQxDsXzRYWdFe2ZcPO5sIHqSW9Fkjt6DLSeUY6dRUV//G3+sSRQ8qqMLg2
Td7MV4aLnuX0i1frNjnasPRq6HDdzxDNhRRjFY3GBmyY0BDa+iSZGQIFml2dadJAq0Fw+wwtfX4q
Esz5z4htl8fg+/AJDSFEGWiq0/8bJMfPoTIX/oI6POv6JRsQssogrlZv26XIBMIcVnI5GhfulyfB
2fqYauEpRqOsMEjgicHdWM3+/F6gZWsYvNOHASTG6AlvvyOlBT0PuAKBLRu79gvk9gWqCAkOpC3F
jRRQIpmn+KqiO56mGLDq688fGp/4Lmce+xHccuo9WHk/RzcMY8W77wrjzvqY/V+xyK8OSDDv3aqh
Zr3mAh+YbNUjiLcpTR5T0HtFRSjsJKl0orkrAeNqPuylwXgP9L5OwVOg2q6nbDHj6UREZDk76IpV
Fg9+UifraHwlRjPoKkNyf9I76W0I13V9JO4ZvbTkRUD6ncOuZb/ePz6f2TBLms1P6ac6HaGb9W11
KL+9Hxzb7EZ3+dzeOlgMo+gdt9YqVyN3CuG/8OhyqwNJRKFI3Senq1CVAg0c9Y1auiTOMsjG912Y
gIt5NZtO5FguuW7jK1JBnD92owkKPhnUM9l0JsvONsgrz38S1YCoWjWWU4xUVbalbCgMt/F6tfEn
wyzSRrYrAjGkr8Z3zZ6jz7uYOkcZlnbsaZrAM0h6RD+GtBDa61Lc7nYFFpVkQh0lRyQKvh7kwH7B
BaWJ4fu93y0n0UQ31rd23Appxg0J/koChh1+FRhuZa/QS+s9isZmyTKJwBRokG9x9671XbPwfrYm
MBWQvNYewBNUxeTOxfwamD5JXkXsOlTXzYC090GJ5grLrxVuCVRpaYHn7ZIVhZbpIWy46belNXJg
VZ6+65hjYd7feV6d7L5LSwfd9Oq9gRvbKUOO5tGDp7TrUI+Y7PBSSJfSg553xUOhuz4Sl9LsVAso
eMcm+Ul47DP+t2id68mF9+wfaz8z6uvuG6UO7hn5lIaXFE/0jMOScE+Z2rjjXjAJlnCobo0zFI3v
T5sZN3qg/n3kfST81Kkbn+Mifh+/twgrUVxKJvS/rLxFO+tJKF3a6ClzxUbDLFX6EQwokxvmWUe3
a8xUFN+W8ibyFB5UazNVe9d0fY8AuFhfNz0/sWudzDmAqs8FPB/JBS1uxu5a+zzb4jS/MzB1N7hq
BoU21bdbef4fUsaZs4zV10ORDYQTA1Y0GzLwiWEuIh3cMqPlThpjLcbdPV+r8AoR4SYxjKfG3xho
+6A+Ws/tOnVICdn7TE25HhcfvhDLPRq9gzgYzScaVN5yVM9kV/FKI/S/781yPl9iOOZYBW9G/jEK
kqI2DDiM8szT+V9HApIzo1PX68+Qm7yArTYJ4uS10VRvxZ/QTud/XaivGf3cRJMu/F6x97VW+vi1
NBqXAyuT1+aR1ylTV9uupeO7wrOg1jdNsOqQDhcLilzP81qAQTeBSFWYF3gOnm3OOJSBn8AU38Lo
UfbS4sQWVBZEE2Ja3yQWes09hx+eaQBwI1Lq9Vl5OtzLuYAfQcB7R+e2WG/EIAEf9Ac6WIpR87zk
zxlfA2ZP6YSyTE24SHutwyzI1I9XmZJ3W80HtmqCYCKJiGkRRjB2LuLG/cHz960ILJyaqlbG2Irj
25Vdf/mRZyzv0IeYmBrKJzF2olkVFi1RCON1W1Sys/6AfMUtim8060QsaIVuZsugITnX7QscHP5L
wDH5Re61e813Y9KJHFSkZatmBVlia6i7U5gO9OkAA3+mdYGhQxyOE1LjmcWXNx8WnmFSWnKrhHiy
fUvvfuDcULyxobhMR1g9Kz1NXLxesG/1ougVISo/3NgcZ1/lB2u1zDa32ulKigdBUOwq68+FGfTE
3WRWeJmxGFrMvcswS6n/MVRcGMCy/8rkoGrNVXtQQhZ0FrQxlkcQSobxwDgiePVAp9ZFxfbYE0pe
tcXBCti4o/vGupYAzony0+gnt9xfq++LhxgQyuJr/hSE6o4gxdgsGX1mpbVLizpWy2UTb1m9bAe5
8Sn01iZAGng+Ohxr4NgtkRcKvPt720M+kEaKymLDfDXVQtJr1V5lpZ4j5Wtk5fkN17qd1swjOk0g
k+scwWG7WIWnQEb9xu7nRrcQTe9GLkc2rB9g8JTITjX5EBnsQHYHij8nikSs3DkqEzh2j7ZgyvTs
OMg0mvayWuV/2Lqy0bil6YkkBgIXhfpisjLGVmX9SGm1Rdbsm9m8jZ0Z4txa8g89tgUaCduaImnJ
sokORTwY+sHXACfr4MY8go3UVUmKyQVd/EO+DqfHadki8VGaOQhSRNQ/VBxg54wgsyLCZHZ3ktUD
JAxJYXPsFDbXwq21OOS8XN3KbwqNYOlIRLPV9KmROEgYdZFLx1AwShDjzhVnTcjx18zYaXvzQ6WS
pzLIBChBzR324sKLJqRR1ZJx2NKVoW24yMp6kIcpw6UZtFIkC/IrITREIoITP4kVrm2DNXMECXJK
D7OBsEEcTMg5/Ejks2jpyLM6H1dPelcYOFljCBKw7qEUPL3vVGR4Tn4DYQFezcfsm8IN7mSahMXx
P4pQ8sml2/BWPNiU1OuPl+0SXlzZiyAeVMMHcr+JahRDmUbmnfUGe909p+q4+xekS8ktZlLGhpA9
Hk0APyLBwV7bZX/Sxvlled+KatXS5XuqfrKIWUbfVFur37R3Znhm7kSvyqrnfRNaS/4I+X88fcb6
8xeWM/DvbcnO8eiEvFLhjfzvxCNxqvd4VoxalBm2BF1d62h3xki5Ih2MOaCT9MEEtwdrX08VV7te
eGV+G2hYlraA4aOk5fXmFltNI/+fZAyssRXiExEsxXU2yddV7Xcz27BBrj3f7kkIVpUdfeRFtdMJ
2mLzaYLEVYuMZ9pp9uBGkHDv0p8USnk0JAQWvmRMu8dI3AlrIT4jwIBjGDbIsz1SWglvUbKp7rwP
QB8COnqs7vUQTILXdFidJq0jrC6kiBlAsRiXQwZ5FxAJw4r09IYZu+9miJ6hrvd+weU8bajyfZV3
/esJ9ESg3yDkfG1+iVco0yZFX0PSCGWyZSiWMvuTbUCd30Kg5zdoAwhqe9lnTJ12myO11DvJcNio
QzmxsSlFqioiKPNCBwfu/oEVuJdIFnwXmPLDWZjAm0KJZ5Mv0zJkjLe+vReEYhINipodRL5ls8kU
cvq368+QkKDV2y7LOGCQc37oxFZEZlYOpuNjcxzd5s3xoswlHCUFmHk4WskMD8Iqimc1NVmsaNEx
1X1VJUjlJdlU/mLJP9m2Zg9CUjFcRVYuFM22ObQAowc0+Woe3OpB5+aiM1zIb2VKFpQg8s1y5lrg
8nfxBeMl4I72yE0D4btaLt5BL2fGY3M046i4jjopIiQzNY0CvmlHRxaVfDbc3XOsl0P2OhY2lb1w
nKCDggBur9j4KZPXczsfHRtePbKTvD9VtNQORFEhW1zxlYJZ7wfwFg4+nbVt9T+yqQxlHY5V9vKd
BNNU0xrAmQ4bZzUQEOQ18CxbdoZqvkO2LNNCPk0f71obTyuOwXQtLwNT+7w/8uXdmQECFnA38HWx
Hov5pDjmF6QjL2DekL1KnJ0IlRRDHi8/b1YJAlMQjC9GIG3LI9uM9ayxW4jYK1SIGuVd3F+kcRn0
KyAVGMON156gNp8KgPJPNK0ongZZRLxIOsfDMCmj9lDURuH7GdxHAAAEmJKZKXOqZKJr217ojqXQ
UM1L8dLneXwiDCj1R0bRpWpsc4DDfl63Wj0ZbME+9ILzDwSbOg78ue+XkDTUmeUvu0Rs8KzaW0Ve
mYq7Dr3Q2LMk/4yBIA8KpOK5XFxmdhs7Uj1oPU7WGMqt2ALdf520A9ANHDJlOUW9CX4vZabaZo8M
eWD/9igvV3r7l4BbSsKRutGkmX+3JZ3Ezvlzb16RQn9GOps2vqksp90Y/OZAcCmNuvFytQJ1u2il
kCE8AxrC7ZNjQme1coscAu2wWebEhcyDmSBtiAuvoQjXCC6csd9RVKXIw+MriyrJK80b8XWXo9CG
/StP94CPcm0Rk7ItdQCMUvlSimtEdlYny57yRAHbdhnvWN8yDx8j9PPJh+Vd1W+D2IECXDG88ILt
1gt50j9YO3ofRn74e5ncxyi8bUt7eryY13a5Q8vt3buXhz4O/9FrdlGUhv8dP7+CCGnXLmCf10wr
pA+OYfEB35rnjb5LBkIvD3oL6li09KOlvmVuyDE3HhwWfxHJkwmSJ2/TiYGk2Eskl0xZWWzzlTiZ
IKMkUr8RGLTiygJPQ16UUfi7SKI+3YX/j+5rV38Rijh2GfjXagpLLlbMsGhsT5NkQyz+adm0C2YM
JlwazG5/DzImMoPwIhkJkOD6xz1lyL0iGD5BFjDqSfy1i8+85YyOZoto8vkqZSlLtfHVhSAn5HyR
2E9PYx81TXwzsKRsvQBZ4Az9TH229+A4Qtmpl1UYBpsNjDw8tSq8kJ0hVsFxre0d/3tanydCNrco
QthfVA9RxHO5araNaUlTrBdof8Iw9OAzYv6GLhHHFNktIA1NHb23Qz5DrFXfvg+e9T1DDuf6dF/C
4JZ8qe+dJ2bpnNIQTS7PqaHQ0B0GirYqCjSY16XHg1X8KF/F0TjGuMSI4T/G3fPpis8CaRDYhwI8
LOJEtSFdT8zAPXAK5qoj3HrYs/ppbUlUOEVwFRGeXJGkm4bchTnlBk6+sEX5f0zx9mRBuW7MACan
lJwk1f5j5wsX3cDBp3DhOS3A6s5nMm+UmST2gyi64OGEAiTGobsWYo7va+RRXIaFWzVkUbsP14k6
bIJAX2NPVS9rELJkLPyMdF/w6wE5fnUXpz4QP+ucW50LW9Liijhy5Vibu83ZLQt/4PeWWNE25X+G
n8oPJkNYiN7gF5GC5sWk7WO/OlkiSj2bIppBfZ7xEqmFfD1uNb6XBPBt3Q0mRKbO4RWKq34f/CW3
lQHtKh4lkxPHTgRMU1DoBdWlu/QWo+RpKH8C6rVfFM+j5DoURFLoI5MwSEUKi1uuUeff20CXr21v
uzxmvqSemRpuqKM+5NU1DJHfVr0NkM+sEywQRmK4w8Lkol9+v9ieOMahaoACNc1Pom5xmFT63rvD
zQr6e48hUqB+CWbOpl6ksuhwIJMWzitoY8nActUCqr2QEEn1xzA9CC/TdwKAnYgUneierKO56ht1
vYRlTwmS0w0no51kEnPoTLWEDCa26SJgSxNk9b6jmroffHuOLB+2Ccz/WG01huGRoACj+RYy4EqO
5EgulnkjY376heBu/DsQx9JtDkakct0RVxsn1rsrVrULzeDs11VBEPczai6D1nVrtNJz20W8EGrh
I+hZ92ZukOERI9xvxkHzlaz6NNonGTUM/yGCzSNOxVTI8v05Rbeepi7rQ5eNmpU/nr8abY33Y49f
iGy8ltyY8zJJa4mgdB3cnsAUf63YJLWvBAP+XgeNdErgbjhn5U+1nOPymKQr/rtj74JlOimMDSoi
IzmLJIrTvg24Ajjxiquy6J/p2yI7+OPuYGOfMYjg6RLYs1NuaY7MB82PCXNlIuLCZ7ZBme/5bAWk
m6wFCupN8g1967R9YLZDjvZhJ0ujBni9M+taVnz0H+vTDgtFgPDvWzMKPmcuAeG60eUf4jaRLN/b
rU9/oYMVL3Eto32Wi/bwJW9kPTxm+aFHtzMwiECbKbxf2N9IhE96FMtkb1Z7TXYqVtj9w5+O1mm5
IUC6BX8nt5CzdKTu4hRZaqYR8vPEpy7yEw3rLPQKzvc6G/hiquVmYRVYJmehwbXjsfDRfiQsfoiq
atqVSLZRf8QSZvPNzyrV5/jyvmusy54j142NJ2JhD0xzamUTTOOqTbwLWPcetdp+E/tZF9WUH5O7
AscwTFmcz54+whOFUKAdtq+v8nfNY1BLbIfDhNvT/pJC+TEXUPkdA7a80/Od/cWg1PFJtYyiPApZ
8SAVpNtPhIJTjgPAvuhrwu/KVWwYhRyK88ojvf8ZXbX5gjEbBlfnNenxBNaeJywl7Wsaiq8fCtC5
34pul8KvWbsg9s3SgAtNrmI2A1YwxpAL6MaFaybh92x7YHwsZffycEiRObsYlaP8S6rkG3kYQ49T
LNnXY8PebNwfpRkg4vxx/2MHKx4/7vAURBu958v1DCO9N5N7BkMvzSy/BpeE13DWnDVs/c7/t7mG
ZwnVCqqcIU8kiamWEqgkGwXmIvfdvJa239L21HHyPbB2G1zWq2JTKD7XzIx61S7y722pvFpHXQ1I
8mSIi/mCcQchKQmegZITRj5y1HA9M05+/vYo5lkiiqu8VJdAbfvbms6kLA2S79gTrd+2y9+ns9jr
/vMpXMWdOPEsbb1Bgu3LKiCzpzaIkU0lkRkL48Iu43SER72k9gKq2tA0c7ULwx9jdwE/83Stx44c
3WPgibaaIWhJkRSrgb5FNg5akfS9eZ2cKtJNSHwPcEVD5P6HdAAGw8+aqJyoT1aPZqbpAtixiV7b
kgDKb6OBq/mOUNKM8ov7CPdtf4gByoNGNxAirASuQkjBq0pZ6OTeArxVJhNl9AJF4Uqmd7FMvwXU
9xFdQjZrkYBGZpXjDqyO/oI36o4CTtstYHP9MCfCFZeHZmJemB601+vc9OSpb0vPu6XAHl8IbC7b
++RThm99lZ1jNZKGSWE/ZzE5cYlm71DVgfIIBUe2xJwA+I4DvKqiIvh2xnziTNlPtXUAQELU6DEO
33vcdX5IMXjUS2KUcQlZKmdTv2OarkOrEVm/zBovJAQPICRbdI9SmnVd47PdRj0cJGFh/xJATjYm
MSvwM7BLEs9Zue5PDKXKVPJx1SzbpKJlaPaKDGloM1C7oZ0wc57pu1UnrhXC6EtwKL8ssxTkM1dl
Mr+tzZzsBUR5nbEBniTVB+uZTw1GaiRJwokIp+C6S0qMycA8yPWi1vw2fqWvqtJ5M+Q+iRMCCqM3
OuxWb/OEM2WSM74+1NiFQYnziMwAZnMZP8UmPmYAG6urMi23yJ3v2SaT81V443KMK8Nc6bNQTxzf
LcBm+nUjvIRNEwhT0T6gvEfr7VUXsVM/eT74jlx0XeCf0QN986C0wCql93pIlv7JjtvTl9cnj146
XcApg9sS1LCKsZ0pGjQDxJEi+t2+nMCQcR9fuVtQ/A3AnHNyn/w3DnxMF/QUYz0qymdcz87XtbR1
FxdNlYWgt1DngKR4ZJROEl9JjeAv7HmqHlzRne4HN+gwcZM/dd5Mz1vYBLe6mX0GxxJ8jmQvxUCL
RBD9bEtECjXexnll40nJrgYb3+3Sb9LowKR9kC8IHNow6gO8d48di0sRBMz2x4vRBgj7OSnUBalH
6SiVog2m0t2bjIYzetoVikgv3bwQbl/B7GQOehMcqKisN//wLSYgSErS+Ov3JVCnsrIGoiXjbRIB
LAAV0/5fBfStCnyF+IHIYFPaFu+ljRYdn7Hzy7krBN+wZrL5luNI4PYelkDd3M40IOZ9nEbhArGC
ScCO5XoJ+8wFNpya1RIGNXGJgHraNiTVRK5gsckQoI7JIBIsxe7Om53EOQyLpLrXBLVvAbIvjc/4
He2dTnd+DPnlH922hat4o+EKHvFcXo96YG+DzsCaCpTIVQZ5h7Xtq04mWHfRxSmDzl9a5IGs+U2V
/Hf+aIrT7n9j76ZbnnBx0ryhTiqvhAnnWXKq35SYFQw8MJAuTpiw2Gg/eZCV3dB+2qof+8QhpoZw
CErrpLDtkECgM14uh+vylobwNcXXXGo4aB8ciOx7bH2rguO54qb8mz/lBy1rnVmBmU2xFQ5YRYTZ
Fi/rA/t3jpfUi7pA3pPtrbXj6I62AJ3/KnxHyL/xD3OuChOeVpLhpdPwNX+SXPOxtZXrHFMoRSnH
Rd0qqIQojA5M3uXbN8E9cM4tNtVeJnpU/TtOr8Pf30IJK81tFLyOvA1Ky5n92bagyJ4cz1Dc0LoK
tcvmCf03Ev4UBX6Ha2yjDBmoGnD/AMDNYyNwY4MgakOJFKk7AzAxvd3u3xo8rHPWGiQYqtnhf5Ww
a3D/R/SEKiK2EXBhrV+KCjOGQIlN9UU5bA51VEfPEXibRkwqsV57vYXY0mpVjNk0xJUjUyMdMJYh
V7fQ0G01TXaRdkwLuqjIARQPsOBcE7PtKIkTEQdwg70GXD1k0dQ+xV2R4EfbdlQ6GSv7u1v1/pMf
GE9nMPvmfgjqqjxoC6sBlIDwHzevUeG7y4AScx+Ul08Ow+IjKvXLOuo8wsJGARyvjT0OG6m/bGnH
3tEmOcA/SQoElD9oPntw2dMNvAq1MMNogRkEgD8lt7pUTYFmwHIAiGV4643+7AGEioP5Oo2BmWU0
CVff2LHmjMarFwAfevrqIGMJ5h3NEkGBfgVLmMghCYpEvFur9K0LqecCTm0HtE1tRdKMHWDgVKfl
Us3BEj97r5KjeBB/r1zAr8v1+2pvRfirxLZbN4MI1QLaaVkv80R+OmtRxn00O6vaaSWyg8bVd0HQ
kR4id4uW+QtRVxfbOLbYhMVH3k4Akt8WXUwsg4l18f4pHKTJXQ05wSwYhL5ENScYE1bKZGkwLCjf
hYZIPIW854LScFOlk7veFok/n4zzUZFIhV+rKmLnrlJxZ9P8oGWJDF0uuIdYAoSzOigZujeRUx8f
QcYsQ9eXLXFk8cdABJb2kaqyC1QwklVW30IZb2kVgijm0KiG09HBz6JkCYXKiqdLgH0mZqlnKs+n
PeVrkI/QJxP62rapTKWhv1wSwGlqROlMd5X6s97Ig8yieZthrtgxa62nqt0IA2sU0Kcx/VYufusO
vbAWFvH/PaPupN2yUKtzCCn3hJ5c34R18LlxLBTiFu5eU2lkTL9STromF+A9Ni8JDb9qOhjmC8aQ
nJnrlx7QiDwJ5q2WsGJmEneflVUHaOqgM3bqaUTwo4/KWc1zRYPEE452OelyBlOPLi6Hzmt8FI8d
5YqpRIlesO0Cs1R5scKVS+leKj76HD9SXe9yeKHkadKtUlMqanya3Dzs5jxSd1DjYvC3zkXFtbcK
+Bu8Lnu6nEjwwctcjV9nXTUnVxHTHAIRd9pR7fkN0eWmS5jejnqueblwbINLL4aXp+Jfizpfl2hy
25J/v5QEXS4cVZNe9ijtCkc9G6R3DbyEiI15+m0WuPrYENR1B8+nhOQ51Deq3TDSirMHIbTUqoCL
MUtiYZ3rQUeuGAA4HIiqVtPJyQwecc73EAlzq+ZZaA4a77FfqnEloZNQDfJ0yDQQChR0nTlvsSKF
RUUbLRlLgpaWheB6JXabM/NOW9NU35tK4DDHO6iUctmrIysvTJUmLQZHAt/guqgxlV7ZikrXsibk
y4nWoLUXbxrHjHfkdfcRVsW4lnaftcKRkNJ2JQYwS58xf6+FDzTAoorSe7RJtm+42FI9u8d8UFdq
OMdWFBH1Z34pCKEaYM5IAo5KnCj2bFDY2xsi7lYC8N9cE0oXZyzSCfibmHZR19qBu9MSbkrrlDOf
35B4kSl/rsSFnX+Q2Y36S2bsaZKhTL6ltpwLhONdXHRfLi0wlHSyra1NCD4wXExn/ED7D6sPULQP
ST8ecVoJVjEnHoKgtAL7Y9yZdMgSbzA66Dv6UmLnvihqZE475+6+xxyciBvelOjP6fHcm3dJWIuu
gVi5G5S7JOTGwPDgP8X3HK7e//7MmhSZKuv0R9EyQF8emb5jyA0iFJzPF2oJcFuk33afMCDe/BLH
F7quHcZiWEj5WFLHOxgW2K9vkz/QB3lv1YMT7Kr4F7Z7BGzrFvvFZSw6bkYzeJyNL/i9Ellx6QMW
JVxnP24Pf6OKLXwab4DBcRLe2QwRaEZp0nDherN2h9NL+QcpKW9xKVlAjLjDeXXdsuvtSmekpGSa
BdiYDCjWYyrGH0d6w0NF0983qTwr9U5dYM622EDErJEHUp/Bg658ONAa0tFXfUnlM70NvIeGvEMy
lxg9N4yfDz3me+137afJNyTkIRlNVQvJsg7nZ9CrtFiuNY4YZ/xouNvCdGbcgXP2+cme7NdM9N6y
Hc56jNvSKiAw8InX8mabifEw5bMb8Wgzl/KzC5iqorklypoXo1vzeFP+beK0cwhUBmH2dOcw0kDn
37RI1ZyZ22//PliVqTX26e+k46O4hUc1+/SrQjzRCF+lBMaz/8CZPIYahmOxE5pGqjHVsmWgauyf
AzIxMqMxV6XAvPDiGMceo6jaf1vCVGjaqCr/bVO1WzCXX9lsSfIa06Cwl3q+jJu9qlsXntIUXM3f
ujqFFZESBWY3vmCCRV7cYZkVdB9W8Ta9b0aEdvrr9NFoxXnIvM5lKdt6kzYPSl5bcBToNAmsqc0D
Tx4/Ye+ML08DXobg9I6ERs7h5FtHErIvUzCEvNulGiwSLhzLiQDFqMZX0MHy4CyW+ilyA04fha1a
gM9OiZp01AqBfTCTkJAUqp/njWSo04CS/O3X9tc8Nnpn4yeBBBhzhYRAhXkfSgRJsgJNBweBJ1TC
U59wyXAWP0JX/m+2Yby75yUU6EA6xlYuaNEgSqPMVJGa0Mi5Vyy0k/A6stKSsZC+x6cf+uyzIqSu
2orAypismf2NMSjeckSEzm5XoAy5ZfDgo3KTl9MX3DvUT69AVcrCImTjzKBUocUMpXzcLmeLi0ym
FI7wQGEfKEtnxugReZqCdLEMHwY07f8MTeEqCHQDIAWTF4t8NnH0Nk20B9v3jsfyj9yCulV41QpG
UI79j8wagQNIS09LBYuCbioC4cBp98ZWIMqy0GD3UOo7Bc/wiTeQLF+Wt2KjxZz0Wwn9vTZVt0rG
DW0+SpMjPaq2vlMsXpRbhLgCzH16wmcptMFT4/mn23RGa0t1kr27n6nPuJyvZcG7Oa/yW8NBSTnd
Z4Y/0IG/Zxsg/SvOtZNaJk6Jx56Qc6IbhKPfr8CdLYJOgO9uslQQgMM/CnQvezcGMfyw7zyFKo/U
EnMUpn3qFaUtmUQbWv12eldrujP4hHwQMCwb9Q6g46yiANDsmzFQDAx3/GPXr6usINI3zPN7maND
1gou6hpD+zc1Qig096OROnL4JPfkzOaeQXotwczM0hIQcPqdcasw8nuFWZ6PSnraDpApnt7GxPzy
GEF8oLiG9OYWMaCimJ+J6CPMnYHtgPW/S+o/9YEYgmLRA8bA2uUZOfHKcohDJvPjK2I6uWOseQoi
Jzjv4X322lN14w2leRVHYmHdMPx/YZt1jlKLkp6/nd6DeCxBbCou0fQPb18YQffJqn1NBscZIiFO
TgJdWageO/clG+FgoYy1SHj0rVFEo4TdM9/bn3T/aD3MCCJ9aUpOOK/t+v3OZYcjH5Qjbc/yaqUF
mC3BOIawEUQrpTaLI2qlhtusbzeOaqC/UoOdLJjAkFC0LE5zVjzQhK7uCUdvNN8uVLfKkVaN3MR6
l5qLbqgEMV/E6bx6A+spJDGsdloysV5Ac9YxomRdrYvP2+6wXBnuqeGoBiJ1HUeBTjeTnDIjHB7i
zjxRA8nKGgTFBZN62tEUEqdbbv99jzYCp8s+AlBxGDrmuqNNgTr9Gz7f8wVYCCwEUilTDqE6JqHI
ASNAUwqq5/arbKFd2QlxUrD9LaTBpL0gUTWQhG2sj2xjNnX5T3ZSz4e9ST3JO62f/kfUxpzNyg0g
6Nw0SLd4mZUnVVYjmJqJIvUSct8xg9DHuUoUXxhVLjpXDAxhaR0dheXsEPzQW7CrTk+liAlW7Z33
g+LG1/xI2oYFwXv5Jdk7p7amJ1cMWjE/+vutwkx+mUS/LY7zE0hIJsSfVhsqR6jyF1XW4dplA5PG
XehK3W+3tAlCp6WoA6nyBqcEY3hz9G+mBlgCMtfraeRHnVT71vvFsxLmnNUSPd31E35QQFE2V4Kk
rZ1jLR5Wp4jqG+ZWIwqwb7nW1saaoDTYnPCMTGR6zB4Zb4koPnZozbCrg28lgIK7E1qtuz8mBjT4
3vNi6LWRHdr4/cTDzASHFuzVFmcTTPaHshzAacZHWkEHLrwCShj2Pwf58uT/Xobg0DSq9OFbwS95
ZWTA2yoix6/xCpA36V9P2rmg7G5dx1DsNuPKk6OG2BY0WbookE7UxfG1mLquzPwdrjuE++dZ+tAK
8SjZjE8AwZZAu2F7w1wkmIzB9p5km9h0exmuCsalnchAGxRyqJQczLd7vgeoMzVc1VmBupbM6e+s
hOIXu56ivMwWiJmkG+8Y/zInH1yVgNctAh1x4ZYw71VJXl7B9CB2kObVbGs5WVdnINnmyM9N182v
qWABRlwOwGQVLE3NCY7eKcRGU/xUoMoSCZt3N9VYwi0PLvv6NX6Oco4CX70GKCMqGMAdDtXP1iLY
9sixFhyd7qRxRvuB0aDdtNgheq1UED+k76G51IHAXYSpAthvNRMt4KxsOgWaGIlKmtvfRdHelCo/
I7zv8XG+94t/B9jE6eXjhCTuFQkx2dJVPV3fxUdWuIPCzHC2ejzlxqaaX+RvLf233TT/jX6Jyy9J
wMOSZchqguBFGz4p+WnqWoGN9qn/c7cxdK/U8f6uq0DUK/Yubcg7bSN9yuLXQvoW0Z6+L3w5wBWO
uHniop4FGSIrzy/eUc1CTjICUF2dvso0a68SDkKTRmoFkFcSYPwr16sBWRZnPf02iJNh/djxOtyC
4/6Tjh97Itc86X8xGOIiwrrhbZUYoFZwvTnLAslZp7z7iQaLD+KJAHge3iPSIiO0ZRGYvJ06i3El
jTDHwoT0RQOWekOo3FQaXaZ49S4HY6Mz/Ix4h5qqmzEnz3WAs6f7y88oj9s6iDKpXhqsSyKQ4BYN
fC1/ZhjAjAPOkjD3bDJG7hrfddOupp1VNUA5ggWwxF7Dpt4sh/iMNLZOTH/7/DFNNC3wTTujVZK6
SVHJrBD2dsTO55ncSkksDeHCjbWq65zP7xMfPYQXX30rN7AjbU2xLwiGsm1z2fzbcW5dWkYHFb2o
oWYKVUsp/ENm2Cze54xQWr99ozf31ej5Sv+UKpnrgBt7rWCHyFdWUMekHs5vIzBKSdTZGTaI/K/A
UI3L58VYCIWKGR6agw9zNvgwDPOsZWwtLb4cfPPNgEJC6CViD+YMQudNiqzNekZ/Q4UYl3TpA1Q9
jZvaz/RdOiyjivcsi/PDfSo/5yZPP8vSp8muzmrxl/twLxqqAOMCWRkCHF97D7kyPDEB4oK3mMEm
mphyV9RHOKAsXdkkv9upMoPSeJKSUXIwEvhsfFiOLVvpuRS730CaMb9n9hWdzU/1+1R58z3hXJ+i
giVKcCTmUz1DwW3AD//XPD9T4WWHiLDbXPFqLC91LzSmj0Yr65+uazUhDPv+JTlthiYN4DuCeeRR
dfWz+qdViN4S6jQGkHmaRWewANFKwQ1I/uppdG2x8K8OXDAFV18rF5GRZrHGhVSQgVM5XbjoxyeY
GUwU8D2YAnVeTxhfq9su3hUIoF+v4ahJkGGk4CNaZNcrMO0YoB7lNfSNFjaSdJdUbaQ+enPwYoM/
Ad7WYz5B6olP3c0UeW37t05pkylz0pXbZmWVE/7k7dnm1IqpCYlCBKybVbowEgT7nb+H5psLzlKk
/2fb86pnbx6Mbr1hDRNyT/k6CiErE91DtiNUfxpTiKcLOdxhx/0m1gLOp/31j7hbU7ndQ82KGaaD
wyJ9IVla5mAlvajGFawXfHqsdn+WD81DnQ4CT0UMcesyVRoLOXbG7KcMC+SiHZc11OwokCaQe25L
P7QNgQJtLGRqN7CqiWTJl8KwVRSI0XkDQNbN4C9r3rY+JiTVU1ZyN0J90NuDBScLO4nf3GkQO4lV
VZulJQ917L4hKuNnWKkDt09Y4w98zbF8XZ1FyN6q0Com909z7g8SEJyZPZoH/o7vUd3z1b/I4tS4
XeEiBHg+FXvS1IJAPWYL9hNTkQBcrMKlsx0bNz/9x5HAYCHgNzLSL65Z9pY9DazqpSJsnf821g6d
9F3h6Re+25rlzHRWcpaWxGPnsYXZvoiaBO1gTpQibjbdlHh6QYytB9k8GHKoBSJsWmUyyTC/DKVi
5bqDEq2X+sJQZyVdPlROag9b2dFgPmfDU10GZdgXhA5SFQyJ1+9qNDzKlG/hoZdlWxtDg+r8OgXJ
/ZTEnlowELahAbY8JF5ZI6gQil3e37E2l6U2smg5m6BcWwoc8q+dhXRXkrFkk+t9U+mLjxUST84T
mc6aDL1QwHfwZMR5z64Ox0zTCYQQmCd/F5xlrPoCrU8PqYM21IZTSP6ZcZ14tNiLRDwRMEplwJoi
sCf8Uk/T0wBisgBF08BSyxD+m4vmYQU/KVK0ybOsrrMeMosxcY/dp3QEjtvDl94AuxaVw3NvLHV7
NQzYJ6RY5bHonvnFyeUdmbKB6ugqtHsTSe5E2/r59KExeqvNQiyIHPoDGJug680xrR3rLZ0HbFcD
smXmdIxS4tGpbtlt1fEZ4zNXCxbZNE4lupFF/e40pZYVc25E1WqRr2hYxPC4cHG+9L+qkFdwML3r
9eUxyYaoS7A8FIA/xkflj4Q7k7hMAnzIRA4CiEVGLzkelqI503UE6d+KBef3AvnIjUSo0/qXhjZ+
sPtvviy0yXu12Z5bOTksP9fgkCKzIHQrg1I4a3G138BJxycZlJ8lPQTb+ECzHY6jk+0RhFij3gFv
p+TRYiJQgJcLiZZDRDVAbuCBmj+NMQucZ8jA62G7UIflUuKOFVOz0WwddtK7cFf7KNQpadb3muey
I+6mLIEjy+egOFvfijLjSRDFUh75lL7UfC74aI0pVgNTI+rxulYAK7gCdhvkQjnoc7IscvZKy1Fp
92EVRQjXh6rTQjCuNvc3Rb2QQ8h4KPKaPWKIABXJrIHH59quOSDo4YylTZWsj9QRiJgxyZxgcAi3
IdxbgFSIInQERFkMYw6/yGcw2gMTwy25U+Ib1QHYYC+x59auUf5fqdp+H0Qr3Og1jJDCU5sQMycJ
F9WixG9QymFQg72N/YSICHEsveA3E05RZn705C4FNxhcjTet8ZupfvCq9fBi9rfcSGuPiiZc/PEL
XtkD2Ckg1kCSCjz783jX1votUdPQcNaZh7DwenZtR/Ocf+de6tavQbf14yYf/YE1UqdQ7+LNCQZ7
bWR0iObNXgghUNH5JREIJ8LKPFSjpmBJLPiMVrWrWpqhmkr8yPo/cKbn+JO7f1ED9XtDJ5T8yjue
/uJc++R043e1VnzRs7DgeJecXXeRa9nf1HyBsXLMq42Y8M2xtdo592b26iU5LmyOd8U1PltAXwzb
19howxQ6vu0VGpvmBfhxZFIBSRXz9ViVF4diHGt1h6UWeOD3eGzI68sgwgKpDYkWi8W9/AS+BctG
It1CAIx+Xx5sRTqwsI+zFgWb4eyLRqhljinrqSE0DqaXSOhuo3Hc/ts1a4OwNi7srYUp/lmNAvRy
7AHdWMBetU8rTqF+x26S/82eMgNcPu0kJKT1JsKTZjxrY5Uj4DiJXsdllnPRITJVjzkVQwkKYL32
92PBXwmQejLFeDAkSizXks/Zpki/le7UoxGiNI8SE7xCKpxzowWEt0grKuVGs50k6at02Sjgkvre
LgGctbPQTxsK/qRKlCrD3SMpRj1t0H6b5+vhhVoqjD5a9ixUemWx6obZA/NqWcDQj1nEz2FP58cT
ehckullYeuzeiyVaNWWCsQmBXLvtTgUuD9ncBUa4q/PiBgbqaDuUfJQ3Ep2QBntC6vPjO7RBZJSi
jrz8r8pn6jvE4UlcBaLnGvWJf+MnKbKhu5XTOjA13UzFbFVTeB7eh4u7Y1558GFL++Ps+pVjPjYo
Zqi3dhA7xoyh5Vvns1J3kkRcWjFuVC2VsO6xzOO/lRnv3FzbnBhKrZyl251yj21VG9RsIVhzSeeJ
Eja4F2ca1At3Q140jm+EcGoXryBM3Ei/8hrLFx89L5/LzfHQZkKANGXftcBSBg+MTCV73eojWymZ
scSA8G+yVpVgoSY82C8S0WnQo0vyIAvJKZlMAtfOaoCwAXiTEYjNTv2rUktlsiaxNg5F7EqQkMXn
Gxpufn3T3CWU1xjbQ26QyXUbIWojwwN4FcocsoytI+s4i0ATMKuT9rsEJGRJvdHp89qRYgl76qMI
WO/i+vtJJU+3V1LsS+55T0ha7rnjiginj5WcNNKsDy1OM78pxhEiJ5pEObHldD9epBtruCCrk4DB
dW34EKrmoz4So/pbgH73xinIJbcJUDpemXKHr4odXvd+AlEyK7F1hJVhd+BJsq8dzWEyuw7sEEQ/
F5B5+x4osUeIQcXESmi4ctFVqQsr7PQrWouYGqKR6EqtDoYS6coNvg4pj9SDL1KZ0wknlCzrt8d+
s0Wq2IQt421E0lOKywkUfiihCdKAhRCeAkgric6rqsBYi4N2W9zBuDht1OwZOFWxnrmBYZNfjxwh
gongl72izodj/K+y79mhW1CQFe+lWnB/JnpbskyfCTeh4hEZ3nNxTK9Pe5qjGXd7LGGmfm2rOBc+
kBr/aWuSS3HRAunUd7Quml/jdqJr1Ln3iIPO2WjcfbgSF0FfAPki8skGxLbCqXrUulAXqPEsnGMJ
Tm4GOCyZ+vB96hTMOMvvWy/bXyLoyPiEHxAa6JMchBWZwJw7U6PKzrzmOzcs3DLeUsLUeIW3P42+
oBJyekwjEOTmFCLbVmPoQVxaiRkjFLTLYFLWkpcAAcnYrujighz1boDX0nZqFRygFrCKpBEpT2S0
P1j4gerpZCctNDsMWTrRR+ziTgBKH5E21wlky/3v6Dikogx+HnkjS88MdKupLOJJb7I3XXwIpZrp
LuztRF4wLvZoFm4dj+14tBlmvUj2Z8pVzQaR3diZtll31K70xLgBj1W5eK/aWIqyVeaYPd6YreqU
FWsmBwUmwMZbNuEWjetEaDPGwpmhjMrIfT7NY7AcoL52ub3VIB+GdzfKWDunNzUyKaLpE4c2kK8O
xTMo+hrJmhJVdlLAP8G3w9D7XcWYilAH7J/FkSOkDvtpSmU1yBxP9qCu5KHvl+YU1ff6tCIs44Fo
ZSB0YQf/6DCsqyrhyjtsorNgEPvI8MSd/TL1OBdQ4VqJ/QKOUXLxEEtGIs5Kow5OoAjh0pCi2ow+
JWVOiHs3jCFhMwMTen/ylyjCIfVF3PDtNAlJ3SxjPyA5wgQ2G6XfBuTnaI72dvDVsyF1m4p5gHSm
eJ1ZsgX04eHNeBDdyvLX6bXpez+GhP9VPHMfZXfTyLgVx3xsFDBhI1Scnq1DE5hT4DU+v8uGImtW
1n2mY2dGvx5t+e2aJBeUkxtEAUfHmGjARb8kBQGYsidG2gJP/g0JLfqMbNJUELgTdPFKV+YfFTgK
Mnczxkze9A+u4KCTx1QoILNm/63GZTKSYhUSkakrVGI3L/OabpDmfDai6eVrBrWKER3E443GgkpR
IcyCrJAOU4doLSjMvLOEmhTbs2JJn/Trrf9Ob2Xz5EdajcJfcjsGtdUqfhqQBiyNmKPn5Acul2s8
spRQdPPZ8v0LU4vvRNmG3BAOZckVP5H6DToCDOoX7AzobSbrtLWGi9aI7L4ikXKWiwPGAAZ1tDzI
t5xLHqlxhJRdti1WoaTBNLWalVXgbWwm0BcXTRKx76+UH7jgmucQCCrEf398vHCzTe3zqECOszSR
/63WBTPoUiBHDzT5pEb0zLNYhlJwNtVuyz2WJ7YmqeINCIh/pJuBQmsJjUkJUHgjgwff4HqUcbQd
S956CtfkHiFiSom+XAH4YEJouBN47baH6PZ2KNgiBLbmD5VHD31b0suSgwX1+CbZUH0rFxe1pBDb
sjN7AA44KadRNNklasQ+FWLtKbi3R1mF63z5LEK/UzvMZ6SWIlbiL3G7Di0KIfe9mj0z3gGcBjm0
avQATrtkDXoRQzUQDqslQW9olIWbVdFTD8xMO9G9AzBUcxng2KeOSAREVWmRwFHM06Zlzc7QadVe
z5m3GawPC8nfXlWfUOtG7BcjXoUfc58YEqnh40Xf/F7tnnJ8FepFDXrjZsENVl0VoWgO8uovkElU
chX+MIHpnUo3senZNv0B2ZSBLKND4NxtoM/zOZmpMoUjWarfKPtJCuA4cB1twf23KHC5fYzF91vo
ucywwmf/W7jqqg+wwr6U6C8fTc0dxJjohcYzbP4jIHCyTS7JlxEAd6GX0a9ChxYVahRbek3WObmn
N6rg8lH4Ec3GwUeS6b89eZjo0TAIubAp4K+73kmGm1hjC9JILt0cbjeIQELMe576UqJ1HZZ+drdW
aTNomaVm3shhem7TnJX3HyHgrROoYWtlnfcCWYHT/w+rziU+YCnPCI15nIDM9MASL0UJkKGDPyho
t3PSs58MileyRDz+dEt1EpHqsRizum0FW/aQkLOa0EkAGxICm4jgzoeSb20nRQpkgRRRXaiY6bOD
ElQ7ZaOR0nGMiT7m34DwKcp/T5JYHmF9hx7W++tnzbab3+O/y9UdA4Tv8j7uE1HSTm9rmapB7b5v
3LR4tMxJlLTQG2gs7qwjY6KXFeArhY/rjfurL8koTxcqSrpQiJ6lnHby7xBWhJExvzs+fZfdc37a
Buf9BbylapxHhqnunS9DHXR2j/2NxCGDnbr7aKnNVUm3GUCBpNiG1muirdEbffYSJDK+etVjaVuq
2CYpb6Gd3q1VSkPe8Z0Uc6z1aCG363WQgHRugVn72GXlnqdIvVTKV5sCOeRYrkpqoOynLw20PNYT
ClCwckuS5B0lIJ4GD46fyjRaM9WLnfvXhlZlchyruRpRBHAu9cOJaVNkGIy+2RdLmJiggsfPb4o8
38uiyKo9pItbpI+Qnx4uTpSg/X+h1gNUwQkCmPRSDFg7tPYt1FrOu58crQ8CTCg2/dIbU9ioa9Un
oPmXpVBiSA1qnhvHWI67Dr8S6Ae6q5YIgGv1RBXEdW55GI7NKni5NC8VdaUK+KEb5zIfgb6nI8/r
NHNDXgS+GYssLIN2fZmW3G/NivYRv1PV6feUjPczYFqck5vmcT+TX5/JYIaW5eFnjUo/FOc6oU2E
kHUjIiii6Zw/VqSOn2LX4EBl89Qe/RWBTvWCoId9DwHnPxIiW+1lkHE7kRj37FxgnsNpsGSGH1JZ
5RH4QZFDd0ZqPiVd84GJkUisNZQpIEwVJqYCsFNScQ3riWJRiDOuI2d6ihfIvtE3NIhKGJgQk5jO
m2O27waxw2ierFeVmLX/2fnsd1scvkRiefypROoFcwkWwkjZSdMDZSfBaslng0pGIoPAdkAn+mu5
+fxpictWGGgViZfheVZsW6HdhuqjvwzGREUd1W20Nl7ApwPfIjLOPdBky0P8R/x2tyUKSaoYwXcK
xvHQGE6Wv65kNwOqvtYIAb5lFn59s7MLEYkTTHQ+LEVRjXJMVAba5tD0xCJ5L2XplE8gWkPUelSk
S5ARXH4C49chy2pNVZY6rCU9y4kgcUrZfiS8VJaYlME5mWMOZlFLB4ztKx5pTcbGQKDbxUnjJXgI
l11Mx7bPILbwyRY9OErTsNvBlyi3dGsK+S7DVhLXMRoqWTF52eJWiag1arycL4iNSYFzRX/N9aWo
qLyEViUhAMwfNlKxEWIZ3UuxrQEUfeB80/Fr0E1AwRd7UEAZKDlvlwTnrP7ToF6SyAE5f8WbVKdi
2EG82/GGJqeJ7uhBvYMEKoa0nG9t6S9KCAYA5CvyhP5J092+nMxEKaqoz5WKPi0FKDs5gS4l5Ob1
mxbmCcNjjl5jQA9L+KP33qKMi/mkacHeSOKWme42ifFdE/H2yGn7vWV5lp5lHIg73d4lANeajV5u
vhHxI8D/gDJ+kmAl9YHPwVcLj8FJJh/Vxhz9Q0q+PARIJ8tJ4H2TfH4PI6aXCGPzR58keFbN2KS0
E5gA9GZ1v+GQVXYxRj2W/VIbKxqptiGQcSoq5HOc9FNonPmQAetqKbPymaanghCBWbTgjAvX2Cnf
NwHJZIJG9eDXMQSiplMPryE2r+D1Un5rx3gNRVO9TLiwYkA51/6l4FI6rS0fAQvsgU70DToybqd+
ydWdb1xtKuNWPHfsFydQluOkEv7dmQvPYQ2C7prEQyDzJFyV416ZMhsDf64HW04Ps5Zsgs1s8Nxb
esSky0NnqRBLcFXqscqf4jMc2E8P+YN6e2KIsVPQvdfPnBvZVK4dP25jg5YofiSmi8KBLnf33jC5
Zss9CrUfKYeJFSWCTPy1CEDJZYYM8wlPV7NKBNl4oH1Jo8NxfPq8Xcmq+4E1r10YGj6dItte8Hiv
Gf/xGMEO7ef4IN+tAHgOB2VjlnJOyGd15gT5IKTaNEDWWgM95gFgzX00+8S9kt+GBjzpzDnR8maE
FQFwmVbgHrTT/Dui4xa4J78/Ahth3wIfZKFskb5uV0Q/5RczHgCHwuUApYlu/6jXz8kGN4F5PS20
ISM/x30f1gLdCp3vsFuV04DpYzzuKxAl0eHSgfewP+1lZy66oQUZ/qAj22IuzVOQ7McvwchIwBgJ
Ov00A937D8scxHboPMQmblsegM5zfv4ZXH2d78IPuMupwZDHhjsZcbAoVz+xl+ydv2jjF37+bpm1
WkTaWsXoJPnhP+KWORy2BEP68QH1ViPzRc4uJj/D523p0hR7c9xFZqsbOEgVnIoA5Kt61GIxuyCE
0nT2VmtQJQItdVZ+NxKRwPsNbRETa3J+z8sPph+kp74zrpiysL85kkoyna5emFeTzRCjwH20xbZj
S0ku11lAk2giUO09KEMeiyH5GwiGqufHJ8zHsdra7IYv/nNH0EOP17lV0PK6wj8SO1ujBLceSoVP
c0nuu3eE4t4qHiuKlEAdidYY2d62g91GzV27vNzqrGCTrYsHtxmvctrFZkMq8eDuJkM8Tnn7vZ66
JBYoxaqcYgLU6N+uuyYjFX6ct3odiuESYiPpgrNn4HXsWnhgmucN1eizghf8ovWzDkTT8dPCU2Yr
w84BT40eaIp4Tjw+kNf8omE3CpmD8YZMnvC3bn8RjgjbBeUg6zCm+FUE9vutLFJhShdoJ6yw2cF1
oJ4sXPY2rgCQe/0+oTb9JKcEf/DAyrXv6SbqJKesNE3uMpaKPegdtqeihIuYkZoK6x75FGZEQGjv
WLy6OHscXYMs0C9vw2xQ4Vr5ZT9xOljw7sd2pDf2o/CWFtjlQzEWJvPCSEgaAoAxK452W6eFAL+F
ViXWXdIIZxWNxq4P4HurN+2gI9yn2lwWZbB1ep1K6fHnpQ9ATdwza3+jlLKiocIn+FeQHyepTenF
a00RzToV3a+XZz2PlswL4XDUXZym+Y4nz5DQG085vAehATOEQ7xNXYl78Q6rIUqy4RkJ9cwstfE5
7sKQ8i01kIuJKA3EmKEQqWcdXMtYNo44mTx7dzMLerES+uiF9y/rDbxPNEp5PU2Ry1MPtCEeQE5N
tq70qHmyPxNq3LUcq5obFRLMhnpxifsgeIn8J4ehRIhzJ3JzPj70kgJeRo8dt30Dzq4h99JfHnEq
zfrj2Nw37p2aFL2Hz8UVSOmhTuRg8cO4ZUot5bF/lGmX9f8ScYH9eZJh3Z1izA0Ytk9TjBBxLSNM
YL2TkGrlcWZnlQnGuFcrXf/CqbSeh++xn7OixyIbE2+FFMOEF8p9/mdQi6skytqh0iKfMp8zIrSi
p80nPFV4RT1eRjnfYZJ3u8aTQdm2dtJgT8QP875c+XhHSZwNBVU9ZRrWo4yBUWaHackQ+TGnYIPG
vEsn/l/xOipVZOUsn/yb77Rac2hI55z4o0BHW8ZQHWoHWeUmhsXh2lX5GabafllC5hBPdlyhizGB
CqsnsMZZUMxwwheU7K5WsMYVXegoccqNeN1aUc/xdc5Aux2qZFmT511HSqJuoNaWOsBa+52ZIesM
VrBIN2ueJNWnDK2FfvZYffK59Q4kUb2OcqV0njBkIVkMc0xpaXAyBN1b1R/ZoImrrluOBPXwV19u
xFRplmzunIywZdUPt7v6xKr2p5jtA82MbdrA82FEgQrUAyRdOtkcJZqB/Q/+y0vWqK+T7f/SLvr2
SWSDuXE/G6PIKNZdRVlnvFSJtXIpwqQ2ZXtEbyOeij+S7IUEpXqx6sodN/ouhrZI8BYXkUyMjCG4
QkNxF7bIfI/jk/C5iOs5uvGXWdvrPrY01+Zd8CPbTXmO0S+KBzTti8MXJ3BHvDLHnHzl8YIk68xT
HtvKSXf1aMuURNzHxR6M4ifHMkUgK+ERtQwLwc8pC2nsgD3O0eAL6R93I+GNVoxlgAhbiofKV9hj
cnOxxujt7m1Od+YnU2S1w9xys6SFCUvFbzBDT/5UQXbsoQMCQhlJXTsX9w9a08MTXbcdzDKmNDXy
9MnQgwHLsTHVI3o3OwuWwqlv14ahqHx7sRaAeBXbTPEvjQM6M7VbnwxPMkGkgVahlw5kdSWz2Tsz
i3xmUgNI19B97xnSOBpTWlzlCZLzFESPRbor1LxDQhd7VSXe69GdfLNcMUn6Yqj1Wuh7ehZsOJcx
fUvcBQAFJp8AmPcyogZq9lik++uBhDoQ3XG/S9ybPfGa8PFglSvOkVr62cfaFkC12pMkDZIITlZG
ljRBgeY438oSjUd/fl2VpvpbYLHOK0BvCKkXfBsdCJw9+JGz3d48eHIo4KewKu55/fUbrsD/YL/D
fZpxU5RpLYoe/T7mdTp3dxmINvZR5eF29DuytoHHzfClJtUXF15V2k4b7IspUlRr1QnOdxQ9Wl2r
y2aPf4wVCUBI8jb1nLFV6hJAIgvS7hAzQMUurF3i6V3c6tuaFIk27mJG8mxnYKxHHHkyrVfeBJ6J
9FhJxrUJceIG5y02FgPKbentMibnuNHpZ0TrEaSqyLkTnM9y90jw03DM8sLXIuEltU5WJc6PT+xC
LBbnR59rPln/xf/WsVLVkEIAqaPlFkImoy5fAmA22K4LIiErmIWDXJ9Ge2mJ0BZbQpXUsxeukpOs
SfdCrMDoJEJ58DtCn+AEt8suY2aNtfpLr3OmAB0IPjDJTjIGv2oQqYLbqZQ0j6Nu73XPQblKJQE5
ZN03QQyDQgcNxLFxpvU8Ie+uLei0nAYyrbE0JUXA2iFiZUCETRchUtBobO7wP5MOOUuEafpm+zxa
vV6iC4B4AjQFHr7GDe8aHBccVzikwgFmffhEkrQj5pG99LMWPuIorvU1WKNs8nvSnTAMa5RrTVyO
41DO9PwlMHXpnFtKNvKhTNtKzquyOak0lqYuRi+lKDRfh+HMw6OULOn9vgl5e6ExXJYRkTmmbyzq
vyunA8GEWcFZuGhSumRJJfeR9S1Shcqeo58KUc0dasn23ea6yhhGrZotkp4tp8omjfiNuaQKwFeU
KMXUvXfkDLm/3hiCrRKFO//csWN8LPKbf+jGXwP73jY/Ivyrbgff/d1JW76G1QrOZBqByfsskuMX
/pB8OgfiM4Rv0zzAU6F4+8nK5LSl4sUdbT/f//OfkeSFH21Io+4nFeyN25gAu2CDd5WIkpW58mPN
Mxnh1lTYp7uCIhmDnla839eCG8pcnBSJLjnHMuBMkKrmDLlQtmWPb0n0hYm5vMxb9BTIzQXfx/O9
jcn0p1ZypPqnmYmKjBoiBN0+Jsu7uYEc+okvKJE2SEQqlVjY48xOvuX71QUWRJ7y9qvdB5q5Pn/Y
4f1f6d/yfRX1sA85WzD2A6I+D0kbWCYzKhVlIz7CZT/x0h3nRPdOWGZxjiwmxsp9AiwUJ/zENGFt
NijWZrGPXPYjBbXvnt89Ai/IlXyp10muatoXN/BjFbSqRYnqXWA2JmOha8gKy4qkLR6rhmDeO8cz
c/M5Gj4QbwIXD9pgp5sK09LwAdb01+xUnj4fZCD699gGQgIFCuTo0YxluSHeeWEj3tGpTmHC4bMp
3Gq3o1LzPnUT506Z60tS9e7FGBNKC57Kpa4cX5/p1/a1V03rtxKgl89XwjB7exrG55BNPK/8Lttx
1PlZsIdsmXkJklUoGnUuwWbBv3k0hV4TWDQcjc9CUUoBi7RgRisSyuu1gxtJNKAUvIJ44is9P+Vn
d1EhhUYFWMVeasIFk6Vsax7h+qpTYxeKFYw4E7YGshGfWuRl6QFnHsQlkRmugSN5zakTVhOOBBMD
CRkGmSC6Xn/NXlAuOr0JV26EmiHALhlQtOrOH8J4WOZbW66u3Oo4ami/AKqDnF9OBrBnxbkPx+nf
5fI1AwHN4ujhky8hv6x/4XTIkv5l6ecQ2e4wEU8SYfzy2T6itNif+/iYMz9NUsxRT7BxnCyR3s22
AbApR/RXujQ4l3ZwFqPiTvjA8kDKIF3Pe/yBmxq3+KMMcIr9UvUj/lrq2hEb7LPmguOvc6AYnK6L
vdX9eQDao8rXdS5feK+oGcw+AX135qH6mjdtDuSKQL/oRJM/2WDzrFeS8dgTDCTIvaXVYe2PRl/+
otowTcdTFRiqQyAfrYdz4fzo0SvGtzajjDi5z6kxzrYrbtoXa3ZLNQpk8BqRuAJOeFBX8dV54wyP
qOxTtU9VGBYCe4l3lby3EuZyzZgNCh44WRPumqDLO8oDtVxdQM4hT/lUI3v0z5lLQlc2xoQRbyvk
imprkR6h5/GmzAbFe2P5M1mNr8ZBYI0k2+JGjRgn0KrrKN31gRAq4Qq4sVrjHb+IzmiJhBkYvT4Q
EoLyVP/roAK32msdc3+iXfCTJMMM69dMTCKbSIBib8Nks9l6AQmiQtIUAXSniqu5UxzHFytccvRj
qzW3Qc4gHcv5UrkdQ+kwtcozmSqqe2z7xARGD/D173cKs0I6JzDPBU6iF3bTQFUw8u95lkswxF2d
Jkc6p0yd0v+8UyjeqPAvUzS8bmAEvZnS9p+OrwdBLnops1GmyzwQeDvWFRVUKA/ZEkHZ+BlzpeZu
KIsZXT00uYRhIpJ4lQYnsOvnpyXrklbX/mi/9fb/cpsi2H+mn9HeIIHPwSkDYnZVFDGqjkmAoGkm
45hTvQbjnqjlhgDpG4tJG7S3ddHSTM4NfdrQqGs6OUXXHUwp4otidBPyvgpSxpu35DXl8KS8aUjl
w2LcjoZTCZS3iR7caCDWBZ/XhcPD5JW58Wq1C5dCgcjotemXndn354py7rAQlYnAsl/BaJLsfP84
T9CN8WC6g/zW+DrNT2jx+5u66SCeraJSYP3qJPY7kyD99xokDUC7U/v0SUXDXl5Y/BxkY4RjTsL6
kUaNyfxd5E3RX74rNzDr2mMGL0uz4itmc5enNMrPDn1VdVzzxds1sxFYPkPdNBV4sE4+TnB5A1l/
MjX89BwlFQ6CvsE2KulzqOGB85FyrQLFcLkFjhN8wMHbfV+rqsuh5mOBMZ3BxvsqHoVW9k7dpIVO
41PLWhhOoSNOfkck2bBQ+cNm8U0f5Slj4HY5WFwwT2rVwn0JzVSu7RP4yYUEZW/EpQUXN2VZwDRc
yA+cWHXYORRpA+rAL4A4TQLFBITx43iVOGx/vubTjT7S/FTpmqoimgj78T/tG5jsg1DO8CLI/C4b
NfKSk0WuF7/dI2aNiTWlMvOvcALivY76Cs7rPzEY8qf0ia1Yso/TBvls0X2e1B++kTHLhs60Tb3k
SP6odcS2eRERTeEmW8gXNfd1CRkskIa3pfDTyeO9LCPjK9qDFD5JmPxZJSYWe0q7zzNc0xveK4Kv
vUkQJnxLEUFrlbMra0ZSSgGanKXmOsWpKlFtWravJLtbgaDcF7Bluqd37HBACuOb7wdHAymC6Vz8
yccZGoi3WQMfIyj4YtWyvKh4PwBDNIRyUQsXdHA7x2AHtcNVoT2l3wakvU3FWfSEBuIg4sJlniMk
zgyi3SZ2racFpc/HBMYzUtsLyNRP1z0/mYLf5Hyh4czZG/J/fsPxW5f7Mm35Ul2XaivFGr6g3e7q
YE95ifynrQvdZ9UOt35qpA+5dAdjr0sO6AJ+otDQQvZ61IYL4xudBqH+zRm/8frWhc23hx4l8+yj
CZ/yTVYHkN554KUV6Kq53C4ColLu2Tgrl4TTbagUiln0HCQc6trkU/Lc3V6q/dQ7EPMtCwaBqJmQ
IO1ZKV7cEhhfYcrysOaqY3iV/Dbp64jhA9gn7KZNVJli53LDMpCT6SC7KC3ei/pRMIDHSdUHpzpq
yBB+etM/hpUE7vfkntoe2QwmSuXVG7y319XTtshUmM5YCqseNBQcOrC+lA8duTCqsY3LJVJl4ZQr
qsaU6dCYKwD2uNmKhkjjkGm7fX4jhWzLi6x0b+ul9xd2gWYX+52fkalmS7kGhCRB5cvcqxn98ZKB
wZhYkC7HfmLeBsAAox5u+B2m50WqQd4QLDI3OZzLl4mt/EHPiLeowFxIuW2LUG4pRWEHxfivpy/R
ZNmCHgMLiVWLRZrwpXcfYG5CfP4PWj/gpj3yYJcsMZ+hdYvfzhURJFOdNX1lRh3pfa7hC0Yol9Nd
osReeuSpuDk96wHjOJBJ/zUylvqUGSn8MIbyiOfqQpaRhUccW9mjDCeO/mS0jlhg7ujSp6dYFlhf
34+skZS4Tx0wpv2iRHVg98cRna+vPS20zMdcCkdYBXn0sCD5C7/TEFgQZCtsEM46bc9QQARQlM7r
KXMzKl8Rg5f+LSBAP+AQZGhiSWXJOIJVDRCJHU+5AuXNkqmQqKYmm5eK3NxmIs+N+HXxTajqnszp
mEZsgfEs+J15DEtHKrCpjAcWSIqg2pqdTeeS41T1lZovEIlOwRe8MdJpG1oESL9NLH+L2KPpn02W
JaMfOsU+BzcEQtTk7E2GUFmnotrrdPFVRICA9D2rSjtrRkN5G+vU71e0cJSunUgKO6L6QOzq9k6x
pmE6yyna32XaeEyfsOcg9u88ZyM7kdyf7Noi9VGiqivh+I3InXCa2BqKdFnuWr37VzurIJfEIpnG
aipRQvXsLdnPR9K+dPSIeBCWjtemJbQslAvuMVa5kwG3yGBFyAlQ6FmUvGQtgNKZe8Yp+o8HsyfI
Ix7pbzJOU9FsTppUV7KHazdGLGSqUS8xxk4x2b3ZwxHsW0KRCnAmIMjPWcnFOkM1mqFCIoOUKBIC
QFSxWTpKvku1Rk1zrsQL4HrEQiDIB/PVYVD0iWEGT+7dAPzovGbFInov8XjezalLQX0rnw3jovAj
bZM4aL3t1jjhCsUOV8eI4+6lMTVtTFH1jRPi1KHgvlIgAOA4XAp0oJPAqn+ZplpL1VQhbn0vbBX3
V+qgt63FR/WPgKDE1Y4eTawp0ecWtBU6LunEudO3brOCykPFznBu5ExgG4bmy6Mo5Sz2USolb4rb
7f/L3CyR/hARL/5jXU7pSajAn538XiSgUM/QUW9p0m537jNbAVHR4BNyJkWwpv9UOi+lAJNNLrph
nlYiHHlnI5UV6S9EoPkxEgXyzbFcHSLdix8qMNKVLice6oiJo9wYzhOjDdYwOWw9EnigeDUeDdC7
BxtXh042E78eqtUNMT+p+E1zXcDP2d8hoMqAV9TmUQbBrfrm65mgprdPxm1xvkOFyOZDxso0gm6a
Pjs9l2HeFZ9veB5xxDyA1XNtymjJUUZeU9oOmfZLEgcFoHuKzT0qtYlZK4ph3+Oq1sHupNX6FkUM
4/RFoJGTyxGilQzGq9jU2/3P96KZ+mOJ5cWyjUld1lmtSDC5frlt9rdSaUcIi3zJVCcqnf98OabV
SY8c5i4m0WI90omIjLlcwkSBYm/3fqC2Ku34Bb8KsjHhzgc3zg40cbm1FqAiQMR+Nbrct7jfghE+
RdDFXSN27rHwh65WCBS2YCnP91RX/oK8JHngl0tU3NEv6Z/RjLEHWfJGlzq8gK4hH/3dZMsQkm6C
pmt7TthyxSG4I9Qj49N5W8xg6ag9llR/IyAvCqwugnKy/GwUdc7tv35h0/wSyaDJuZ2VU8aH3vhv
8fViUy5DWoXTS5GX4ANaa+cbdECMVKQLwMGUDNsvTobLXqqQfqtPjDPVrdZeHxe0TgiBhxKqd2hf
ObBZXvEeq0hh1IWLiBWYGgHZM9i37wsdCXxdDE97//3XcAAqmASKlzFmbC6Q9+P+LnaFCKIGp/rT
gHL99swELRYejk6Y5upOR32bwOKXEVhelvZxUfLzjBs5R/UgoLSMzqURTHHjNKjVQac6xkz5U6Vj
zngAyQUvEvt/gZkvMp21dF6VGdGFHbtTLESo6eOoTFEtJVOTYKN9cXB7Q+t2Qe6Rv/LP3P1oYCrR
Vd1+Aq3V0wyNFzCpr2pifL1kYz0I0Gy02epniuD0lOfN4sOekS621b+YZJgAr9NKaQpbdK6+jsiN
c5CZLLkZmgIxDy/dqqMwBVOInBivQFlMxKMJRBMyDpAxFdbuLmRL8jsst9Wx/vVS7NRcABeA+0nN
t+kfEdyiAIHrB9dm3Wgj4LCDJoR7IdZnBJQPCok+46emTC7gpIRgabH/K49ydRcRvxswAxrwBJ25
D0KM2JEP0BDXij7JktpfsGvsP/ckrUSH512I/zNl6trD6v1jAHcuu1Ev4WVT9wfJOunpnO43Gxnp
zPwdEoK5CSiT66wKnzOAuflukOeN31930SPXjmZ1Mlp6wuRm19kGExSImfgKjt0PjkDnWRHVwJ9e
qQsEw5Nlwa6ed95aIN7yIeZ9mzNO0HO6R5fd8w+PqvgS8u3B9MqxeQ7DlEduKnJ8XbdEq063BMv5
lvgGmhXHgyT80McTJusWyDSN8Ios37HTpkvTSVqjnSFJjBQmDqaW6d9l7UWw3TAC/dFrOKeB3MUg
byzYrrDq5D8Zvip3bzHPgDXkeagysMrcV5hKkpnvRJjSb/dRxFiOlJtqiGtRbxTVxDlkOVIu1py4
Gc3KquWMOxtpsuRUCj0U4W8dVvEULoxKppbX8FkE9Piy5gDpkgv2mkzb1gGi9cnPtwRAE4hYPNYX
x8VBlxv+QiMm4+bsiSTq3FUXV89IIFJvYRdTUeOKfoZFDdji2mDGWTrZp0lXG52lYvG8Csq78LTs
1NoWzLecK4LHt6dr+lNJoRSvTKjaAis4nyfRpAdHvJidHlRJ5L1mhebzlv3QuoAvcieZ15JjiW7j
+hRgzOPbdTq6jgrASztSbJDa+77RNc+atDCWvufSAO7RXIbXw8yO97dCE4EGbqH3ro/KrWGSR4aA
kgdihpbPEoBqE4DuCeowhAOsonJalYvuAsTasKtRYO65Tp/auSAgkKY0aNlOdtX4SHdgWvZMQIYB
P/9bVpgaJURrLARlBp10F6APcqWBM9RQXLUY4lE9DW9JXNRYUrtoUYYSj92DHhNgoo4jfT0e7/Ey
w3hZsg4iUoXxoiPdE8egH9xD3l95Hn29a+Dcn8qp2eJrDwfLVKjBTrM3XXLUg8LqMvHA9S6S0DlM
j8APeFUY+sbnoZ55OJ1GkoD2jcTF6SHNEq2QI65EnA5Jl+dIlsAF4QJwWUA5Pnd2ODb09jrgTH83
HgQVDPGSaFtlh4KZ+0oUR78KjRMN1puQHkWn6d21s0NSyGFT7u56dMSc/p0DtVHDNh/9280pgNYG
X2RW1I6xW8NjL3SgI4C7QH/CUPVOYmRUOi8+aw8gdWlFL0xgU2hIB2KcItOaqYufSEjmgTxetBYQ
YMLYQlk8rN52ll/D5pOve0t6IFLT1v6PM/zEZQezx53ak7oOwBBRt94CdJfRbgyO2sjsKtJkQg7h
HVr3Y4ieab3J3ZzUZA64owbBcsiSrqXXnkH763x1kUZN756ZOhVF79Puq9fz55KHvx6cnC1u6vBw
EXHttz4J6CFipV+ikxe4tGkiRiffpgklUXRFRkNsZ+GnVq/gWiZFrSBsIoExIoTtYVUvXxB11x4F
kOruQxytoRqoTMGlEticEZEKOms4oEwkgLOVDJtt7lJ3bYdzMmmwVg3sKNv8Q+YX2x5hB08fZuRu
Kr0Wgb8BYLhqHtaEMke0PEMhkwTknj8MycHdVGvKtdGIZvkZExcS9d2dDweiHTuHS0h65MftGhSh
3UK/gjVeBL9+ACdXQSC0b/zHegbL4hGq8RSNCc0LMHYOyDnQwhhps0CFk7kkDaOlzG75lT8DvIAw
pp0YfWSHwB+s7OHEUvSsAi2r9Ked9yR7O/DBAoyPKbSlhRTrs705wEObFTbFolJ4T4prfkkM69/F
V92lIlAQHr+Xa7KiXYtn/eTdlDiRQR0c7uax3uKfhp90CWZMVTcmYrpZfi9Ge49NEM31J9GWEwWl
NJm8vYKgsywHW7NtzR1a7LbAaQQnfLSjqBmonJFhCLvrm563ZjHpFhkJt7F8tXs7SmWQuu5di2fz
idJuTme9azITuRi+UZo+dGCAZFIx+3UbJKHpLbAZPidQoPw7Mvrbmhkj8q3hm40m+wtprd6aeIHl
Rm7WNesGWxM0fsVAejsW/B07sAJblkMV0+kDg4yibTJYXdWjil3V5simn9qYDpMFrJhh3bzZYCpY
fcZVDc+2zOAY6HN3njv+2Ey4Zju/BpaBekZfEWVdFbv6UQS52STfkWZK3RY4RA6dY0mT7kfUJvMS
38oAspeUGGZFf0leslO20QKWqgi50FeNtqj4adpQ7tVo1cQ1BNfNGgi0ymIIJjmzBDhRN0Fod/Z9
gpoWZJ3knbsge828rzzRnfhJ0ROxj47dTGD87MKIfT4xCkFF3M17zwTJvgGA4VETZonFMMtd2vw/
RL+A+7Bky7Pc0r1aCYl48HDzoqK+gqTPwaTl+RrRSHhMPiZ7dSKKRm5D1BRl7knF3C/mw99Feopd
T1MlyMMTvoEvmSPGzmqPLL+VrohS6KZiwpkO8ODE9IspIsigsDY31cpF7XEF3z2ZWlJo7kUWHcRn
HQI3GxS3MivFYqfRLlNTh2n/F95fEAR1kQ4wrvIzFLtbT1j1SycjIDIrKa7wfAOQB7ZfKPYTJqUj
VIqVgeKPNXKC1+09Uy7GRWrqkV6Dft7M0yUTpbBL2gDkCVImXS/yvYPVRPtOEYq085kPDcG1dEJt
N86sM0/Uc344wVAbFWjlzTm+cYg2p74jEQX1m5l+J5Y18oIP1dH/VYEpEGtBwAOIUhWkkK1iHHuE
IkMSS/SaP1l0PBXIQ0t5o5Q2XpJ8FPYipGlt09OdW2f55NzkmA0PZneHJr/MEGx39agVamTDKZA5
X74AiYPOVV01qJXEoIrk/TYsi6vSW7cjws4WfheO9kOdri+66sTwNfv0FxqM+jWmTRNywbdL+lxu
edE7vf+qHelE8KK+5BcAJfl15USm7kiXNqVWbXls8MIh3nLIYiosfMs4WoFy07a3ig3f1rlgsatk
K4R3DNKBWj3vGGXrEv3NKdR2d41OaJKpxDOS1Ss7nxKoooYtHKg163zonPySqo2WpS6jma1dRAzD
dalBYUsh8Om1sO4t6Ru4NMu++2E/Xphc2IzEeXB5Khyf7Nxu7hKkxm99iNgCEt6P7E3JM3Y86dI5
bJ3Qg9tPOTmqG7foPOnx6Bhzv51iIPQofQJ/GEcVXpAj+2c/ufwDg3lNJgKIGQOX/vZYpDcT/+u1
19rbOavlnZVo/+mrqGu2bpDx8oE72Ebr9dH259qFDVcEiexwDKGR65+qW+BoJUAdvThsQP/dmGCP
u8IqLJN1eTRKlDEbO54VLeLWe+L5L2Al3BAQNlwSTr23+zGXowtSFJUIdC9dnrtNuqxb4oBn7SUW
AOiI/ZXLRV+IuAV0jgzWCLYda5YAc/TDdfi+XdnwqOinC61s17hzODhEIfZbtZik5L0FYqdHd1M4
/LlF3bcW6DZfdAizYsPEhB8Nnb8XLVStTNav9lH+BRqpE+Yy3A632jBTBzFJNrhI9jFy6dE3RKwP
PWWtV/uRetAdZMGFYsoZGYbBpXjPkCGxp1BTgIP5lAy4MX2JPW/bwYL38M/jfZv/a3hCP7a+91U/
+RHUJKXWRdel1TL7ErvK6mmGZlCTlGI7KNgdLGE/2qGVuZ5Ig8fl9loVEmMBqXtoPLL9KE45nOt8
ZQjyVGPZ/p8M8jw3TLtPlgNeRX2/ohnSNh7Hup82hwdNO8ThLUuxSoWKoIb+4jnvD+Mqg8UvU60x
/a5fYHqTg3WeP8eZPH90Eeb4rKj4xX/HVsqqgVl2Xksa4qi4yXDBzhtHnseBj5oOm52OY+LhzD4E
UKUqL/rSmhhl1luv1JDL7/KMRfwNj0VTn47ir2Mpvfc/63P8p4Aq0TSlDl9JWzSfZBfO1Zz5lOMo
/ongM4rMkKBK0+SoO3PkfNiQso+02NFu5JPAF5gTpK7mkTGsohbKgXSVaeoYKW1ebwE9xNA89rwQ
mZr38Xo+aUQPvX7HBTHQbwZnc/426BNzyUdlnRrTw6J6vg70QYCmGo8tpQLU7DOg4JfsUxyjvrnn
h1lF5Jxk8sP6troE6cr4v6Mz+A2tTZ9W2lem7trYXKhwj2jvXhIXUp3KvM1w4QANhnLM066aozxH
5/9/a/lbydTFMmSFIu0bKyChCzrPYampS+pl7nfZldv3VZpi7LVn9O6/lUNW9KehTSZRYUN9/ldA
/oeebsuWSPHIH4F4nzZf9G5/c8lQ6AsovEoTenCDB3D/Zplj+jtkkjR08nj0R5rxHa+1kQf+UHYb
PRW1/ZoMQSok1GvKjHV/Av/mPBOPA8j9H2wS5ZFIwO4LI6TVd5AED/AM+ONti1qRH1hJQRlJ7Ic0
bBItEKQ5ye48C6AXWIunkA8GTnjH4ngZT9bJBRnteAFRb4Li4emD8GoDw2BGE/e49Xuc7pd0lSXI
OCixC7RVF0Olk/Z5kkz/QWCkmnnA9aH++eU32yMUkXNa/fU2MwrNcRW7OALh7zEDfOgOsrt2S5wT
4dDk2grdu2ZaZJq2iWKDqKa6mMypfRV98nmNF/fBMGv42P8ZUX1AHTSKH+4YjDtD6tymAD0Xm1JY
lqqYxI6MYji0mPqKgVraKsrYq0uruUxK/8AkcYZ/zyMYQoqyXQ0bMX3W1VPYtbFD23kYUcjk20i2
kQi9/k8zBrWvuKJrPUpG7PK69Irr3ay82MUaw+C1vpP28G0uoRx95ZgUf/3qR68p/OO4ByWlMkbi
t1TCicGpBfk/hB+IQHJIx9DQrVdLEOmIZ4c8LORFIgrkEU4m/eBj/Z/TVoYwRSz6LUdI81l7Fijf
EvZzrVapUd+Y6v/fFGLbwWe/kpALRyly2L9vggjzz8O0whbbf58kqAXmHPm4PpD55/ek5N09Zdai
f7bTtRW4QjQINYBCJllS/oyjuDO/hRlS9pYtcooiXX5jYzHvNdI6RKF+GRNqqF9D8l90hQ/gd4S5
2KT9G9hrQVIEoEA3pXx+AqkhkMGEG2DiB+0E4P5OuIQd0UHWT8fXFehoN5PD/x9XQ2CJI9dsxZ1p
gRCj/tKFxw84YD+KNSPXT6vJ1HNVtKRfEfeeEBFOa2ORihIx0uN/4zHdVDz/WvU6iLT7pV2vCgoN
zRvKGSTxrcD53VMDoQ16rbHVEYIoUdPd+ay18DgG/5nEbM11GZ7Y7pDI3+SVkpoksbhlvFzSKGmG
dSzy6pbkqK/M8CSc3gHpeiCOAd7Q5vqYmsizmuuV5bX3m30et9h48VZST+6gr4m+5ghVWeERSnrV
dBfLAYc/Z+9Mzie0ebmjtxw3m9HCiCKZ9uyhk1XEYiXrOzExMqWJqSC6LHTaSHe236mG4woHAFXE
Y0uQikHy4lDq/0W5K4GrxyEKhJlmI4fNqKLfUUozIKs11UnjGstrP+6nQR8NJvwpyIspTSCuubyF
UXnVjJBk0dqIUJmpxaDQSrPMJIv5SRLjwoaAJYYlx1OH+9T+EMy5SowG1RTjero7/Yzl15LtL+Kq
bC/JNy0ixImZ2F2wrvfmsC31psD4/hwinwYaUv15xxNMA30+G+SS+0oLWFeeiAuf93r48PdnSFDX
c4GZ+X94KqC+jHstmfIr/6UMF+Wccnf7bG33vDI/M3cgTwctFQgevibAw28FTv1bXXT5NWD0bEbl
n9ob19i2TNYCa4Jd+M4BIyE7GiLCEyM+CsuAM/fzzF4yI0XYa1/WRCncnXopAcEInFtacubr7NXQ
9fLpCl/+feW5lTPxQWomUXfAcbeKzYkPuyIWz1OgryVp14MO44W9ym4rQaiosKBNynQsSi6EBHcY
CuRmaw2EsH0Fn/GjL1Mk3Dg9KM3IbDGPRilrjPivBonzlZ+1eTuPnFJ6NkJr5tc7Dn6JVbQMehj6
f6tu4AkiC2iOLGMasHAx1giXKy/GOBcRFSisvaZWW9Gd6PKfsxXpiGtxws4ECW49C802MxCr/rRY
kkrqz4WYXnj3NPSr+D3MI5GIpmy+MHlFlsvm4JRbT/MF3sVzx3xVvI3lQynyECvVK4FWfAS9kZvV
Fnl+EL+f1+73x8KLCyYUSnLXix8GpSLokboq8xk162Rkiv1Aq3pIWBpE1f1vqx89LBkORUa5IKUa
pTzvIqIITwMvpivMWOA6dpsqYCxUAzTcAlnPwuSJZ7IFg8S51VqR4yHtjeMc8d7F05azM+wy1rW6
uok0+ZV2I9BjswAU4qy22CVi77cYYwzoGVxAxq57ks39BgKz4sOYHnqhHhF0sjZzW3F9G3jCTGN8
N9ucAyFWWYqBGfki8QCNacH5CYIjm/+ErdJmr0fb4gIx/Lp2eRTU6KXLCpDOuCbD2yGaBP9du7qc
oX6NKqHBRSDqeIvrYG64KCPP72gi8rhI1rmSvHyYMdakLrrnr0f54cgQYh2T2PuiNoNBFe99FDZE
fMT2NJhbeA2iow8MeLTJ2wmcN+Efqzob6j2yBagGfITGtjslyOfQ1U/ElG/bml2OQvtbqEcyssNv
HhFigseplvYiqqg5qumSTzKVkyGmP67hcxouw0cIpb0/NCkJX7YhpMMU2kk2+cqBLjd7shJXiwzW
Df2bO6j7kVqoiWEDytwvLXassj7yj7YixXIFK5gOLFa6b2ppYzzlFqIH8mwPlh3vCvQYhJ1+Sths
FHwOOsVkbwdurf5T1xzxsB3S1wSlTgxrK6a4YbR4ErpHG3BiStiCR1hMhR+D85j1Arf4LHUmms/W
n8e2pzV3QZg7UNr5xyLg7S0XI/iT2RsHLFp2mKlE1LfeSVlg4MndAP/jfwi+s0ejqSzsvh5xBjRW
q0IGdGB44rfHyUF9fASYPKfXOGA1Rc/JOOzFw6FA7i39tok0/VlOP+RKhGpIic0foDOVxqxIUs75
m7BZ1kyxboH9JefeQ5qR9Qmpq8XxuVinDINBqhYfzgtTv+Pkbdb68rgTTaIJMlJSHiewmK2ne34O
7StuHgXRH1eQ8WpqjfFiqIRC27CYccIT9WBiJSxSbEyjEsaXNA5+5PdNnS81czD8JTWCoNEneMQa
qHMVHsXxe8c3FPkOhhAhHZb4St+txz0eoJPh4IMAj/vck3DUwiLaIhquOfbLu2/pZ4OoFVkLjFDw
zmy15jDTjC+8ka6M/65p/YxpaP1uk+Uxzhs+cOw77xalx5AiwlaCb6WoAy9gH9E0HPFn+A34SDYF
YdaKGSHnaqh3rOsnkzbJFMwt6DzG8mTeSRZdUIy4p+yTXrN81mg4TSkyhQ35+aVSVw0i+ikiZUO8
OhdO1wHZfKCuD+6cCTNLIOOVgcX6libzU4sUgV+5SrZSakgvHSH01x2NGLK2tfR08EzVY/zXByuA
Q1kBbdViA1UCMcWW6taGKlgKIcucT/UpKwSvc2cSKmSoXSpKB+24h9P63qX+4cqJ7MR/1zkYqjKA
Z4OHtyqR11yyDX/FQ6eT/NXnfhZV5tBvElWKa2pYrGu4c3BdPfQHh6PbEFwjyNHyXyPaplFO8HaH
HFhAK+S/CP1mm4FxVmpd+ghy35XtI/JgChJMxBv0C+Ywc9M7ft8Eb91ClfQyCm8/T+WE5/T/QZXj
+MapWhvOqUjyOk6NHBoi+49JPNO/Ymhuo2ewRCVezIr3KZFLrMbwII+7tiXNjxbnjYMTjhDh995i
QeEMIJ9hna5/LsGRs0tpI13JrF5MnFt8AeV22vtrV0OfcBN5e5CgOSHROr4pI0K43mpL+0NHBJb/
ntXxKc4WB5Y9Y8hcj3llfv8vDrveO1xJdAPLRDzY0EHVfWddGy1oO3GaMDUkYnAXAvj7OdOKBYMd
E8az4h7Ioxe7BZiEyYy1m28ICpbEyFka9QbV6jVW+ax8vydRNw2bJlvuGU8lG1JfuhsUDCAaPEQY
RJpCHaPV5TrMmER468QwH8a52KYTYis1MKpP+6PTUQi2HFgTvdxwjvmAL490MsIOVuDp6nL6sPnT
xvSkob9Tt5n47s6PgyVZp6Ybffk7jodmJGwEG1Tk0JfIPd+DPlSfl/10CYojIR+6tG5Y4FikdWBH
j+XqiHtlCOZwZgt51FVYfS9DMAbjcAEq6qQhJuAsdwkPX5pCw4+wpV6zhQn0slJZQfRXngATd4HC
mJ9Ro4j425gXxD8+HKIck4VKSuiB5XNEiGqTcYOJJUzexlIw/fAaMTdl7J+Bqwisuic6VvMeb6yt
A8mGQ+JCi0Hd6SVLSoF8IbBvJwVp0HJMPIZwBUTXAfz8kzQyVIuq0lQpszkniKOLWf0Qr9bx9/o6
JdwwwmEIzF33WCF3xbCGEAdK2wj7dbO928dXNuxl5zPAg00OXs9f1B6pJjnEMG5XjqATSbgnxLvS
UQUYv1scGly53jrop4sdA59UQ7edAJ2jJRx2gUsxDWZYC8CHXzKbuSL0sw/d+Pttl/wa1Mv/WFTC
Vn07JEYtWmI+kpGP/6TCHYhzgiMXb9LARgxyAsQcs87WXydTCI22mH+IPUsLTSBuLT+HR4lsfLHL
njfaDbHb2VLxsbb74RIbg3L/7YFABrIq04nn/fw3xMnvGwAhUTFjSYiqaaSzVkwfmSWXIOp9BBnK
vXUOZwonbled+ynM4ZmbjRWx1HYV4ksOh1JUy/kch7J9RydBhLCDF7wqyRwayoBguj22HUtqGOvQ
c0FNlyTm0rBR0CwpjoO1e2QvHo1FVuOPAOPj8l+6/FaKLvIZEBTMbAJWb7I41XwPU4E/hxqHqTCk
uaBnNPiTcdSgo5XYYQNxcgSgPSVlfoYXRNZVqyxatzpThqCW9IP1yPBZRCm8ltPZe87IPlCJnM8F
cnJ6ofL4AAge4K0qoLXnpRq9qPVxiu49IJCP2GRNvF7Tvlk/qLBMFGLNCIjAn77QXzOWyFAKySig
XVZ5KMMtSOiIUN910GepsZJIIu4NP2zOZI0aYQwCViLr4zFoEvkpSucpzX/d7HiU9sH4D90Urv14
VXWVcb3CzvXr+GXN+Trbnm/Mkv84/P7qMpHuI7D8Q8ZH+bB5rJdzvmCh+oGw1bJz54mhrRVHv/i8
LQJOh4bGdMYn157M9bEmlhhn92c+5w+p0noyMjdx/8FiRzvNUwwfWl7N1rklKxxan3r0s1PS59cv
kxl3SkrGPsnghMnDbDd7Gb7d8XOVICWJ8E3eawiP4PxnjrCj/jdCSFwM/kjvL6So6eOJQ6AD2M7/
nB0gEFHD2xBOOyNpmhe/jB2FBryBUehIURuMPbGcQnEV1Gi/44vpsfp+pyunI9aLJqeL+fV6h+R4
3UuNvHJ28QK52iP+5eH/3PSjcZzj3u8HuAlpsqYsyct1/VThcXN03ppqDcRSP683aRpBVTSR15X7
75vj9CrzfTgsqIXfLvTndg6Ivmi0NwaleAawyi5U17y7NUCSft0N0XvnHD90zIFjU9V0lgpAUgWv
mhad9gxd/T2KRtYd+0mrCHdcEjHHYLla+LxRDcZb7aiDIdhnXFOXABHxDelO4kPhWPHSeUYX4H6/
AZ/VKusXChiIS9WCC828FMxkAjPMHGxnpOl4E9G0JRwJv5osSSH3Yl2QSa20kNjdv2qfiqLUEvo4
5mrOX9cGuldEl4aar70M0V/VWZxCaXdxujkbMmOv/wSdfgfB07DsXvmnx380uNuUseFtt9StoEzm
RWlP1+aJHDLH56Db1KP71hELZywKbPaAdK4QfVYT5C8UUTs1E9p3QhPhAh9R6fx/yTAtlOIxPSJr
b2LgHrQm7ybVAoRw1F+u37ZzxmivIYiMXAQagF3DWGCu4qfFpSkdhsvEtmWGFHsL1FAHzEBSmIUT
rh+o8toG2g9+4yNILWdik/b59EOmapket0P32oCcJRdV24wK9G+vZc/PXn2Ei0JIeUWV6jHT8IXg
eiWvJYiHqnSyXq0Cu2TXdniCmc6Z0Cpo1HSFVnfBNgtvvTRYYJEJVd7DOEzFLACHuzsGl/lQGSya
dTONTXwdXTBb5iy5iFPg5cLHm37EqCA+sAO424QCKKfnnYKFitnBHlwVXcw1jIJ+nqywerxMf8Be
ia2AHuKNWa7UXKVwqRs9XXOS0v38ON7jsd89dncJsFN+GabUVou5PqlkFe/nudfCnozWQ4zKmSFA
quX/oNlFht8Nhx6/w/Dm0kJAhsKeMYHr77blpMiu6u3vkqZhJGra5zFQV9QpGnXzKzyD0+ahEDvS
r0X3e6VOqLMBu0K0q3UkHonfz0DxyeR28nEEddgbNfwihTpuq92pewV+uBVdC5EurxRQLw10O5UN
plh7UYcJ+gjFnDTnzXfBtveXcgY7RRd7lrb/Oc4+2SdJspGHuHFER9rj1T8/cOpTOuuF9rzSohwh
8Sa8LV3eMxPF4nt322KIE4tfDYeGUw1Y2DEFCln2NnUZOgZ+z2ELOJ6JAtKJgpSy0scTNBBC4yv/
VoXvPOg9p4H/ajDLf8ozCMGIVRXt7BeD9bhxzk2N2jitUPmsr4sKvdgO/Dcui8x70kigmtsEihRy
dt4Sm9nQGIe/Ii8p97MiLNG1QIQg1EgJoG9Wo56Ed5QVL3CSTQaJrkrrhHYXAzEi+cNX5z5GrN8/
h/2gUNuBkStGgR/heJPKlsN4ymrtnpAJo4xgWI2l8MZPlMIxqhrkVl9rLYueBAW5lIS9GGecQGMS
0FYh+LIvZz/cNqmuAKEbvEO6BJypjsOxi+XxbFybpyZesNnEMLTA8wsrKtFpoV4nDwRt8tDfE/y+
mlHuleDnDdIPPDXM/vDgTxfWI2Yne/xV9/1qj2aCM91vi+nO6cWTS3q8r6SU6A/UMQ5CZ1mGvkxz
10mpOieFF2z/uzXpwmLpzsOYZgwJT0rlnixnzb/GWfHuSzAeDjodh1ucB8/EjcHAEvAL/L2r3LC9
TjKlXjjVFhfU5jKg5NLV7FB8Kx6zo+CMesJ6L2Yc9kwPWfgj5y6ZvG5RLq8eDXvbX+LutuZdwxCd
ck8lB+84i/O/+FwL0bUdXFxex0dn0FSwYwSQnTNXIy8NFewPOuIn8EQB9iYxPBVVVZux2PLl8t7L
Bd4YTRXZgpOkwBKCAnpVB1Z9NaGq8Ex9xTmWuwbqIq4IFlrfDyS0QQp3IoHiI0lrCed1HbOHwNUt
MMvTMQqXxhJw7FJSSw5yrnGD1Yx/TpUDJdgeNYuAHLgIxRH2v4ZvVjuSyTENiNrLayMfFfa+B31V
EzNNXB1xQ5sAi8+S+I0cGBvoQF+UjR0MR2XOcVNpWoxyOs4aDiHo24LDQHO/4vWF3AVSc9H7m8sf
Wxi7L4W2maEXiONlconJ6ukiWR+ipl2hVjNw877ylIozmj0uoqaqFN6REDOVm4Y3wczIf3VQXLm8
h2iUmr0xXq/pCgibjhHsEejiZoUE4O7T8cIho+JW84afa0rZejNsmgpunXCvvprrn23LDurAIY3S
g0oDJ+hnGcIUrx0sZV7bN7B5vDoovsW42Pwd+DKIHNC6Dx5+vm0J9qJ5BzWBq45UihP2or6stXmJ
a+cEIjc9wWlmlAZ8k1gZQJWzzKb0Hom9tkXrTmwZBM1QDb5XZZegGpVZIfsplL0ChvqUSXYhnsAB
hH+XkQC9o6MtfWitpw0wT2Vc8CC/fgJTP2UuVfCT/OyF5OMg+z+7KuYXW/pvMxNHpy4tH/n+pypl
u8diLY+08NtTSr6NpBItZ50f7X7pFszszT4lVLuh68V5hhUP5K4x59F+8Ae38vjczCy7dOYjN2On
nmyrSNWR6hZRm3imJ76x8RQGz2RGXUSxM/7RW/A8S6gxB2goJnTXyJePTB7tz6pc/o1So/BGf7A2
VXEiSl+NUPFCT59cRadn4ywDPNIm8grBDmC2r+PvCV1clGuD1BwPqPaaazy4JxmBuQUO3KF6uxGc
Q+Gd77EEu3oosjRiv2LWT6CIlSJ7IIDiVJkdM4THc3nPHANPnVNIjxLgKl4gDeOz3eMjLtAjajfw
O43nNjiIZE5qFZLOsWcxr9A5lcAUq1nMyyO7vD3UYat01euLK9Eu9iJJXoIfwhV6ehu2MW87X+w/
EN3T5FJsnMIOFfupbkZkULGRx1XMhr5aUm8PWzgDOpRmMKOLqJfF9UYabsGOoGDFSmjXdZUkQZlV
wmpW6CGYMYfwKSK710mRhXPkZYQ9It827oYrs8icek5wX+WkQHhk7Mp9AEeNtjENvrTLiRUkud4s
8nye+KbW50+H58NrpPehRI0OBBKLzbNAeIBBiz5gRrSNlBilG7kdJNgWNy6OuItUzX7qKQmco2pU
i7J8jA01yL/wb7IM0xx9Jir5CTP20THr8KCpD/ZIkDf1h4jWTKIvgdBbDTHwCyCY00bk49WeithV
PoYxI5jtktPWFvnVI40336Ecc0l2+bJALdHsfFkyMlqZ852qykvLfDsNJYqc7CmAhiKs66ubSGq4
BS8/n6EAKibemwZWtY+e11f3mA8fFgGbxy9Zg07EolxJALjD+q36hwOg5pich7icFtn9iLP5twi9
ULF+G28iOxUwfv4/6z9LzhfFDMy2tXscv8WmReUCRVYVi0kyzPuFdOFRSJsAtCMQqs2NAq+Vr5i2
0SyqyelN/BNbQkVylrbbzCwZguKzLcAp215FWV5kyYNXeLRSAXI6frWX7OR8E8nP61ZaBl+g+/ql
0FiIpGA/tXF8FbHj10zcaDKhSr0cK851XeKI/qcONrE7QYsXOCd0cXTa94WE2f47iOcjDLaBg0q3
znIKUs/0uIp1XWxG+X/DdcOI27gq/Q9P4PetlBzTJVaBni7zMrmQtu1epi+BELKvhmYcDkNRIa03
OeX8PnXB6hhbQNL1pKkWzkfboeB0g9ZpY2qxbE60AZcmu1GLCmcjPc9PmyvwmX6IH+/boCYsLzy7
0UNlV0zkjbyqnVPPNPZXieHxDgie2D0wqlReHCmckJ5YTMCQm2uR2hBiZof/Vqq1L9ohgaKv/D1l
j4X59K4/tPWcACr5oMsyv23Ps8k4+q21lhTbiZx3PP0ab7LYKcMLMrXDs06D2XzLYtlq6EAFSkA6
Cr4EJ5MTqPqg8XZP6bnPFRzdTemouWw3kClIy0IVSohI6ikaU68o+nd1TOFfugJA085w7vpOtXnX
TXiXf305luxe35bRQtHdOAHJMMrXvpd0p8fRflkBNOUhWPLlQwg4o1rkxAvODBQCr+IM6rUpVd00
I45sCjN05abmpSFsXquYcea7M1gnKnL6nmD4q2dJn8t821JI7iqJsNzEC/TMATjxP3DNbRIOqp7Q
3rEOgo2KB7ZKquapfKVR1TCAgNjeTBcDQJ148nPm7bfOqr1ihBPrYLnZ6jryLNQBdu54HkXbTkkC
zfmNaIg1TraVAI8mawWNZVCMyJG3VBg/mX9zg2/K+OFS3GnC7TTY8CkMF4gIWnLrg29NL8VHxFGV
/N1E/GV4j4doAQ8w47lQMEb3T87KDYIZBXfcWPqFxDuolsGReMDPQIOs5kcsz9xpQSdPDp5wCbOu
/QfeW294xE2PGPQsD4dsNVaMA4s1E5Mcg8p+jKkpxw17ijlydcXycZsFqPsjITylv6hjnP9WYIWI
CjAndAOXCzVCZMTrRp1a6yaVGzrWEa/z6LQP3dhdZCrmG500VqiAChDkOieGV62aUu/0ldALsgrM
QAQYt3NI/iFtvPeS2aPAvIXNbD6+f6WrF5qdF/gDUbe8V8z1fXB9HEwhgxk+B/iOXSxjBF1/hGsY
ORkgQgij9M5IuZrZmxTzPyC6jI4UZMB0lOx7ueE1mRWn+sOtT23FkPOTr+zxQMajh2bhx0BPnbyq
LTU/I9CHHbO1NIM/2PG4JU8nP9NZWvxuoEyqnX2xE3HS9uDkMydPJOlH/Dk2+liXTydnvizjI3aJ
1XVa/xcZSvA5/FW0qrQrs7Uso8eswH4xxRV9OUwn9o1VTfHmM6hO0g2O3olzyvr7ctIx9ZlV1Miw
S0nM20DT8n15v/R4bz0j0J/NmbzbXDJl044bbwP/+l6vjOyL6W7Qj8DuXPEblcbdlI7RKOE51Y/1
CSUSWDq2DquVoLpKS46pNrBpW8Ih8luwg1ys/sESwd68wYdU/CiZD6fdrtwJYvCQFSd1FHKlfqu1
wYOB65Tz58b7ISy9tgYK7FeNy+o/yutYnjQCFDcCO5Isb7VlHApOjZ0FmLSrjJiO/8UH/sB9cYiX
D9wH3l4b8Eq3f0UnNLdfCQHXVvBkBQLxn+i9qiGSpfhyphC+vR2U5oL3s29gjdln9ZozkQtgLotN
5QL3z3nBJKnOgCe+4OaY6bGwr6qaPyFxfJmN6znrBjjTNBM2VgRJ0A73o4b6G+veUcXv+qbbnyNP
iswPKxHPLnv9MVvfURvnnUz68D9tsKtPAjLND9kkhtPix2oCZpXwaFzOHciCVrCdddClAP8Ty/Sf
2Tk38BZSHF3hr0LDO8aBrFfa5BajpAiZfWstjcvYpNAu1V2g8umz2OVt/b8lcU65r1V/BK00GAcR
FcKadge24pEbzbXHej5qzL2lF+06+yUvKtvBOyEmMdazTMNZishZZEjZqKzPb5BRqVDIoAhfT85/
JawfVqWvJ8dB+NKTN9rCfhlYLTJgkLQ0zAtP/dG+Wxj4NsAKysu/ThzgtevUnbGqmhKWiIPu2dlR
6rP7tG40RM920sfSjTTleOJ6bV7b65imjhyQmJYW37Y0gKm23DoxxU3SqaA89vKBBM0ZfZcz698v
2lQtC8Jak+EJjZ9eqLpX+gBf7QJzCDOgTqBPEb5ou6kqVvJTOfhU+LXIaWn6z2JTT15IqkKKDEK3
SXSwrm890ghT2rlrwE1dLJvLtcuNiSEHZp/IG14vU6orN7SxMQZSdkMcp0G6JJMSOAtpXWD6+oz4
zG06AHQ4vZ7mtiVTI0dYVNCiRu8m2uNWC8vge3fPYpG96aa6qqone+VnZ1QBAbEdPcg17uBcFLxT
qS8PsVEN7vMuAkyGGAE3cEE0wZZn9QPjk9HyOonXTbAPDG55EjOX+cwk6znunl3qUdT3M/kR0K+u
fHKgN6StD2I3ZbBHveQ2qexZ0CCwRhsTliNXijmAt8gqjAcWRNzCuqK/bsDFSGLQJA8EzzsOcFAi
d6JNWCadM6QuHKTQOX3G2TxeU9WZLjqe2jaUk6RdDAzfTl1cvD2kh/OKiz+QvGn240QIPFe3WKAN
FQCvGrQplt71H2K0qtKpcHFOz0GS9NEFUQEP5P3u+G9DM6FQU3IwOnRWYwuGoNYG9N8069fotiFn
oFAdI4V9s8r+sq5FSBwg6YQHOpjYSdy2r9aMfQj7ft8FxvvQoKMuIaJIb5ZiMQw5TZczv69lmwPZ
K+7pnn4nPm6TdkKZUOaA3OahdSzmFqUoXgVohz2GP9BrnjQSGsDzhU/tNdCdwLeWbzTbywQm/xKu
xucw6svJABgQZCMf3S6Mv0aiVFXf4iFsq+q5WBviI8RQ2BYeE5eZF9KYWTy9ga97McbOZ7JtkJl5
w/DW835c/A6tsG4CehZjl/ZvC2Vjmy2upTQqEyvet3AMtaSsBkh0jRvXGg+ofgxiSmCtXafDplf5
tBScpun6eZvPJX7RvgF6efhLnHRghw0ENhWYNEPjJ0Yla4JNSZgVeLZy9T0G1p7JyHLjlJoeGfFF
R/xpnuekUGBYUvPCQtR60HU6DLDM4SlEMBrwdF47HFPC52yPAQYN1hAfc+GHRcNOK3FTkMicfmPu
7yfPgcy1DAVzwfcKN9pjhE+pwOOPixfCFO2AhBs1Mdw28iGK5tjlatLhhuR+leNekd0jP1gL0D/5
GckSrFQHZoDKVNONH6l+QbYpSVMMHZna+k/GhnQmTmGJk659zdv+Zr85kiB22DroU/QUm2Cnk5Xg
7abhL3u/jek0MnzMJhpOZ/LXjEtkXDn+Kx+smBVJRMf+wdVY0BOotlkhdtuKouAjKHGUkZD79pe9
Hppwz3Xv5lqi2JTBY9ut3Ay2R4ijeq69X9kGJNxZFfT/7KhlkcWxI3ABqWUhW0SuIPTubMjH+Fm3
7V/ZQBbtbk2zugXpGYcjfwDvHsuAf6y8SQm33F9TNky6pN2ymBfeNx77arbCrwy+hoB118ORHRjp
PBzdjTukcoZjiSQ6LtLPPhGgyxxYj4TCTBow7sJuYcMH5RIbG3u3zjzEMxIwm6KdHGv10N9Vqg+6
30EJvKJopCE3TOOSdSdaJX1IBK5mSHAVBXHFWrzPrPkr/yYDsT9sUuxUiLSdbt3ocR/TkHiaKv0S
SeyXv6YcgwBafqLRnc9IqcrHCOEPSWDC3EHqHB5tKXCk3RzundDCmd6CDE1xWAMLM6fapd/w0CFk
rzpGgOsTRcwFwIKMGDjxUIFAwizg5lpgGIGchdOX55UtXdSyKebMJZzd2jWYPk5apnh/J51YmCG9
DK0xZMUai8eZ2IrOYuvg0kM8k3QKNu/A8OEEq3vkRGjyXwqEukBs+vHnqi/9qGoF/C79Je0FQkvd
gZce2meJ9de0pCTOm500CZ1VZkRp9Tue4w208hZulPskl6h9gjtY67ScV/gXCemW8JlsfRqKcZdP
ErTbPPCpjmDN5HMemiED/z5XNXkDTI6sOR8Uo0ZfjF8vYccOKIOV9v/YIefHgta4Lz3i3ZOaIpm0
PO+YPjsUyBdBRUCAVP1W2RRud2j22ccZGwF/IVhlJZv8MLDQYke/0UBFUq2I1tOK8rvESTwCPqqZ
7LzyIFlbi8UnfVDy0cWojyXzUk6/lXmIAbgZYbkewsgRXJXrg1tJh8v8pN9h4EuiH6dA5fTGKBiX
+BNjjol3VnLlsV9d2XJrkufG2CJ1WmMQbDwR171ydTHaMMepags2bW9TUybnwQfXBJiVV1iDTXQS
SNJFV0sko4oen73nHEYEuJsmOGMxRaUqLvCOZFQ652QRZzCgoSzAc05oDHyjlvUWrZViXEfY6gn2
S+p9wtB2zD/yA8s2f96cf2zaSPWov5wJX5e8CiKhajy2bM5vA+Ftmw483fJblys8R0KK4hOHBHhK
t7DX6q3JqOgIOHFeOJUPVUgfADE7r7u8tJhopRBtdBK2NwveL/ngeqAZ59zwhCQpHA4zh0hGnL9x
TYnafLI0skkaUFxp9lwzivrZDJjRyUR4uwR5Y73k1vDLmOkFqY+CQibxkv2dyw7HLjpENdsQl098
b4Z0zbcXkjikFdTZleWzbw79Cci18RWeOKqWVyEtF6IIjtS7m27d+uQ3VLrzghMXl21qcK6WbMjm
m0W9yWhIUgIuUIM7O/4N67N9UJ99hUlmllZjcNTovtv/SbnJ2Fz+S/5SNj6ivxitG7Pp42NuuYzN
NG6yU1J1o+lMEZQse11HrIRJpxjVgvSsxL+5eXuAzbhel2ycQGAQtgQ6axPIyZ0xiXIun5ktthmA
srfhBmbTTMYnXH2NblObgUOWUW6LBvdp4DoWxfFXm54/b/7Yihh+4fgNmC1HSuPXDbUBB6qmad4Y
YarJzoz/UakK1m4d0FjiQvl9QS2zuzIfKWfDQU2nOJfQHDdieipj8OD6alMjuPWIOGVDSMVb/Fwk
ARnD5ykEsJ4Zn5t9Ajh+1CMYxG5uoINpxiqvk4DXy1YtM1tQf6itkIvYdbCffWERvkBbEr99SZuK
jixcPhq9xPkyn8Pki/OVIi5YVdxRCnpTyr/+4BuAuU8RPSQLzH+/IhZ80xEOtTnLW8YGq6sqM+CQ
G2XVciN4Q7kMPClHzaCCIi0/U5Fi8xW4jOV6P+/L6M5N1cl+3jFrax87KNF9YrYF2HhwvjSKRDRK
OihwyxyjWSK6HQt++MclRUDEIaTQr5EaGQjtAtJMbXtG6uFG9nENezM+5X55yYJJ+ZcfqsfOobwU
W2xj2AVpyktX8pcPvMVP6cXARxDgWEcMLNOObgv0DsHgLFhZr4IIWzOy/NKvMAVS1XvvnrtQ/JJ6
nBEuttOc/eVY9FeI3BRtWfpPwSHiCdBJCHrd2gSlAR2KTlrKX4KYCI+NdwxyUL6+dj3ajgnJjFYF
Tn0KRRvnMdpDnYBOTqgNqQjSzrN1+AZwfCU/MqaDHHqYN4BFvRSodG1IUAXbvCHUNS8jGB9ExuS6
Nl4UQ6qSc2OQEAut82ZAxswqzUl/yaq4aBAr6MV4XpFhvZh1enXgxaIs+Dt3jun8UmGsJAEYomqS
OzlxzvMIDkAjZ4DJlG1RNQ2sNqzNWjCSflSYujY1td0ZCuPXha8Zahk203hx+Ckc3dFcZ3e/wLo0
4ksfOlnTCjfvPmsSm9AdwxCOGFHGYibDxeytHhjsi8Bk4Crtwqg7YpfvxLbVMaf3/IxWb21/G0q4
pyOxPE0Lxt8OwqJB2MT3fao454MxE3YPzhStIxdSZj/wwf0d2UI+d0PGVmRvGDc9ejRpa9yhnkSH
PNKkS1Pq5gCwiMfxGGDkALyxpHie/LxZ1PSepBEx8vmHagfOzT4y35WwBhjyFY31o/IRnrsZwGKr
JMH70RD2RrqsGubPRZzazZWjkMIyBtcR1/yKBxwTdIb77FuxcPjlZsQD1yb1ys6yPykS/+K+lGa5
M4UagjdiBS711lLGMkcJ6uOZpO9Xsstwvb4N1rl0XnDlNW6foTMKzBIURbFfMdpjj6efahPOSsKq
qsGfT945H0i7in4q+M07kRGxK/GWXaMtBWVrV0Dux9s0W5lSlRkI10jInnMtFLd4B4/jbCKdHhF2
Tu3T6aKGH/z8klLRnOUP3wO3uIIwwcafJOFV9qk2Yutd0HUntrL823Krgq8r2vewgsxuDg/Xp+23
jmAKm8EddEBSqbqum4cTkWlMnUEm+ST1Ukwe4wZeoD4mgsIz9GeA94dgHHckqVpLYOHOUqnkm/Fs
rOM0QKyV2SPJss/7JkxABgM1aHR29ZoS2ISytsCwQHCH9TvwhLhfw0CKYpaDYaPSLUsEvOjmv++j
DkBDaPO2fXQpf0FboK375WQmbmVsCkJlOUPaJ0L4u8FvQIvO0pUGreohBp1woOt9sLGMEYaFNULc
MN+SKwoksKhycpyyGPmCwS3YygH17Zjkeg9WY8u2C9QpxwlvQSMcgeFjbDxra8NUFNXInqWujSiq
O3bW3Q7y4qiOMMFwTpCThsURplg6KDGjvdk9iT2JJlk5x+gbFlD5bPM4rxoywc1htJTMFu8FQk2P
rhUmft0Ot+mnnYxGrzvNB848zimtjGZCEHYFpShO5kvguP6sIGn/2jwisd89kogcKH2n96Mb34lL
TbASeZM44mRWRnJbdx2JvNytmYDSjaztCV+LDldGIlbuJxVFz/s6xnPiTKCXPnNW03ht5ixDvnK1
Cfs/4mmCimzkm07abQS0g41UbFYD3t2iQZpnkmgC+Y1Ae3IzTeZkO1tNEVrR/Kfg+340Z8xiF9Ra
YScrWlseOG71L3YuMN8SHD158/pzyNxLpMK4wp0F0oeJUxNDTkBJYdQfnJjVZluYvnYe5A1tlqWB
BciphLlLdtW4XNufK0dXzFNh9vd+YBXRf/qzrt4UH5UGv8RSuIC6yyyPW0SYrOkmyHO7kM3fbn8l
/PFDjSBqLJVDM3bv066LsP5IYm5kfQHQyct390fZkaf6kS71YnEMGKEmmG/wXJQ2HehrLVoO2Mj0
NyyyQzNJU6PM69CQ412x4+XR3DT4dwDIbzUTD5j9rXyKstBJ4MiiIngiQ2lWKCAfBh7I+m5IWPx/
IA2vHDCYdFz8ehKUXeZOWawzrmvzEHkNxEOlgf03J92AxVFRAa3W1iR+Ulk2kZ6QC/fUArycB3NK
wq8LQiBSG2QwdKsRsfdwJGoQsOqQLArrUmLV9hdQQlGSEz1VdZAVrxbeaOyqfEODGgUh66st2bVL
Fu/PxmFA1G4DCQMgkhFQDDnTImshYYmIHeAHbzras88xPyQv6mjbj/Lztqw24NFSK++LcvKSR5Z8
dmFBt8FyUBuVjRsDj+4KnAZd1InrK+fQx04Ap4qzB0zpu2USGbNseZVSbIYAbxM8XUlrCcPSSEtv
3XV3KJuTNvUpnkdwuCfnotfXTZmnvzDvB+sDwtyUCTmWWJWFnlzg9JmJWglDFYbyNP5FI9lhUenw
zRGe1DgT9JY6DZjqVnj8oxx4ZJsGPgJNQRrIVN45Fo+ONXJmYCZoIVIEGtcdtXdWCRRVRgskCLp0
nm2JzWLK+0kGl/Elbdv+jgg2sUulSMGdHC885D4an8kLIhrCnE4Gmm6GTScIfy+MIiDmx1noZuzv
Z0aDX2oRpcPuptZyClQOp/mE5gZr/w7A9e00w7J7harSOfbsraMHx5cpKvTsca2Oriu4Pg/hvFiq
r6MBRirdNFutF/R/1bNwr2pLQCpvWhdVyaTPkQz0q85c99uavqQK3Uecvr2vPcIZ7+oTjslmVGJ9
KQjFIhBW4iBaof98BabwrzyNMQRU1IhDY/gciOE0zc/l/zBJnTznU+AlZGu8J4M5T5rqmW4iB/AA
t8gRbHcDCOoB42SkLJbUV2xR1hpEeAqPbQWOZQvI+X5L9jodWXXp4DXJh2ln+MxoArclTUFMIfcP
EwPhuTsbUF6duMotctZhCS41koi3cRiVuwg4a2HSlTZ+NLI5jZE9I/GqZQ1sWNh46E33iMwbVN0z
8VNvn2ieI4DVh63ulB/SXvbigJ4cHf5q9Cc43m5YaHBVkhSPQXQ6GPBQQt6N4wyuZbuqmDE7WbDY
9PHy/lep49zHxJ36KWBpiB9qLfPlTc5w7WHbGNFzMl/dKiwyolqTHgH/GL3X7pz/dZhTWI4Sb/fu
KihZFd1jKImpnZTpVpi6Tt/GywKSvxauURab3UI0AYGqOpoRzfmVRLW5/T6O+njCtCcuWcAch84T
x3t6CJLyzP7pbIHiPBlSzDatLErGDKej9HjoIfBIrEBXUnbQvRFtHtTXllPNpxe46/bjxEi/EDF/
CeF2oKvZFAYTT5eztTfvH8m0P4o/qAtkgTF/Tj/SpcwuzfH4RIIiMJejvSvCAh75/WtyEWV9bw/M
vUP37O5IH8vXYPM68wPBlr//qbq22Nbk9xzIrNuYjRYHVkBAsIoF30SrSnbtWOMX+j4aALi9TzZP
sqon5YLoiFPThe8dZByWvi4seQM+HDKg6hfGqSQYrW6PcJY6171gWOoPomqxJOoQb/2Xr8N7+8GT
fm8cUF7G0azI8JlKAmoC7GZUmoybwIjI/ds9LJsoW3ZeLtBS5MG69VZPOHz8eB3+RJXjptuG/O1X
kbP2rPUuPocB2xl1Dbe58wIBXxE8dO15zQjF4LKzWFPF+12UPKY9dAc1tZ5fJihGbBrfYYB6QK2/
AtVXXytlsfK5N+fpW7IUdQW3QY/FuA2EZWYzbkSmxLgvvxVDo7BKU/3ClIXSgi95BoXZ8D6B0B5i
4V4yt7zDeCrdYLNl4l7zNThoiyAaAvyutbiD0qpl3kNBhPKT5ekYAf7S8m7qSAOOE0Abt4Vad7mh
xGy/xW4dH7Bj9DDB+nKwRft9G8Nn/Bbj4MDrx3KVZwqY22y5ItHpm06dezLQlHW9O57LwNEwUmg0
Y96idJYysmD39oAvI6iKu3gIQEuEHHhQr2Fz+0LnNLWuofxgPIDuGPARFi14wrRX9Gbe3vQguLp8
Gf6nXvyU9Ry0rO1IAVnHgvwFD1EkX/StkSpPME3At67D5ptl1gf8+pf4JrgOWf3vpdfFWJ/OFJgy
cqawX50JrRPXL1euRjFPpbOwsoWDqMzXC2c0+0DUgqiBSAwqHatjU4KxCEDIzm0tzUuDyO6y3j9o
nhPY6w+lV+qJi3f0dK3Bik8U/AFiWgo+i0Zwsh6rl9hmV8JCl7nrjccOplDh/SMw73jfPKmsJE/X
7tJzEsz9mXGiCouJ9t2P4pK00n1V70CO2aiFM0SL7fHnPpl0a+rUNR2DlIwBsyglaO5Wg0y5kjob
5Dc+PYuM/PcMfRyc6GHS//oWBNUPn8f2R0lnTPe446bXnh/b6sq8HwMW62Fdd2uqnN4WSJ+XdY6n
T44nvfm1skm7EmdfjPqmhE7PTCGsEp1+qvb1WVVhTMbqnaMXqMSZ1vrBWxTwM1A4WrwTsFtPjFO2
I3S2Z/7AnKeNw4Hs6eEJ5E7mTnrs/dYLifGTigcH5ETKb7dJSIY3I+68/FWDeIE5sD2rxC6rkMue
ClYfN+z58/ZzvbjSD4mgfr9y3ReZwpH96lsajC7OUacbOdkubvbsCeN48GBhxNSsx7ay6cxea6rO
iVgg8ie5PhMt2tr31ICG9wBKwzzaoi0hFBZ2PEevlYgdcTLXgI8qlPyRvm+jztKHJEqmghdMDQ0o
qGOVp+RdQBCeEd0ZQYjHTPS28iln9MQtQmiGi+kY9zl6Lb+6/cy6OI2fkjV/uGjkyzUY0z6xseqz
SaZ5PmEL/KbLPrfS8V0ZutsPBnRKzAnuFbZJtOuRrgvbEHEFKB8M4o0eMF5+FJJJjTtL6JMoTz5o
R3f8XPg5UMQZsRv8/OI2cpT7BYBh8eAJL1e8Ct+ZYKWv+YNNKIv9gpDIuJyMCwo2+SsoZ6sSdP96
wTgjgpIfa6DceT2ehI2eQSTMpsGvrFX2zwvxG7RXvkDlkwU93SNYbUGWXrdx3JP/0FEuZIwgRba5
IQ+zQioIFXPYomjt2fP8vduuQ8PyGRqmkhZHICHBN9iQfg0KP4l/v577txwpPEwImXqQbYDel+t1
4kKHAVmm3lPUXEVImVEifFIMw9aeitMQ3DFqLLAke4wbHXKMHvIPrpRiW58Rrz7L5713XtAbsBy9
0UC5TpSRvZ17tpwwI5AwEeNdIza0JsfynOhUxRRrGEByX2nGOO/UQpcjh38G7CpslzVvLSdDmnNL
7iEqgLgsfLRhPGivAHJCfDaZAa/Bw4vRLNuZ2DoNdMkwXH8kWPzTCtFKFH9txkbwO7l1qUfwUOKb
LJ9E1h/zD3ywhOzGIk+W9g7DuOwtbhDJtAgiZCxOhv1FdxioeSThdL6pyOKkkqzcTSkF4BLOy4XQ
x85NmgVZjuiad4fdtPLLevnb9JunrLFNTyF7izwQMwhwI4yiAxIA5Woar7ShL8XBlsDdB6H/uRQK
e8RacKSjNLpT/FmsQZn6ZO7ABrHpGMlh0MT7wQiB2Gy9x7SM1Vyg6QyVWU+4jgLa+R23wOm1fTaC
VH2gbsAYgFYk+PDM01Y2bJX6SJa/pFSAqa1Y8KxchfF6yp7mBHlUI2HCbcH6X8s1CayL1NzGNCDs
/ENE9R8IvLVGEP3ePTB9ha6cNrkqCWxu6vX5tUMxdAYzD63M2wu+iy1MkzuGxN5hVBCveFNZ49e2
PXGi8lS6Vae0pKHuMtIIyhDNfTimPINAzoLqTSywpjE9muX9jn0PfcaHDG1JVtyJWR8p5b7ncf0w
OUgVzhrX9KXyuqXFWG6ChxKq/zeg39+RUdxEgS8ek+4AFcvlQe6cfoUbRZ4kZ7huJrOGoGUjMC2l
xTpZ2d3W3Gfc5PcMOOWITcGRLAsAG3fMbsdony+xu/RztxssU0y5fWqK6NUXeGu7Vo5Ga8LCEpp1
iFsSJJeMKsAwM1lfLyz7nBJVVcmqnLapRjUQeGYR+Xl4jDLIKZV891HmyQotHwG31+x9PU04tKId
/WpvxGKn48YhibyFYudYJdAH9y2wO12IX+/KO5Sz9nlg8H9Z9CTXS6SkrvuqMdtZGJSfFzha/P9Y
MImMLD4ZiRxJjMntQm3x+DiXsrkFjjzB3Rwkl97Vd3yMwW+YmkbAIrt3YeH8cJIZk04MppzEUpKa
G2EMsf1ueIQlrbbzJnGFLG3vyk7RU2yDY8JhkOe8n6sHdleHaFasQCk1sbWFBaxkUq7wPE7GnYzD
S/fCKlTh2pOCcHnoZ5LrnJmBAP1hcyM/O7w728liVmL6fbhEc+0ySwn9VpjN1gYRPRZAPNnX6pfK
/dgNc0PLBorV8lBli0utuhTagKL3bZfPL7JT1ldEMii1JIWRKMATdO4VkRYPrDg5NN4srPzRO6cH
gmeOqwqaKUd4+ne9VBtNj3sr2UubL6wviBL4JReDPuZZPwvErJkUDHQsi++MnjNrxVV8tPZ6T+t4
iaDIJusjWuC+waY9grx9XNp5uQeoKEgfdHeyDHGJQ/DAWKsXUDiYF8QJwJtljyu5RuFeTqmrtNRB
+Ezi2H+HNfB7Q5YD/OQ4eJBimK7W9pQHqQKAG9yw7xHAcCivF7bXU80ccUkbkhT+o1ipsWuoHYHz
EglWevzGhurcHazJL6/wQFyo1nuESx1I63KXrn6B8anUh8RMi2EoJnCQIPOTz90/XNGWs4AS715Z
PEnN2n0xgG0Hp8vT9+4KtaUnILh8UqirfIgBa6cKFn4uPVdx5I/OQtKLR1lvgj/Yrm0Cmz8zSKf0
97vVRE3HDX5Gi4ssl8MuukbsJXUAc04rPdkKfa1IqOzZtgcYmRO3FDxdow7jiffke8KvGQzscxVi
O10uQTj375oraIg5T6gl4PtVF7i90PG5gSFn6+Chc1HT9R3GVkGSSmy4My3bcwrxQIZu+Tnlkmn0
R9vfVQo/QB/te8DuJ7tmsjFAS8FpGEcLAwjWpl2fS7Mnvl7gNvVLJT85KXtinZc7lzD4jh4ci9Gl
HObqdO/byyAESkBKWborfvh6A2OKCOH+Yef6fIpUCowkTqGkkLSqWBCauo7MVkjis/ngiOQt+ppm
6JAaOc+g6hIxxvy2wNrZihpdy90DrRZShMPeQxu3cKECJm8GTK95KA/bb0rVTKqC89nTmCDW5N4R
LKSBFYnA7Uu67rn0tllVEivUVX2H460yw6t91uTH/DSnhHP/33u2zaVH2aLM3DkALYU/odSe/yYz
/FpBq5LxqXqZFAAEbWYpKdkNnNnaceStzRl7/bKV+5iWbngxvVMamLvoaP2qOtK+6cARSpCBVXC2
KAFlB+NYhOG7vMyDHeSc+aDFvUUA2S8u9QGgIDxHpVD5MP2XQU/i74OvKru5I0Qhdq3AFlG1TLTi
QV4s104yRTCWfJks7kGGTLqmRU6cfUL6Nk3wVLY644BmLsHin5WfM/sRjRtmAMjLDT4imu2tdWJZ
40Fk419Iww8+GyB+wkIAfY4RIvjGzKIJA5fr4Sw+mUzWHnwXI/zDlNJYndlijrw1rwTnSepf/qMb
x5XFXXn2t5fqp+NVL6TukFJHm/Qt+41Xg7i3cWiTjpJdMkRu4Qcp7E4rmwiA7g1EI2xOqt7KhBmo
h4bRNL8SV9pAx5nPUAr9Zrr9tqGR6axdzZS3lyhVdudCp0//UiLm7bLDBlb2zx4DaGvqy/9+RjGd
7vg9CvhX9cHwP61p2a01cGAPHYIFau/7hLUFKcL7pL7UeXgZBvH9dhG/QfVZm4xlQWBONFCSHhCP
8MOe4aUvKTZ/mAcNLqo8OgJtuDTbPovSxNw2NORnZdSLQaCrhcXVuWZVVjS68H/KKQCBd7z0lTP8
/l6vTJHQ7rJa+qPzuGwM8pjyfh6qqaLFmVA/2jqaKM4UiYEJw/1UBY3wAPxJZOYTPUOjMu0bK7Ru
DKlG3fbp9E6KC1BSY0Dj1IFVZOLCTK/fpiUGAqc1HEMgghpiArD7xxwTIimzE1RiOs0u/MxXaxnn
GUI9m7Nt3R0Y1//W7rY1LB7JBri85wSpEdAAS4mPc/lEwHz/zFgkivjKY8rYgfLzHC/VLwXctsFn
Ohl0HcEctckRM2HCAHxDAhRbiVjxzRd4DuxCjK8lnoHVKRv7dsMmsdT998TPED82vcSIO3fc82R8
tLE+jToMCpF7gLYcbWT4sOXFEZ3hfO2tyi0rpms5WPhM0M0bvi6TbWLy0pvvNgnANqL1EtDiWHHl
wk/0VUQk7n9NFbc6rkhZyjF2V9ZANTBInMh9LN3CWFezdnzpmZke6Ihai0ZreZSj3qqp81SWfAUq
P3DFqo9XzBum4DaoKzpJNw+fntQu2ewwgoB9FYMgPT7AVtfG4OWdlPY2xHTkFADF9TpeKQnhvwwV
XDgciBdiJAvjBeT1zonk6gRH/94wPVKpq4af/Et8/sMXPPPUFNBRqJFv7afopJWg7+C2+PCBoBjW
JnSz0thbDM5RmOfD17K7rxWcaQipYZ8TtAuV1fNi9BdvNfU00g0u0c4FmbpZrPxkgfAkyS6qTvNK
HZ0VjC4hI3/pATsRwZF+BCtgvBxWa6+h+mTRygVwrZ6RCt96M036w8F/62OHUl+ruc8ClIPbwJ53
k9rGvUnDF+pZo60DWBiEUVkirwGGNAyEYT8vR94PC3dqgj8aTPIRgkLvUfh0iImbr35YNMQAzVW1
2nBw3bjLZdPhsMYnN0X5aUHtAJJvCgulq5DSN0q3CB4p1qb7Eum89yynu9rg7sqAIPxGp9+v7XbZ
TI0lJ/4fnBcB57GUjW7RBb7aSkDYY3DJAyfERlRSyOvUHiC3YGCbYc29ihtNiaTAPVJ5pdAH3a4I
Zc2YFZWAZDGx6UdIM6p6Q9O5M2GIxoioc1/N6HWWIgNCuVgvAs0A5rhSjzZ/lQ724IxmZX/lEUyS
lspGhpLIxwecx2H0rcTg0i6eBPEkNFwvzc6luVlCBH/HRzlBh+L3vMLIJaqt9EZpWnnpcXnZ5BsY
5WO2SeuyndXrhQ9BWegWGCBrExCbuB7oJ0Q24ku2GlUL2nxsPmoG+pI1C591WJSXeKGm8tMjpPOT
H/yEsD1cnNSUzzF+yi0AcYDMnPzsK1MwOI5/CqEvYH+TAciCtCPkty+7N1PTMuoB1eSBTqUok7eZ
4DmQC5BjZW1p6fqhRXZX1r9mQ+YGM4iv00WRF93XWIMXcYSFyqAQVXuioAzzDJC64pnGC4a9wXAE
ZmT81aXoJRTwvTQ9ixwyG4pvm6OWpD7/xcUQrpl2j9TlwxP22/UcFFgFvzMvhUX4JoF4IptJGKLH
uy2wahPtJgB+9KxWsfYZ4PDBXDEl2V9gf2PZ+es/vGMiJ6rXfrVatBlCvU/YL2TGAyfFX4Pc6lkH
eVRMu5xz8k04O/xKET0hP1QbDR/REx/GyeKCGGM6tF6slrNujgYLItfbmQ8e9pmtyzLIKNXtWJKI
jWmF2N3UgC/E0QSU1Doxy68mEs/5W1RSztOYsnkM4a4kOyrirAxekA9/Knp+qC9I4CjkC4PU83+v
bwC3xEdaHnH3Gj5agKiHbaPfeFOnnQgcZF92O6yZeMCANQLJjFbCIbUcKLfP4beKmREAokOkiDJH
F92aU7Rq1eJupyxVk2f1aVKSma2cNaYAA1RsUcK5lduTMpWV8GjTS8W9Ec1BJ/ej6EEks6rdBhsT
oJFzH2teOT7YnuZdlPBFyf0Sr2IB/UihWQDCRWEHuasfdWmOhNqvB93Dq5hFi/EMyuPxKc3pRCAF
mpZP0BNjwm4AnAJTw3FlXCIcPAZnNSpOX4KTIYufPK4wCzFJzwBStSPhxObg1br5MIYyfzgDEJIe
dt/2ova5Gfe9iXgEQjMvIQmlQ6iFaGtG3SpvKFQS2qWZm6nU648TJFopbf9C6FtoO0hUZdXOff4I
PJ/NjGzKg7HlaKSr/F0rgtGTIT+VRZXIG4dbYfz9Cx4JUtGBSMT76/5ECEzt9gMjBCMVQJkpZhdv
fF9L6gXQ5R5LvzZTvDRmsghE0z1fGkaKXHN3vtpZbF+dFJNlakYtuPvwMpQrP+wijvDY23RDE+8g
xnDVz2hVsgUnU/iY3XoXooyi0Dvu23FEu+Al2b2r9h9X49of3D3ayZqa2RJsVIdc8sLUBJrjTvW0
hGQuC8fSZsbzqmmSRkiUBZN0WAFTlhxmm+m/f05ZGZ5JdJO3hqMyHZIMkD5Ubb6qS7xPG+uTC4Ql
n+5pdBQDEZMYgdVzpgTeCUuU8TXjriF9PiKtzTMoyAj5g1uubjh06WbiGICppFfmIsYlxywHT+We
D+4NM530RMnKvzg1vqP2WSu3l9f/eIvMGiZdwN0cvzDl9kcod5Gx4wpNJXvRxmrCCEUf9QJecdJ9
YRjHLzaY4+eRWn0h0/ckZJm0focnC+suJpRmi1qoH7LspWADJefYCP8DJ+lwmOZmG//wB45WFIN5
Tpc5vEWD4g/KW97J9WpzIE4/ztZR5btaGlxF4qYjsmkyC5d9ZRyyRKAho/Mqr7h++qonmMc6edEy
iFJ7p7BWhiIvYgfYhxjstimjI8Y06bViXZR7LOyQEDOzSebGbgxudIIg9dRt8cgzEJtcaR2y/Wvf
eN4b9Pzlr8+tO5n5+WHcQAO1k7YJnhwFs8v+9bLULIRA+jGx/JSELN3qb+7bMOrjnWMovf7pU1U7
pb9m2fuKZPferuP/jhgCLIlq/ZHQHvpQL5ryPhJdbH+AN7oRatLmln4wdg3nOBoWjdgQQA14K1pm
w9xxg1PS8e9IW6pDGxv3A3NVzcbqhIay6pj+cKTJM11K0jZCYssdSsYFiOaRX3tutzVC4s+LWfNK
GnCAUIWIZmlDYmPu92MiZegg7uQhuGDJD2WhUj3/S7SUUAXN+rOwHrhMZ6v1pIC6W6o9bk3hefdO
ef2yT+WWSGcddkmK0eZ4CL6a0W51klEnPaBDt8ZxgvyQ5Ua5LmuTNE8cvqEiE047kIj7ofhNDJL9
AO5/mZR6193AE8sJDRZ225j3WNm6eRvpVthD4XnTM7zfsUjtCysYzx6v4/PCmn7FybTsXgTDm4Md
e5O8qbNK+ETlp5mlA7ce5r+d+cDTPlOyw5H0e82eq0BJo1TnlKGRUeOi3q85+rpqKcDT7imwbe88
cgnMSeDo+sXGs2o12b/3L9GMGnLn2qnG+mlB+peR5sbMunER6JXJye8IJZv1tCmf5yYsgbpoOOFC
ifbOmMKDFKQxy2gKS8/Ci+NjbPYxiM0L6jCeFigGSutLAWkHq7DMbCxYHDNcmw/BQNzGW9vKRr3U
fLsF2qXc0YjMj/+H+IV0JIeEpPzvq8QdCRvFTMXdZXN3MpXpiSixZqD+COTChJPHdXiZewSern1/
eA4RhdY8urojZsDlzrC1DcK2g2lksec70nsd+D+VUPnCWAnU+/MbyzLkqIsHy/Q/WSlsF75hqykr
dznv1bCDKRLnwDMHfLI4EwFJCWHKsBww+HV4hM9xwt8Rb4nl1cLW8g7pYyV/qEoCWO/XtS98cIRa
jv2iyBjCxI0ObznfWv+uakfyjDrjyj7KP72i1maOMbFtx5E+qfjZsDaiT3AosfwvN2sNILTPe2CW
ajO417IXeLwImJDLUX6wKmh2SIog1GQnwL9WXHSZN98t2KOs06zwEgHEz12KIYXEQZtGijafgsJS
AJnmYfGfk1pVd8Bh4Mc6GNsdGXjVDHZZtVedvPVHybBRIMb1z0fbFllvzsEHWnQQdBYDhUj1lyqi
K1xsugPmrp7VCRoYNKl6pZzqrVRIVS4MrzopKGISNG0VeeR1cex7ZFVsyMiWC7GcgUhYM3mGqcxh
1kPXDa7V1fMnAmquf15vpBCi2Mva1tXzSlbnbwzTo0uBBrxjwkBAd1u8/f5hECegzbhioIXgCIAN
jc37rb0ltgjm7g1CvYUfkjgdL1DF6emnM7j73j59szz16kwmj8fXjHnvSYUZvr6AAJ0/qBhjKsSG
hWD+WLWHt9gqdfz0uXq/k6cHWW9Qw7+WTANkUpxMIHobP/7qfVjNLis7wvMSKJ0FciP4XPL/sa8p
qmk+MvIbZ+dfUry0XwKwbRmLSrwTyqMxWJpRSkBFShNN47xcUqE4uSXq0vWIp5TjnKlfbaRMfQFw
9lE29LlA9gvo1KK3qn3ZqT9IZjoSOJTrF4tq5/CGb3PHTncSbJ9x7zDhSoSgcwVkb0zqI94HZM1M
PD2SJSC0bEPBbIgYYwpzyzAUe7IelMT/DA3jqXQeLcOfFw3y1zKLn77JsF1OMru4o/2h5fXl0xOB
iIFYjkJDnon6c4qhGmMlnbQm2X3P/w+DVr3tu3gRHQMgyDiB9Smxz/X+OAuLI0RP62DL4ZN3d1v4
c9ToLydxyoyHAZ307b1KVe3vGPlzPy2QpfJDz2GMsB+agHtRA8WIWdfcDgcHhwRs/NW3N1XF7gAW
46uxucqvUpFeZYMU/3SWdL1ahhjY88Dutzzyp3hieJqIld6LSPnU6rGYAhSAwyBSnS5/KRCi6A4C
R0CdBM8wYiCeHccMBqz41lby/74DlJkwlLJTptrdOKdczHNmRCwo6JKf5caGh3+g+OsK8apmt4zp
a62tGCFKNN6NE8hfzDOKa31y78OUa6jtsOiJ0jOsv+SDaqdoDgg8Gc7v4jRD81hE01CbZ/QAv8KL
kendGSWRKFcGNhvpNh6U0g4ukHeWzWn8waHrLeMPHhK/R02LQhBk9RyjzNdQ3Y9AHa8Mq+rQixnG
02DQWm/sQzrBuwoMyYeCEnISZjCvNEM11c1X9voY0Lnu/2GnYEsL9VesagBZuF8fp+o3Xqh4ra0e
MHcudXPb6PrM7bCmkEXO0yl7pMEXSYNai47as/90ibud7iwI6cF+N4OZXgTkGkzAqvnhUH1v5UpC
8M0RhhNbyUMgbuZVYU4SVakV6Z6ooY0wnJjamNbYMOgAOhkFRz2fALw4+15lz34NBuTc8TpKnuzc
eSfoPepUUjZKoFcMr2KTZmNQFaTkg6TzbfzzIXk93i5o2GrpTjAlHA0K8/K2Kw/0twu+pVNUTeZ+
KxcfkRVhwfSIqFs405zJvi08KBcmfQR2+g7n5LBxsE6M0HRNtfl7tACSL2fHfvBz/S5I4c2W0ODE
tbQE6HZjShP4MqPrz/Z12nreLczQknyMp4O2b256kJT0Erk5j+3Eq8wCjT5SFiNrtPQj5OspDedX
EQFoy/XWciXau5iiCP/kpw/m8Pv8ge9h3r/hLLUNTFcREuDYWAItTJ/17vxe2B1F9bXXAoB0S6h3
FrPVyn3vc4nGToW2CThsYaRaikx9a/NR/F+2NEOwFEq/R7a1b3rJ+8W4pK5JRYcLBcnAlhX2slSE
vpk4fI1zodvVq0NMaqqiTICukHD/63Feuoa14lJ++COrLkACHJv/uB3oeNsf9ZscDdBS1+/9TTQ1
V1Imu9niCzWgak8eHy4J8uvgDEwfDUIzpZxD/wdsd+knR/86+uOhANe7LCWYGagbnjdo4sN5k0Sf
A0nCypRypL1vuPnXZxnZjyhgvUPvwVRr2ZdZNlz8xCs6IxyE4NOtvEpbDS/2KLja2AHR5yyCzjcz
+6L5CjTqssY4PQ0XUDqw2buHPcBlsWeMIRd9RpY+aQMoLt+YS3p2AJCRSXMUZ8vfjQiZu+dR2msD
6jHatxWVfKoMoE9DWtR7rco3M+uI8U3+TA9kJlCAhDh/xUIURU5jwa+DLjiEgdoz5HOmjyyKQFwP
B7p8br5NXpAgjLnaET4DHR9TCOJ+qicsmlotsZgVhZmqyS8297UbLLYiz/EpnIB6wi/CORs1I2V3
UivW5af/yn4Pi8MyQ49OqHC0Hzk1xlL+ynN8U3tGexauRT/qCmmGXn6xJsKIjXu7hb3WONnT8l6f
bqqSokBW+SFHLzEj/kv9+o6j6V4JybFtYCincnoh5WbjyTmxvs5cRW6x28iydn+WQEjkwHaHIk65
KHPOS9C9kLGkwNLZxfnq68icP/IC9m0TdpEpo63dB9b29u5j8jau24xp+WPpoLEvjyyIhLB9Kix/
aABYGV0zt3iaLdd9hwwDQPmWNoKJMphHoCahq+P0eoAQthPeiUIqZpq4qUqV1Q0o7b2gEcorcY4T
CxNOX9QaMrPxslxB6vhN484Czyd4plwwvquX8mFJSF5sKlhbYLFKo5jmoR4B+90YVMbxLX60f55K
TYYgVjbmrSBdnKpkXRfWqZix2TmnJPLB8N2SZZH24kfuPK9sRfDE4fa3o83BlNx2jJf6d4rpaI4B
+48iE/nHhZ/wCCYuoowkIDpHqkoUxsSWDxOoWJ3qJ2WQ+OU88LVVPHqrkalXULC5Pm6zXPpKt3Kj
Mgp7F8Q5nbx5ycR+dMgXU/aEpr3OVceiGC4LvmXMC/EIdWuiXNSF//i6CfCUTYkgrK5hfV0GeYNC
G6yHfqcsHf5GuMhfQD09MPrc1INOrIuy3dtGGtLHfnI7TrFvtrXLghYcoLL6pzucNslyBvqOysAh
37iXuImR8tQy62DlrhKJdvSl8fleV442H6/r4Fmo/FYswSG6/QOk+IKULec8ACalT0GWFM4mWwDX
ZxmFCCD9vPfI6FmF44sHhMMrcq7DwiFYRf9SCCHU7a3GsWuNRbdnljX3j8P8HCtfuOhb9k+dj1qE
GaP03hl77i/TaZe4AXaqw/CdGTKWjVFKZVOU6YUhfdnM0D1IePKdXDTpQolEddtMnsmVTexZScgJ
yFTMfNbi5Jw8WcOi0X8iR2O8LWDRRDBcZER16CiQin/hr6Twxe3+PUqELw2Gt4q/ABgyZ2g92RGo
MQIy/KB+XbgjnKAa226jTtIcpgcY5B0r94qF1/XUqsyh2s0sVR0yK4iZohQYs4vL7ST3q6KSX53/
3Xgji4BmnRAZDYrFkmOVo0QNhkPUoLP8od1S1m+FR/uY74rg2c2srsCoK5FPHwj9SQJj+i7ipKYZ
ouN3k/vwM48chpu0ZJoOx+LEGUeYiSHF/323W0TtTbaGje/LY5s30lvd3nld7ZK879YnNlU2WEj0
6IdMGAMmFebSXo2WMtPDAdManMBRefGFLZfy8mUFarg82b/+CVqbXIfzheSjCq6v8O0QdP7Lg/Q1
n7q8ixGQBpzD+ndTHaZ62zAm2niOrL1uMn9CQ4SPxc4cBJj95dE0/p0WyGTM5qeqjrXxtREQU9Vf
E71CmHmH67JLz7vbkn+MrxEONua+k6CpsOn8UvIJcjJ361GOQEPGf4MZtg9gmQDLvq+XqHG89bRm
OPEOxn6wfwKIZipiW1Vp3RsvrhxXAdqKcPQ/EVd3LIqcIkWjIR6hYA804klUuM7iRxG7ml0srkaC
C2VoVIuL+RIWUvTefPAZJeRNezIMFxMbnxVGpfB2oPjYrvpMgrNU5f/XC0QbE0m7xl15D3kgFcfk
0/LSERpUnIdzBmDe7NPhYnHlGHeFAQuOthPmGFGxer5P5f7mYW66+1PguM62bzxHHT7DY8fBPFlD
UnH7mQh+NMUxXvZaAia3fsaWk5wbAQkqf+sjepO06urkX+W5VihIdAac7ZvfEGfDlgWQdOWgvqmi
cmdUZ05T3meyIJoiebER5AJzZPAxOOM7frPyeTXuP9sjjNDeksKb9yPlbkKbp49Ta1ML0S9QFhAe
Lrglwd7kxSS5T+MJCIgLJFrDYmKTL+5sa1oiax+1KD3h1bmWji/uyxgVT3eowcWazPgheRdSYG0+
uCgIAGKzGV0JXe8FDJpykhiSQ3KQhexm3P7NqWfx7npFbhHB3ahREwHWuyCxYcVJYA6hiQylvpA3
Cy/nW9PllkdD03XoiAVh5ZZeQkqkhh/ahSGSAOCSkSrVrEs3l1+lRsqR+qns3w/VMsKMSABPKp5H
JIayeLJ6MRdyKCche7p5K3xPkuc7/QtopXJzkJRxX1KMdAvlizfaTYNg/9RJsJRF9Zo8YP6KjXHX
nsJUNDNH5RbV3MM951vkQv6vSWumB6Jwf7SmLI7eC8WZIIBlBI1duJXDegDLRaOGN0qwi3jYStO0
KXfCSqT488xneGchirg2bTf6iDSSe6y9qC+0Aa3rrBVBQ8kgBYJF67P4vH0W9cEVAqyjSJpkandX
5uj+bVDorHmrTibE5GGAePYr1t2AqCH0Yxz8sNMdSjDcizDQlycjt0GlmQjWRimFmNE7GiDDhfkI
WMfoUqLJ/ltmt/fQMKr+B69P3pzjg+sunZRf2RN8Y5C+itdPkKyTNZDYjCDbwOeFzRQyAO/aSz7h
QTeso6JG06ntOebbHPyNzR6QHxUoHhq4IR+elbVVA4+VDms3EtYAWmZX5VxjoeWjaY1xpiHn2PG0
vSuCCfwlNrQOv6InO0bOZ7M3FMIwHCVPIOsul1TI1dRarXM6xj92mrCw8Wt6B6MqUnreCokB/2kT
7rilHsPVOA/j5w/wvvz4/EdKZ+xCT9A27uT/FuaOIO6DNUMb/ALpoKsZaIlIGP1hcvmiNl1S/evb
p4dp1098JqSQLeaX0K7jKjSUUSb57ZnA7qeZwJAcQDL9nGfNmIKYbMJ6WDxIuV9Zcm6PtAsIvZdg
bK0loSDaSxaEEIz6T/Ng8ro/771wkhyimtBoZ46WwkAuKffxp5fItJ1HtrRrWP4GqaMEGYaYnTV3
p7qkYKqSN56Tq9pr6icldcl2rOpLLm82GdAYZux5lfBHMqj8ZHRJZ07HHVzjPQJB1eZD0NVEQQWF
qUdDT0QfCJFEvdxSDT/rLX6XnoXTegz6csf6GbOh5m5jt9b0/OI2aQdvhQypuOntHhYcah37wYbb
ICBsP1cK3AtkdZvPotVlUMfFB98nIYoGpyFheHr2i+HaBLSZ0Z49ZPoWu45cG7xDFaGyWUZJmou4
6ZKAuPslyqHq3xxhU4e0tp2Yq6xkS3vCGODYWLCE62qv9Ri/3y25ZULpkJcAeW2b7IyXoybHDCUO
UuMnTihMFAef+j5IoxWzlsMIXf4ZRnuGI8LF2gxWuV4Vswcb/m40JYa/DPS0ybA7xROPv5FbbxEI
P62oo/FH/JjIO0YsByTB9+uen05529x03ugYZDTHRulPRcT4uuOvHvlj8Z/t2RQaMl/hpnjz8Ir6
pHQYDvrTwV1oEtP4Ay6J2At2lFm/mHNRWKKmKOY2eihOO0T6YiK3yN7ufnVaFHX68stejVa6p2TX
iYXGeQ48iDZetTthZ260TUIqDhtCYWOkNFiAJcv9BJpFnj3iisdnLyOjgO7txpMYtSiry6Bv7j22
ZMY7j4/jkjfg+KQZ8GpEc7Oo6m6Dqe0LkactfXCgStWH+o12iUzwjObKUqEnkNpPA1W+kEkRzRoD
YhV7HZ4pjcS4v/cOr87HeHWssK4xawctVR/2wArbxwU93O5PjMAnKt8CJvFBfCb0hLHF+V878yWu
cRY8RF0Zd829dt++0tO90+BfAHbY7mMs/fzYzQY8JQx4wVplZ+RT2ppU0orL9Lny/m8Xca8vUlFb
EfmHG2xhk74hHsAGqc4IlZHGU4dS33LY46QBjDw5aJwxal5R8nnZZujPDAxML4EEnq6LdbAFvAPN
IWf1V6oTELkeOL50W/+BUpRmFKJuni1pU8J5hZ8vqVUS9E/bde3YqKlHm59ZcXm+njGzWbA8tCxx
fKcHSpyrilv0zIbati8EBCv0DacX/asTjmP7EVtqMX21E7VHuoFXNnEfXGRF2dPWexFgkn0jjBml
DF0j61d+Gi+c9mfd24vb10Dcdm5d0A1EjgVcbQTejnF2d2/t2dnx4G1pnttdyNsqpBCP6hD29TKD
wVehnUj+PeIpiGmPMW1JnzgYetE5KR4yvEje7feF6boQdLV19UDURT0+HkK0/+msQIqOfkdVDa20
rMwTlC2n85Q/nmVRSORRN3nPeZyPVqqp8IgKfit30KfjPlODXvulu67Ycvbl0lY0jFGHyKJUCveP
dHOYAXLtgIRKSSG+21atG4KePGrE+dW4Sxc9MW13XXhpS6MHATsl5deWUHSTZ4W5BNSHU68z7bsv
RHibOO0oiwbHtJN0Qdie6ojFZlFmEvt02jJPEBCLcVX4LzhaSK8v1PQPfU5cyIINOLQ/uWknfBom
Xm8LY5kVZdG9YPdzs7vl9CNzxj8DqKLOuEhmtq1Op+vQz+6vXUZrKWcsGaZ1NQ9q+/eQNj84G2AC
Da1IAZ/R7Q8HCe4FNaIWa5QblwAQGIRT9fypoChhryy/rU/BvGSZmmQJY/xCH25cjqLVJRV+rbQd
HzfWGpmRmSb4l9BulwoufOfsAK7RNk37pjvoVpBfOv37qHoUm7sf5rC4wbCo0pwfhGISHW6kt/Po
WSVuZw49xbrf69UoLaP7o5sDqonF85tJ5ktVWfBmOPstEkekl64d1j2M8vAFpGgkn3dyVC0ZpTUt
LLtr3tpAnENZ+OEVLO+FkgDS2qt4zFBw7+TD51y9sFy/3IQsKSHy9+gmar4zbvWQ93l4p+9PlqXv
tP2ZqOwMGUP8g488XmKw/hMo+UN7b8SvyEKytinXnyKWCycx7zQ3Ar4TbSG17bTPjozI+FvRfOob
+7V5DAZzmnJxNkelpf1D84Wdgia070jXut2Gc5+cIt2haLs2uXCDUqKN2zbHwE6tuo39aus7iHX0
unPACSyxSBca5J4JMqNIvwxU9YSe218j4itIhc0eQg61BOI3bTV88c5sNsWl7Et8tyc8b0U0vybB
Xfb1faBf1w+1ork7Ovy09Rzd1/gf2IZWTd1MjkRgwKhzjLjGiR+Y0fcwVdU2KDtmoFA940FnpojG
A0Pjby+x/K0hqurodrgzz7UAWvYFi4NwoGMdY3jlGQ/NaKks/RcrGA4r503JT6zssEGT6j+Wn/2i
7ZGJB5zdvJsLZpml5V2GCf90bGFlgVC49zsM91s+JUy13eNc9RATawVQGN4FjCRRoiFBZ6vNTOM3
Q0/0og35W/9PSC0FDfdIi2UknvywPVFyKa74YAIZGbNVg+U+UtpQjLYf7ne9Lczoo4pHm6ZisBk/
nlqsjRPwFCtlefP8aQCLVEYhQeqTS3bzWFVnzUSthspReBE7tved577w3Nt7bGmgczseiHRHufPq
N23itthkxZSwkFzOHaW4wzkFi2K1w9Wqsls3SWwxha+3yoW4qmeDunWCAY8txP1rvVM3yaOfPvRk
oDwqr4LECw/xQ77hLQLpSxKhptAw225PqZweA8RuBjBSdNhR5+p3u2tjdlEWlBwGvg9NlAOTcVE6
/JOmv5DKEbDOGpiIUDDtC7vfmPdV5pNEmzlA1MNHgyUwbRTIF1VxxhCarL4ToyPxMM4fSabetXvA
kaqC+td1QcwyVrFOYYFzhMFlEtNiRyBM3lCgPqx5c5X3VtdezkSfsliDzqSMJgffinsQrJEXi6U9
JmJFwvx+ALMDRiFBQU4q8v07qGdYPO/SRNNTVb2EQGe6DOh1AgM8/ACboUFHz1glAgS1Bjrf0aBr
87oNsCOBoI/9dbNzElx4oLEDbezbsHaXvO6qoEu06aUBQbz6Cx/V/Uv2jQ+SjAhnR3ztWL5vIQ+4
Wew4qLh64DZ6uTQXbwHbMkH2ip1OuKAL4oe/VHe418mFHQzb8YsJ6uykQ920NcSAFRU8ATeDzXP9
kpurB/0s88ttmL9miH2pDtY3GoeP19i41iAtwnaZXWW9TdXSbZHoeGssd/TuaC+NX0a8gTUJmAyr
+W7jlSWP7xewfGg6CP7YLALUcc4cQtjnOoJwA2baMNpuIBhuKsBz0/0rDDICI6p3iERElCPboe9b
x6NmMlecm/NBnBlGuOBZP1aUCa0qaiVSoll5Fks5K5HXJHQ36scOnp2mN06PWSyyThB/JpXRHHJ4
rQxlBoJ8olxHVFDJyImCQRfnUY7ohbcgMfwSrlbWjTt4YsSnEYgnHRQkV/vv1s9YObtxQFhuUz6+
p08SAKwr8A4vMbzbgU28Eua7jT/RdBC+8uTK2t0QEsaS+Md4R3qLYCMY1Ikyun2a/cBhRuKy55yx
sWB9x0m5vYqiEQkghLJkk4ZIWrzMxbIqdgILxoRAv/NmVbivYGDlPVGILQrEI/4Xfh5BI1RJ4dM0
G5EiPa8HS5N229L2pgV8e2VlyZjjzgzfGWHhIHrHlQImkxGFyuLjAE/gjFFclOU4MlQ7LdF3KEEU
iL1RjpEGUY5AHoKWG9Xt0pu/tI3kFMPyyH5dbi0DxS2wQy/xJtEE+OymhSLVeKszX9J21jewi49E
NkAiFCgO+491JFB2/w0ab6WAAJZ701qlZjpDcPVxGEiRUlOBxy4Bk1hndEtWlGNBDztFt2BbVzdY
iGKESnGOAnEhRZeyz/5hqRW1TK6IUJ/O2h0pyPGax8/Rw2u7hMj9h491EpA5hNZzVGV95KNLtA/v
4Y96oYCsfaPf8ZFuZnKGj0hTf9WYVv9CXjHriZKAFw6RCzt4XEG2pMalS6SElE/mOaW7gkQ/5N8C
BoIpp678/fWtSm/aq0w9TGVtsuztpnIcLywVdARroYEGnPBZBKVW9TzNQUgNFuEhiEAsI5AlqJw+
dXilFx8ta11qVEweXLRSFjCeOiJyzZLA0P3xmJ7qKjqVWcnuRTEJuR+TJoRkohqq5AhxE8PIvZ6p
l1NvL8zg9UNPIy9k6ctVGyFOTItQ26TxH7eJQDtS7T4w8eU9gIn0Wzw6BlsduaffX+33pwyLB760
7YTyShic3SnhTHgDYSm0OHoI8t2ue+sWVCQAR2ZHSkjuRVI7f2+C7dDATtn6fv9eGx3SYTXmT9K/
cX56xIQSezakD6KiqqLvjq1vbeD1Oz4eJ5+KSRLxSxJHL8Zy2gzhWYv/R462WY8A6LISe+bGHken
Psuj4/F9OHXm71Z4sEp3as0bx/pBc0R8zw8h9BuEuY9GLGA1fOV2xbRi+XXpicJNT0LYVzM6NN4q
hoUbX2ATObZwACR1mXUTnTYbCNzzEHthL7kCedO65vNSDjymuatm0lOQI5WTdEW9xNEbNqHv3CaJ
oMmWZv4ST2nk7MF1F6PYB2EkO/BGMQDCR9uRKeaW3yRaJfpfnTSq1IFMuze2pFzTc4svZQrWnuRA
LpOrDtnrOBJDFJYFWgRCzxiyrzM+2yljmkBUqLEi1+4s6w2mWhC/NltF4B7+oMvYYa+q5Swfrudj
+YIhB/iuJyB9409oIAP1re0f5deyJf1DxpkzHRzs+IHyIKUiJhx8BwTYzE2wg+v0Ctwn6mNuAGAI
5M/IdR+v3HJyK61l1VGDeah4jiGjNa8XsS8tfu6EoZVrYBRUFO68WAWY4F7kKWCR76FKya3T8fy0
O0AmuoBMu5Q45rz0+RLxPohKFyyjIqc1HeMaudRDjrjgt4yB7kRS2cI/AeZg2rXaSbd/zHljK85b
aYt+MNVSZ3ytDAd5BUqWd8UW37S3Dkfg+JZFswn+s5GsTRrrqKHTdO3xHyDHZmNhqHd25eubRg9O
/DJSK2fDUTqNzcso3Rd2/JP1Uu+yKAIFKCPTJeJMggL0g/tUlL7wkKfcoOY5Alv5ksk4u6QpXrEZ
fjJiV8eMiGpkJkQ6ge8B+aHLpaHmHf742m/Dcm8f8GGmmBLVkXKGGAufBTXGHMM7laccKE/zyRnf
Nk2gYrWaUrxrnyLWkyfWZYuAEfS3V03+zCnyN51q6+WmzminSrCbwXcQpgNkUMqZl0agwu+1T/0g
ddELp473gTzh5V3JK8XsCulpNNy23yYfJaY3qsBAXvWzUpiinaVnWUIVcWjWx5tGkuEkYNFg6YcB
2jTKb2ChspElVTgwTDZ8+1hofcdz3XXfaOYn/6Z1qByb19IGqo143QwyRGsi9Iw5Rz7covh0xZdF
HcKC1Iaeq6fPTKbh3xKGQ8338zU9FaQkaQrSVe+iBqRYwlYnXrYlTOjKIiRC0+ge3J+cZF3wDNXG
PMfT7UKLgsusut3tCCa5WFDywKydGljcfNyx7bQT60DzI9chciPwqdFrwkqM2ZyESz3M9He9TTKW
DVhPHHSqj3/95FwoOx/u+SvHs155vz8X/LQ7J9hfbmw0m9ZKoSbOvtplPpgmlhy71wcNUU03qoxq
5n1u7F1KveNz54ZdSCVcQSzyMJGkk6OYLfA7wrt+SSqVrXgCtcmFcykL8g4gUSqJcxLIvorG6Xz+
h9+d2SOuGFsnlVkuLdu6yypiLzr1etNf6ngpwKdSTZyICNwDCnOFnliH7IUrN0JnaPZbe9QDCIpB
pArVjEaVKzEd8UsnpSCqyw+iIqt6CAxa7RjNFXPoZJVAFp+pGTPzxukP34fbAmoWoHdkLL1+RK98
EQw5Qn7RmoS86l3cycAKWBud68WFykHtZxZcGzobUAgY5WAKNAhe78KUorOoKGJGcnzqkWn6V3mq
5lJ8lZfiKiV68p27PaxfC3/joXMP8qkj6dW744+Yh1gMzkSo6JsIBaz8NNkNevoN6Vf9zSDR4VCX
cIggQi6u1ghNoam2NAdcNa22KQ1a22QRAQbAkLbnd5SyLtmOA4NKV7TDw8D3nd7Se8VJhkFgk66R
cYy91V4nNsF5TyRI1ilNCXu+nfl3QqGJK9SPuT7f08+oz9b74Cg2ejlHCoJ+JSbR27y/rX+zzLoM
lEtzrHFtoRch0f+HmYMVtV2gV9J4eJLx3aAD4xMR2ZB4icsFLfhSrLnpUJMmJthtl9gSm0XLxOK5
nxvcLy3cUHA4SSHeDLmmSzFe6ZdMW0ENcXdtKs0yoZtq5XvBwc+lbIQzsH8EbSv5VclGOxp67xk6
8IfCCGMyLU2Wxv3LwT8pt7Tq0gibaGCENQhpVI+2auAnokwuohqHRkPmJbGjvEgTXdvzlsM4QdIG
8EZ+8hz80nW0Cfb2DqfUc2KvsNbFzBeKFvzFQheXtqD/48Egje7Fyn24XsFBZczdRoy0hfvez+eQ
Eii24+gXpKp+cVNOfn32OtBOu1LzfdrDHnGVzqGdtNHtqDQPfHq8ZvlZV/kEnDjB260DrKVykAnC
SxJWU0Dv0uEiKo/bCHdMH9bDkGLAVcdIaS1pPK2btyg2KW2nh1cGZbgOvWYRVPr0idjQht0JZm1t
8QVm2ypZ29oh9VKe8JZgqANsJcU9oqJjLEOKew8qCZR5E7t3b6dZaehjI5ahWc22zVfbjUcA8Xf4
PEVTGFE0c2bEJzZCeDnCAzsg4VD8GODW806seFWoXBBOglMFTSLxj/4XmY7p1HJs2xfvDOwKr9Fu
8QegNYx6wrDH9q/WAvy9wM1C3SbUdLh+FYrFaz3doOPJpJbNzWzBZE86BNdXelCyhvF28AUuEyeL
usDXuviZ3M67mcmjz3Owhou5Vdm2DtZa7eY0YPfykvXf/oqJOEYN8zu5qZljWF3Leyq/ECL9ukjI
YAkiNOI93I3bG5fvcI1kjHfEc64KavD5O5TsTLsjOx3R4teOmr9BjyCf3nRe83GOBnD/0NfZxXDj
gjADONQgV8pbxbwrD3Q+MXcNE6T948tb0KgKsTS914XAk5eNLwNNQZWCV5zExHcI3NwW3dhI78BP
Kr/3mqWepBB2HGenNk5ebY6pbiTnC/Mu8X6HBeKs5R/nLQhRUnS1SWRllB48yBeav7kk+zOmmDFq
9G1wJpaNHhTnSIH4FOxshtqBCmee/klFz4NQUVUbm9uBY/1ntpeJjZicLm3Hid4AkTGZSxYX0HT9
GLzGhhuKAqrcb7ja2baSZyvzar4Jnnfq+pB+YLLoLa9tgQ1ToTPIBjZwRTJjiJTjWM8ftB3XpQj+
gvFobkyg11FcXDk6R585xRm76kMvInrrvz5f2wGTlm1PrBPrVMloucDaZvhG4yPuFuW8L916eDyu
Bin0xjzMHDOlkF1JuBRuMxd4YCJgPJQXa40dNa/uS+B3++l5X+K3VqHhH4DkLlOXX+oj+Mthq5nJ
qWejO4ELfHCK+JN3ZqDf/0BdSvYQb/Wl9AAme/bWoC+22pwl1ITbJdhmOsA0Y7onY5+W2PppPyNy
HWYQk3HZYZODvn5oCN7z9PTwndBi1CcjnzC1wyXbW+ursi24jHqgB7qupfrYhv5K1hHrZusmUV0N
rO/xeB4Cm9lPVD8JXLdasudrR+YvwOd5nFNHj4JibkdyREoEchpy92wKw3erF66igsbScp+ddCU3
MbhDFWAZNpyd7c44D5vZyzYTpGLOyv6EE6CSOgtbqdY02+viXczCC2nSYNUIPhQLhRL8T4v88qwr
VRJ3wS/NQlxIrKOL3SDHeQq7Lp2lK1ycvjuV1vgHzBYhftBdC35N05ojiu84Kr3G5r4DS7qup1au
yH+PBil1OC7lC+WQNiVSGFfeyjYT9eWbuMZdjVF2qRlAS8j+B7SkbGWtnH5eWpq1QcNmTcF9G5xF
0TMOIxRToH1lMreY7ZHA7OTj5WD0uxHXghgvGaYEVHoBobNSqXqQ6tHz9vbIfAmDxZbrI+hAAWDS
MMfVlPZaOHIZ1EqQflbBVMDoLPePyO9FpFasYzk57qyiDy8gqhzImnFuesL8XtLIAQ24CCvrcYwb
ewTyBA5AChAfUey3rtkZAWy070VPz4vgb2TormYUX7dd/Wec2umMrJiZXOIXJvGLsD9ooFAuUDOK
ByyZu4W1dB6XFoNVkUyQJpaNCUrK4pCq/Cd9+mvU7WE7jhE3pygnPV1FPzjOD9RhA/zKzslm/lre
VZmxmOgfQ3shhy6AY7FOicRpGUx9LCfyxD5rHDjp9BFk2VgG8vLu7Et3eIMLW5J0yZs+VwhzJO3X
7mpi262Ujlt/Iu2Sww8oXLejddxk0VJs5ld/LY3/kUjXCPrLl1kOcxnB4NMx5ARawcIstauWkNGb
r41qMTgsYI4hHsaHh3csY/IJHn3LNooYN94xRyhOpTivbZxceUGxynrdN2iSCU2hnZutn9L9iY/d
xjcLwqny0evaAxgKfprl6Nu1zpa2Jkp6b2U8SVvoavvtaooAi9IAPq6vEBMb8ewjr2uCNrGGYnXr
96Dr1n8XK5c/aXa7QRljcHA+fJXLl7MZQ36Axz8r7Y6eq/dP1CE00SDjVmsPLC0hvaGTo5V60zFp
2JGe8Nhp6evQ0xbQpc8uufdSUepJuO7z9J9Hhl/pYFKuhE3RHZ8/w0hlKdhJPl0d9vu5p8SgYLSj
KRzZJK0wWN7OihdcnJiMAGv8HpVHAMW19gDrVKk6BasL0Sa4Bj7yJ+h+NWHGfIIfshZfAwmOSweq
eWQuL0BYnM7U0NAVO1bKUj2FwYPEishHu0z1yR9wSNqklsX1RblnXIjA3fLKo6X34yOgxBY1ZHTD
E+KungUv5TaEyHF7lhP9aMLDWRZD63vP7wlReHT9r6kaaA6LaU2w5MHpEwNhZzM76bR5yZFEHwRg
O4wQJ9xSkWh1cc0Acixfdq/YU1VBbfYanbPDjE5vD8GvzZ3Cgexg6iBFjx81mCuei4WE1oL9uDE7
Ro3FLbjU7OJl9NYOaII8ikw4crKakvcxUEPPSluHi5cUre2fe9H/Nv83lwVWw4XxZtE95ef46Bvo
nqWKYPUIhkkE6r20UIYPFITL5GQt6na+nB41Hz9QuV/u3LoILLaWN5cpJuUJs4vobVhYxA5E6tfB
7y912INsAwweY0ShP9/8fZ0ylKm9V+5EgN3aMMayZMist7otv3vdT0WUAPNCFHwS44MmP2V8Eu5T
4MNBjrn4ojKOFT0vsCdPkB3oE0MLjEiC7OP9XJ9/iqsF1NSjAPz+jUfHO3GcGSTllQokS8mQhTEj
X4bUpR5QNZZUsaYoIfSxj/Ka8MiiSeNQt17+dNYx7Ops5gzWZLYvJQmkzOVuawIygjgDw/FNwDSi
0IGPQ3clpZZGZmbMEkEVgamSPv6VF7KRoaS8ZDYRcmbglItxfr9sTCwhcEmAqnQ4B5PoIMtQ4FZH
OhPKFY6D4lUPI3UVU63NjLNJOZFkQaDUtsFH6oe1tj9mSn5uX4hs8d6Vd8hg3EV/NPXmetLZgAUs
x2ysyZfAWR9gcVt5eEni7GW7emoUiBnzxwF8D/BkgYY5VVPZFo1ihWrhFLS3f6tJD4EgxMdvZKZ0
M81nqy3Cmh8BQJHRd0vbcjgbgQSUQeDuZ/4N3a/P1VcJC/v6qT6uBRjQn7fBXQjRQ8xCj4KrQRM4
d4WlP0InaoTLLxrZKoPcUJ+C6Yo0XD1VcUpzuorfy1LPfUhk/vg5UucBafYmXeWdRJZkqoYNHubO
28hGOtXt6KiATlu55WZ60xcGxgqRxM+UzfiHy47fHDAUzRaWXviY/JG6qxTRj3U/x2qrl/2IYD5j
IkLG2biij3z1u9i55B+YwRrLQkTD5w9ckUpBZ+tHZ7Lu02FL/jWlJz1cVGgBt08UAos31mXP4IOZ
VM34jTm9CNSoIfLtxQWq7klzK2nzRKMX7mpIOslHEjA7gRCO1RsqtWlhWgzsUoUN1AD2Mf0N13ut
r4/GNDHVl74NZ1CvhxAtIbfVsrwd9SCUhmxoYYBkxZ16YzuKTQajLF2O6aUNxQcI2o2qESUJz1KN
EDJdME8zjOod/2BAISxQrDihmICTx+6VzBhkaoIziqbmYgy9Yu9Gg219l46tXJuOW0k+Dv+H9yNE
kgu8qhb65ykRsgaoxHQqzR5sIZ9fXjSt4ZWYEDd7lB34DARTkbG8i1sNdHS1W1yl9ZiCurYLIzRk
WnhL/8ppY+d1YMvFBB3FB9cY+QCzrUAg6luGJgfFpvAT8XwW+sMAhq+z3A2RmA2/dfADf5fOOhfi
DoAfczhdy6IpZwBn4jbZHioQWTa8ZrVdG7oJUNEnFkAufN+SNM8y0sxQP/rkIL29oNl2oFMyXVqm
+M0V9mTGXsSq39qf8fLEbqLNy1Ssrpb5qFo3EwF9mdt1ax48FkbycPEEDMKNrWDiNLOCeqKmJY/d
cpqQ9k317pH1+RA1I9dhs4rzzD5eStvrYf9qamORoVuD2XP1BS5BE0C/atvz0BGHhxT5NEmPQOg0
QphluFUsiw4b3UEoW2y5CcBqrUyWl0cyz39Jr79PGiAYjAgJ1KbsT9Ggf2e6AMcVPuVMdMF36J6d
WJjQiRisJ9BwtU4VwbaFP2owOwnlo0BxqtDThVz/cxuc+G+pgKDqigzDOww4248tOZqkOOkZuiyF
KSuUOfW0or10Bzk6HPZ2li+cWX/toW8Caitn/bTMmXQOej6M8ctzOJ5ngOx419kXz7kv8+ZaW+8q
DEnkEmLzcmYA/7JLeoZsJDscwwFI29MtA6cKgfiFX3OjTbmHHGcpxV7ll+nv8OvmCAFol/cSJKBZ
bWeE8tvgErg2+RDAEsM7nPd1uiT/RJ0y1k0WGmz4IMy1xsULN8qhPwaNJvi6Z/piMVHEDhJH3ygZ
X6hMItixTg5HHLoccGckHH+Kj7JK9CWWOEv90mzHGL2X7YmGmQTUpqJbzzCqimp+f5J9dLaxrGNZ
hGFhI3l9EIS24y14FNzN/TXxPLoxVECkwQ9q47nF8upBIYoRPlnwqCoL/2ps1cFUTd3B7d02XFga
KIuU1SCXde9UO+9Vi5HI8SPRZYz0vT/Wss+QqAkXCCmge8/n22wbGsRtJjVn2/tjvyxowafPuLuz
ULo4fUPOv6wEq28uSoRZ7aSWEYi23fOw88ZRgRz9qEW80wmvBK4wXQlv9HLCxN5PIntOICS839A2
dCuu9hlQWn6cIhuk30L89ViZLP1pvy3uHMD4Oe5JWCPjemUxGCeVTWQJQBJjr0qLjUxIw+Mqsa2s
xQttQlpfCTAbxp1PD4Oa6X4erXP6EDTRJC9wXpMWg55tNwmfkZViFryqMUJkhHwwQPMZzQr+cxeG
obl1FdnOMKtbSN7/kChbqjhfMGX9ljezXBr2GK/WFoxuVz5eVbKmqMRf2yX1l134wW7piigCVqQn
WY97B+UETOqewlFiW5O1KnduCAuo7IUtDMylCqVEvi4+3OI8ws3KlYdGjttJ0R1cmI39l3Na9C+V
lyWCS8ofdteR1kAovCxLwlj4NPySj8RjHr4yEhg3xmPGVpFXcdPjbopcto76e2ho2t9S6Wg1fOxV
8LCipEBwPoJQ2GiOcnIuxM3harbhzLJYhLJosi7dHdR8iLob5HFI4gll5WGndx+sHFtLZnsWwZhv
iqVwncBdFe7d3mByfQCbKQXo59IE7nAaYtNkST2xlAyv/MRkabYTiPlb5mvOkd5Xo7SZRkow2BpB
w2NCBMJ9O3BKbl8n5T3J6VpGl40+lRibW6TAhalGTKRdbftJS5kU7yzY+Hh5aaAxWZmXJBXuvMFL
jcehzBjc8/TIb2zZPOMY97eyv441oXA+4tJ3Uhx9TUij1lGarIMM7rZUBdNDZM+pBvWUwIUSX7Qc
Ymg0Y7BeNQyOR2MmWatrPqDeIjPuKPRySrdS/H6TjdTi1afkt5GPoCnweS8Jft0NKL0Qii18sp8s
4qfseZkSA1ue11FzQwTz0Ot3f5zivRKW4v9LH/YrESXmji9hupDsD515QDmwHYdRnBklpJc/ULe8
ck2liBopOB+5fZn5acFPyRSm3Mg4m5O0rZTcg0XtaaixIC34s/aGLx6MaUOZj0jMz4A46qp8RI5N
UFcq9TDMZJxaMwp7ELwRfgrSahyNxx0+axPcfpZ2kCxvgmQ54kkkSNAqgDMFH2Ln3jS0wWtQgl51
ZcAx0rG8x9KaMnIiXEWl3eGGfBKYov2+hU6vTUje0Hx1SZtmzUjNBPK/TAqSAGcrkn7o4ZAkSuJj
og981q8yPKFHkZk4zzRKKhO0LiX4QPF4AoMBDqqpKgMoepxbj/tm86pj2EBX8NxnZ7i5tXYcsB43
B5drsgrsDVdtelH0HVQW4I2l2ZqbR1Jedh4nEKgRfqRRad16EaG6/GFKm2zJ0VEb/eU0b9Kk99Gn
uxB4q0lutv1uqx24Qp084nL71N//som1pL4fBYm5pTCL/ayewMsa0g6fe4Z5e6UGO/Y/cR0WLgnW
0LxpYpq6Ft79OXR4G2XTIyKSQT1xJ+bB7TJpv2qj5vNl/EsKgAcHr3f8m1xY+2Aeq8kijWRRFhLq
QU46VockpunknV6/ugNsQJXU6Q0V3uDZgeFcKvNFhOYojeTp5b3e5KCpfixrQ37RLOvLqQ3gz7v+
w2M4UkOWj1UUKbUh32f8NeHWqeModgiqzVnAMTVQpJK87ZI+FT2uIGsbMASkiyxg/eZ8yGlPrqgy
RYMTKo4+KI52wjx48yfJmq+OgtPU+Ssi/GNJkje3NVft+a6GvMLTSuQqAGcQFTxSnr5oLNY3RbDn
/CJRG7v/DgCLrJ95CuSdN4qkCBRha+spxFy8sP+OGzzTkq4iDizA9gflDiIC039Tq1eVaAiQ7UKd
DdS6rH+QmoTpDKdxeXxl/bKJXa0SiqPryQQ6Y3s+tGh6aq8AE4PwMpXjKJqpW6bumSdNl0NNpeRu
cvyTEZAb/2+sURicdp0nHifq4L9rrDT5rwF/thO1Z7GiiMjxEMIpnEbqyRpr/iX598hCKFtH1aF+
t5LlgaiU5YgrOgB3yzKHYdFaIvHe6sqOtLU3GGZbM/Ha/U9Z0pPTD+mYhN834czwnBmLG4nAuWq0
94z0sHNRtDdDY3SBbRDYeOytsqijVlZlDIeS177wQUz0dDq4eKhfVJ+S7wjP2tk1tYkJeW7Fa4c+
Lq0qt0sehWneuJaA8ZH+S5FBkWE36WYESvluApsLEUaEeFybhVj9+sLdj260H6Q+Ac71BvIhnLdZ
o5xVOpMfJLf36emLyXT2vOTtwji1ijiZpjzBkz3xs7r2UkWlMdHrhZqQ7piFPyiMbYLv6daDb3n9
a4/tVZAte3OygMs0tr6EvnrcZdz/KvIxOEdK80La2BoDTCv/4lYQqfE8I2yWwc7jW6QeR0JYmO9J
1MuE1TSo38lu8mEvjN+ICr/pLicfQv/qR2CcYy6sILqrqKADB+r1xLE6mFeJlDs7U1IKnkQ+8uAW
Ezlhsv/1GDz5/jRCwnJeGA5A7vZOpfmGvZr460iVwsRj2sQ+kLjfUkciRHSMRMOkeYwBGq60tMY2
NNQ8NLRlpYpKRRoNYhDTg9GPswAWcX0FyVC5cm2gLN7JaBXnPdwB6VPC9czihCORxC3Cv8toyAz9
E+AdL/NJDucjZYEpiabqrJoAzrWNGxnHDaWpXlNA/un7gCpgHp8x3QU+0Tnztfvdrxrbvz4nfxMm
gpIYaMyr0hjjLT/MRy24cvBY5psGpi7EwAiYlYpPCOYPCD/cNpCATaUQECb9kt4lrAWG1Ky7wS4Z
EaoMjJR9vIExDx+DDPqsmv1ZiJLuEgPhvti54EI3RIqTBWLwPI9lmWgK5XaqLdt9jRUUyac/navX
icUiUFh1YAUWAjzvGM+pLDOhf045GeZPDj8Tg2jShlE9qbSbHuM7kbrXeHnJFE/41ktx5bQmJCNB
U2f0Agv4S6BU31frh3N80AVLI4u+VB6pPVYUJRlYfK6kPVp2Gla5H6cmJT9MXnssxmD383TmDz3m
eQxaXcw3GEQYMjsXjnu5+/tzdBZ4UnUhldxC3HXkKCCdSm2wpkX83hZf0Wx3Cs/7A+yEMVv7Bq6M
8U0EBEJvavApJu/PUwjM8UgBVe52nwXrI6sSQmIpMK2B6LPqQvhyq5CajzTb0DtmZULFkNY29HOe
nkSQUyLwNmJOmOTXtfaKnWk31itIPE2lvMTwGXvoEk2w4DvujW6M8T1PhUSna5aYXVxCJZNjfWKK
OYfgUqXv2UZwJElE02kBLyawUs1s/xxFKCKHHUQf1DqGC1CB+YV9/UcrrrTAiSHHgkxYP7ii7HO1
+Ga980s4s27uGKtZYflzDfnZ+JORKMpWCwS0jR8vooiFFj7nxYSIzeDZ+SB0MRJXS6NV8zkN9nWS
v0Q+7/6m9dabBbXh8ZR2ft7OoW5zImPy2wV5UE0053mcF26pvXd+xGfoyBrkDCtvEdWR29cKMWTu
E2YadDE//GWuWT2cmCDOqTctpVRmpMEOfNr4VdXqzl/yWf5EEk73/8ISM0BUDYUZNTBZuLFoOxsw
nwij/+TgxFAewX0bl6qg6E46RreaDJtaYeCTCRagqnosvtu8BXx7UKHyK7UtmCayHt6wxPUmenyv
U/xJA/KdlhbS9f8mBZ81EdU9cSQt0GGJqPENDbvLO7ut3iETw+09R7/hMa8O0WAjMYLypjQiCrEh
QBMfl/3o262z2td8u6FJ5Q7epUvEBRn8zEV3mzGXrEejZvFrRDlWxkOiiDUF++golpUYOAb9mtzm
mcobqwmHbzcAwtmpEpR+oKZihCf489a48enSlUIeKGvixWQAZ6GsmuNhUXUu8seYD519KymeJtXT
G25PLC/7GVoAAdnYfFJJsyqncWTjhIUbK2eoohvvtLJmAtxX4CuCAKDs8krRR3maPHwwMXOET8uo
ISI73/Quc4gBTJR2Xp7uLkxLE30LPtBVgkwc4leYtyVpPmiexcogaYr5qMt3jPpmy7KTx1/nqfWH
73XCuDoQDLV+Ru3V3NNuUuM1RqtkdA4X1Fuc0OGek+vEssbuZlgYEgkXc1q24ereyUQmXd1LONSg
uEAGX2dUiPWcM12OBpe5yqnWyAFHrWppKNUm5UWOUsNWEIU1MLFZDu32bERmcVX0bHyqokL2XgLI
vpMhrElsc8FeSV3duSWTZLq12okxBH5dJRt2bCXOpdD7Jp17UhMZLN3gkqE7BAWWvZwaRmr4lA8g
4fri8xWlxjek8GPoKOd+KOF4HjJUj0I6GNXFUoEEfzO/umYH+UVKrhCSQhDs/vxG7YupnclHCJBG
dN5qS9gEze8ApKiAC8qQdkmMBsb5QtJQncFjcnOhFtlXnWVyLZhLBdS8cdLCI7S2fwEI2K/YtlXZ
Sqmxxzc1iDKbTHxZw8SbPleHWO5kwu/qKE/AzVSBjdW5c3uQL2RmxopQaXAkHdbE6M+mDQqugLSv
r22xFmBHPLafiKKfSpKXYcj1ylXQCuCt8+UHbL1I0X0+G/f9+M/mW2Xl+vBb3MFUPAIMgpa+VS5D
4kr0SDwaDLTZGH/wZUgU+iF1zYwC4XxtddGYhR8hKbqZ1XlLpOhtPC1FXCDj4bOL6k9R70QPE5Vr
c0j0msh+dzRi/MtKpMitcLCea5vJtKGYDZiYNbMXUmFsF0Aqzz6KlYXBvuQIr69ib3xWCfxiASK5
CEcXsh2nhhFzpULbCDb+S5vAX2PPv4kSTZSapQQD31SZykMhT9xKF0q6wy3Ay4CpYz7/qxZCRefT
0KjRN7ZqtQqSsMFcqcSh2UF/5dnsO04noozitkcb6X+yTI3I3aDmp9r6sOSLLqCvEt45PsoQn/lm
dFCPiEsemmI79SDr+uUR/dNwweMhDfKVBZO8xj0mYNcvRHrE8NrvuxAk3K9TxasWVGtllWESKSi1
Ew3WDFsLhLAsZ4eDJYl8NWL7tY2MsWMYszBM5T+RU/odmyX9W6ds5+EsGhIJ43YI7wyABx0HR0QD
r3TTuQRI/FrHaa6pkdyiF7diSDL8b73Q2on7ipRKYabgO4omxt5ZomAdyQ9/Za9ilcxafR+wR5bD
TFeCpV0nmjg2baqFjjaxEClIqzmXvWdj95frQ1xwDzfB+MzCSbAEeLxFbqycYyOtrYJYtaF5tv7R
uC83gN0nAuVTBJwHuIv4b3vLlZ7bG3MF7XC9UipI0VBKkNUd4swxvT2yLws3SuTKuzEYVjm1QV1c
LyI9o5ZSIloQmKI1VtTMbhhDrMqSH1NP5+Yu7wUSB7bKTU4k2+jRIktJsu8ZzqvV0nJpHf4PT6vS
H/jRyzYfyyczU2Kxb0A29uWOWwIGKGv6woYL8jE1ABw3Ko1Tf64qAcpmmvO1fgj1N9AwaVbx9sHH
fKvWlngNWfwLn7LdYfiy0PGOkroOvBrcijddC5U0bWLh/VCGH64Q4N2t3l2g9/P2UFjq5DxXhXek
N9zd/m9mgsslM0L3n4omqa4tfZuh7/pYcZiwBGPY4trHclWV7CxkT6lCexZ6cBpuMeXjOUBAxA0y
D38BXg/NT7ouF7qMycHkQ+ytsYL2WCxTsuPFkVUddUOyTgayH73hOnxyaPE1y29RKc9C/R0IxBCb
gnwff1bna1nU8+FXYZzQ6nEREEUBjg3bh+WgG1EGWK+63w6un2VzLCS9pZDA/9LtijSfTOOLqx5p
h/m8ZYvsgtHUJEs/NFKGyzWjdeVHbrVbD90kJNn+2jgmevgITjtLeXvGzfOGnj8S+7ZDyGFyaF4h
ZxMRlEga2mg0mR79IxzlkPJw6GHuIIkx9LlTZT/rp/ZTAxhw2QOFIPaKvKlDsv5Mt7V2eCxptiY+
wMJ1J55akykFCpaMRj4Rvt7ehkNbJDNlhDiU6ByGeAve+ev4PMjDVthmQ9F4ad/JolfQO8J0hAli
otJdKGeBoV6CZY0WZuXVpKi+9NcvgHzsRE3SYLQXEd5r1XWIrBnLpMSsbt3tYV4ru9Z9m6nXcUKL
XEYK0K7jZxk98n7nimvx7+Ren5DNNwcKgnb5dhpFSiKxz6le14KIabIFKMJ2lGXgZPbZ4e0uyQKZ
HvWzbYZ270AFXXT2dkdhj+vYq42DvfH99uEoN01eXdNdet3zgtmpEcI6WlKuiKlJvHHDavI4edlg
sFyHJhzSOdt/KYuyr5ScYuVz/BZd+hL/+VNikaiFZIBi+RWl3j9fnjgURvVxjGK+Zv9SXRjsi/nb
zBxO7RAWLMQuuh/mEaLDLIEkJMHl3+UqfKnlmriksjOUreECfXNYly/bnGAVWH3a70r2dDXYlU+C
XzLS2lenxdp8/K92hyG9+qCgJFvzlmjt02uLCKtX+LqTqoCDdJvduydoa2HW6YS2VW8AG3dwl0Mg
Rd9KkUUDfSGbWqq6HC+VokpSbgXN5VBv2zAIbdONOXDBHFcpP/ZlDqWGw/xSOlsqzdDsex5ZVRdr
NRFy2wsFYWvjJfFMTvB6k6Ap9K9otIr1OPhLh5mbMRKdgPDeQ/l9cyF8YNUVPlK3JJSkl8MPx1BY
ZflFjRqdhT2+/4VodyDbdJGaFGH1DbzkhbLUaDPuE32ddJALn7/G2iSO3NZX7GBHIz1tDZn+x9bw
IxJ0oIElbJAQIagZiwV+GztHfoXfdbEt7qa79ojUMYkTU7LRXIjfbryYc5lwr25wc1V/IvEYOlF/
5LfSqvqol8Cih9Etbi080GLRceqDQVEveLI2pbUG9zDaq51BMFZnxFfPi4/yhUMMeLIJ/Q7saV2G
bHc1Fbn6SeAzSAeMxubY5syBG2pWthJ5kxRJw2mvd5PHL7dua6EyE4X7w+q5b5c/SMWp3GuAyAib
u15p7/yp1uO4/PbW4S8JprDtXHysZtXac826wGv+75iCo7xzOtfW92LUbNNiUynEyCE5yJ2KXuX1
0SVVkPF4Wr8uzE+KZMPVlvoncEjoUQ4+gZ/2nnuvvSJw9UD6ZeQZeSkG+UgPumIxYQcZW8VKdyCw
ANabnLJyjlfRUrDNqEmn5EC0DSAAvxtHakmvV7Anj03bilAggVXS9HawvbeJygD0A+t6tTW/2PBt
YdRaXYpLs8ulgHejrMOjA8GsfIFj1sIG3PnnnWj//iMQkh75ubKCr+FjGHmJpO4jtmo0Pg3ViwvJ
cVxSIzUb5BP7AU5NHPLOQixcEa/pS05rjeceXGX+V4kcyxtQA2Rd50usgjU9f8EXcBbDCWstunmV
MTPf1yZCyyhIXDVk56h7sFWuF+HeMTF5lYbaM2NoaiD4ieXbfYe8CSBWbXIAxJN4IGzpm45vmRFP
RxrGrnTZFfcM/EDyDXNfYSde8M3sn20USv5yFI6byFMWeeY26LRPY8+hpFkYrEO3I0/iXtqkFrn8
vbF0ynzUtKQDrBd7Bz/6PlCN6BGf+Q0rdLCiVUsu6VzQXwKLODpAFjwHIXWNQC2HoulGkJloIpPN
HAhEbTP3uwYl47JO1UaOgSJG5uViw7U6NN6CYYTrC2m/+eRhIYjeUJB9yZIyMLiejFwCiiFwDL4+
V9NT5tRWT/7f2hDA5kfNdjWnsGO2LAvH7cjSnjVtLoIJrlH/bZU0S3rkS8dcj7D4lrg8OO51k1d2
EVK3pdRG467EPTfTL6+Fln+R9Z+mIvG2zGglbYHvhMTp053iAF7oJQXMGoKDDCyBJW8qhg6Ut7Zw
KToo6OyHK2qtg1HW1pjWhUv71vEJEIGJHKxT10EDuRPycYIefl1YApl5Uovsd9BvrBHMpH/vF3ir
pIhis655ELZK643czfkv32rTYE7trpPYbRMhivejakUPEKaSWllmEok8cqqcW+ZpO2WTwcxzAlR4
vB8SzpthLL6eQKaGGW1QaUnkhWgJAavqOo1xMLvhJ9LVq4ex/f3QN+0d9Jj3gC8OAEbCvJvaM15H
1/Dr5Aj81LXJHQHH/IRR1c34iB/f2zYzZRTXM2ADirRDzlWerZ8FkW50W5QbYB2wkjbSCUNzWaCg
HxOYU63m2+yst7B05GEk1AFKsdc1n49UtORzUOQTzCYbdpl6Ykk+dIGaCxUhDR4P5Grv40DZIsve
SPHUdKcLYtydv9lpRAZ/koTyMaNnWM0FRx7V+9FtiCJsdkJTCVi3fV0nBKP85PBXjyo8YNQEFU5+
dNKWHA/T1z2V//JcDWqHHKQLBFbdgojhadFqIyy9HqMkmwhYsmS13i088olKIGP6f4Ybim6g6/l6
JXVAywni1DJv0uXzJh7Go4aa0tcGjgnOcxMvhI4Pr0rEUmwZ5dWqfByudxeWAUKga0u7Av97j3Rp
5v6+T8296Pf1qmx6qqprsITsWkHX+S5VvmgUaayWuqj1A7PYe79zD7LoOEmdr4S2adJoyAahm9Mj
rPu0e886AtV3XtpSRG5RdvqcxhH5w4K6tz0UbUCr1PYFgFos7OxIiAWn8yVDqrfxaj/UTXdxCFQ8
nK79wDC1ibovYwKQG3CyCLnymQLWFHnvB5xIa2VMV0FNHV2ssYwhMnaIluskAG28D5AtTPTIgdrQ
HaXMUsGWEBGNDhRAjnH1ucLzGnwM4HNTEQot8LmU9nooMP+6f3emIanrur+4giUFxgzOTSJddhcJ
7cdkrYrDW78iQBu9p29eZdHzmKB3IC7su+dEtyvgMbrflx2RHwJe3R9ohdNjzMJvipcx+G4mzFC/
RTG0mJLmwvCSp6Gt75cOZ0aPB8C07J50S21cZRJpfr7sorJmkF1OPqWKBV9NtRzr/0ynESsL6+bl
H3tQLpOrWYnOV+hGxZd1nnj0aelUFT2D6NNVjMSraQs5iITNCa9auC6LeO7pmy3Ckz+Du2whyPZL
aG839F3ZWmKETWsO8Wh/9Im+RhlLOAFXrzAAd71zLQui92vGd454XId7d/V2qYywBwxbsBQ9/2Ip
Q/NIYu5LVugZZVrCOrQ/Lq/xRldmcHv2ZJU+kyyVF5NHju13iGDusb7hlNBF27Ey6WBcHOpycSbI
/AuwhVQu+IWa2OGtRPUiQX45fXHD9iA41oBI7bzTCNIHnnlqPxOcsCFHbvlUClHFvj+YuwdZ7DYg
rwSXVtPJDFlMEfA/hpmBwER8ZAY/8/wjF2SJZFiCLdOgHYFiC5rxLf4tq5M0aw6DHq41zMOWREGB
UgOHbQ5dgD5RVzAWygOTMfQtEz/jdql7v48E5B9bKLyaqwBt0nT7jWTgczWp8D8XkpMa5S4JhTmJ
2T8+mUnxGbVl7Y958wEfKHERLZ9tKtG5HI4w7ylzr340qFpWSn8yjY6IEqo+6kp9Zvoui5bdmtBu
ROMx6XN9Spj74VA12NZChfwUcKrQWrvqNJgIEGAZpW+sO+DNl1q9wlA9cEt6CIZJlYkWGboHPs9O
YkKAfH6/SzeZwQ38rxbqWm8MCz7MTh4JLc+vJukuARRZgFBJWNkWyctSVkqhTEzjGwvP34kSNcNI
upxdtrsseC/5HnIUK69pXnbZ+ga2950AVYu/3xiZYlzLkz96NxWRDWabEwiRYJDAWt2xGNpwrOGa
+cFNxADcdon4RWL9/DvbCsI/ltxM6jxnI+gcqhhRSeDLPjjiNMjN1dDmsvUecOI/CPK/Cm5OuWUv
fFwsjZv9bx0zq8c1wuUp2X/zpd1w4dOx6Fbwo/BP19DpUctGcxEzV5+W3wrkjpl4L/m5cG54Mr9Q
qKEHwdBk/CPNYGvvp2WWr1JL5zbNjQtO6oKjaGwZtcLHFmxvNP3/k2YiX+7zC9q3pJlY5MuulKqE
iU1Utis66MIBikeMrCcDRorvBoPXo7jT1hREQkEpH39RG0GI1+Mlomk5Vloh/SMiccnlUQ6rXFwl
HOSyRGNe7miaS+eyaPv3RP2yc/Xhpax5FN/Yfwp2/fX55wtaYzAFVXQgoh/BkUGDFT5yAOcrXl9t
m+d0YZ/w86PNTuTQPl3dW1Dnm+p/+haNOFCw8AVROfv5D7QLl+9h7OVphWMbD15rjAC5OqZpIgEq
PcDOHo7NLl0a72rPrcQP8C9zPeXWlc5TqwwFDQSyNXU1PzVzKR+3CKmhGFlC28qrQdXZ8RZwkgbR
fGFVpFxgPzNhxJ8aEdrwJEH37CFHya38AYGcP3ZuZO0YZrjt04z92TMB23AXwdA+HnZNeCX4wLWp
hgrNVuqGh73mpm76jgjbM5iFPEaYmOuY7/KitrEIh18gi/LEFDKpee8rxZiG1U9ngCaDkxuj4sj7
YKj76Zga/I/k/f37Op2lGKlyGm1zf8ypVhaqZlp41hEm/AaepzAZrKRwP/1PB011ilUq0opKin1N
UeWn6REhTtMWuPm5bq6w42yN6IQvw+lB2kYKOX9Q1qeI+Hdh0mIzy4Z0bvqj2fB+oaRt93RKW5/b
zLL6JyT5G3j7bKb96tciWk1ZTKutDQHfloaJD3PIPSTwJr4ijmHyp/DOnstGDZeKF3c6Og6KZV68
sgN87Snnvf/+kSofUVO5NWiI3Iyo8M2R6ZrUzRsmih7hwgM8Z+wMbUoeLXxzgVPvGbNh6YIdKkp+
kZN26xHbpd+3dxm1oa+aPySK5J6RY1Wuy1mZ9wqQmueIQs9x3veaD+c9IYCSUC9ix3PkZjxASFND
/+LQyIPIxeJk9/s4Nfx5c5ESE5q2JKAiOqjZkYwLsVTrKSu99YQoS6gEDkNB19EoaThe3xG2ewir
moqgH3E0bAyLgKS+86I2Ut/xmQWsCQ+fElGhhHiWEmZL72/RtTSvjI9TmlkyeeCcWSlPTY8bWCcv
UEL9DSBTMXx9RxAgZM1MjL8fblZT6URIZNoLcbA9jLteWRMIrGAmrMW+mpHumnS7bVee5LnIRfqB
tFiAzp1zEQd5SnctIbH73yUr9YHaxfaWPPGhMY3UrkJeB+L0xlsi4h663GW2FA6+/acWN1+IR+L7
5PQZfPMhI8qZqnJlvTiaDkV+f9FnFep2KbZay+j0fKtmtNV1Gt4T3/TYU5qX91XzmOHBiqWukegh
JbC2KX11dqdpvRz17/XvIUeqAyEwHEgMhAP5m4EdWd8HxJd+w/C6x+e7GXHQNA0J6uIfLmw/+yGQ
DBiTS6LKgKi4kofnACripIHzVCvUybC/bX4U1FRXlOzDtmp9kxP8VR1jQm/VGMqQC23pToIhcYf9
RWShhX5GK1e2pA4iJ22/onLKsbf/q+pGpVqP2tZSifTc5SMW+HDZm3x8jY9jfypg6PSfdk7WTTT9
zTDCucdVTTZjsVejQ3DEqoWZb86sLZ6+S0LnJlRxyC1s3BHcHWz6wnFIashlmtWIE/l6/CkUtxgk
OTVTym14+UCEUCyIdWhEIHXtLUf6AWdMe07bPjrK4SVOfuJUHkcZlLvmyiFwFakijWNx1d7ZVmT2
NOGicdZgumVhh2aWKKMT4hl4WS9yhhsB1IKbwzvpOFgI8BJfVW5Nx9uE4F3WKiy7Ruu8TXC2ShtY
7nFtjmxqEO3YPKz88H8miyEmxRJtM4pYZPJQ7Q9YAdj+Uafj/y6WmKc3z7HTGzmjYGzjZ+o4ijMp
jTnLcC0F8uRkW1IUTp5WfjJ6nFPV+6Phg+Ggr9mvWK5MxPYsm5Euyu8DChQpW+KyNa3Dc1bFMEHn
Y43VKuoX8+gtB7nDN2D0L/bA6Vt/8aXCdpWpLeU+QDabWCznjULkNQE/538iXDRHmLm58ONrxuA+
nFJIQXLPJIH1da6SVBtS23rgA9VGVm4c0V7NAsGuPGP21IIhz+BOB45bfViftv1dubh9L6T6uYS2
/FwnC9ex5Aq8R/Q5CVM9S1mYN6GWbh6HWdv8YmhXgDpEUikrMiLuS9r7oesWsGkqoAY/5l9ypd1A
6nP5uACE1Nn3nX+1gTwenur5lfxwUmI6n3sNpi4xGeh1LceDpXZL+6jrIUEos1STHmIOfl1IJSfe
wMoGNH8Ii2xju/h+YIsLGgmAymcG78RMjyXZowjR2uiTvN0wFLk+dQDI9+C+ZsuETUMZEUw7ocAI
DPrQrGXxINoFjsgf0CfWsaazmagappgPTTcTf2lgolUzg3fgoMMTehgXmScw8/L2CZERJn6qpvE4
PKWC+DHUWWetvljF6kjXwNbU6AyBJ7zeIWxPiQY4V6N/naRnmiNPp623oWT05DUE1UVCDV5v6c6s
EQ+jwitX5z5+OhRIDYyq24hxpDZ9lhJ+nDs0O9/HGDYwsxnCyMPvuQW+Qdb3TpnrWU+dLjd0OwAu
4AmNamHdixbZ1i0i2adjlgQddBfL9aadYdX14aRi9ffQK/43GGV0TokqW7pHeWkFHrAuiKTa3lle
C2cQPxN5+ftcR1gAANfMLAHfCs3ISluCTh3m0en9RT/A6+9CRs2S8Q7uPyH8Cg9cP2MDSFdNc96e
euiC8FJ/Ca0lCeZwylXqFjTfIS1OpgylBUD/YeCGQATQm0HdilqqpqtyVBsgJbR9tTsPpCSJI6yU
+M2SM+JZ+KnY6U3z2N1YhHmyXc85dOsiIUcyjV6O4cr22HGvjHKohSDHoCTPC+rIoO2WA5P0JF6q
WJv/PpK5b5XXfTVqo8Kf5iF3WeeoEu99BzEcDvEsZl6v4PRxtitBlowyMai3ARyAWxs5Hjo+jend
Y+qw1SzXui44bdgqO5Yaldtk7P2QCxOhRNeah9SQ3KLAiN26DKtDJrT4YnCyEacwhX2ENAC7fcUw
koIMGDG1hr9VU0gNfmRB6wVUIOIMKQRId2QIiPRJyJci9MILCdk37832qjRq6g20cD47NOX7ytuA
6+xHzdw3bn0RAXzXWgEjBtejfuynHmmsf/oYmQUFL5FDkMkhWC/7pOMANiyjjCs85cR6ftdEmNj6
0+DEABS7aPYlV8dF1doAXIelpwrJEJfEcdd1Koc/rYSZarZzo1f6WDmLbgIUerReM85Pkf2T+ir5
f1dmckFUO8Vve7e7RJz1IxtpxWUDXbVnzTQk9YJSOo5sxMYwwaHCv3jDu+UHrElxkqb4czKMviKV
PrbInH/rWbY2+iu4oHOuHFTt28cYy60B1R6jAwlwkwpdK3/nkQdo+ssZzQvrfC4BEvjkOa9tn5JJ
Fhq/p4sWYtggGmQY9vqeQ2T72qmtYaMyDvC5Mft9H7GXInLU36yT7/GnXwR5qGSZNpQ0s3LsBfFZ
izABm/OeSvU0nZvsJtxYTyZhGAtCMPcOfrB8He0nUzKDYcpa0lOvp4jwNtCeoRSKxVXJ7n8/TQuH
zMHsjf+aiBwaMW42y/Ugc0qa+ss/c1UTNi7xdUQC3ty5rQTukAYEnl0Y8AniRjql9kB5uaBKQyQ7
xG+Ptbg/V9e++7TQ81bL4fYKZEq7wpEPBR+4EmCDkE7ZALCleCQea270gDshNzcIuTOhC3Jjs/yB
5saXhAdYC/G2O0y2uCUiLsqdALtFw7lSXBWlJZbfgBW7TKkzFv2dvAOq7LM9rCurDw9a20+okzpr
NOL2S51FNFtoBH1uRfzra/MH1o8nlnRwhQB9a0nFOFJCF89+MTQDkZGbmy++9Ct1uHQNEHGiRV3n
yAigOJNP8RAqfa8XiC+BNrDIBDVMFonxIARxCVKoL9xoVyzdNS+yuKZu53guy+ayO+bvSwwPfs+a
mbLhTgNwDj78k8+cXLERF2V8ENbHj42kvFUmpEMUIh68D+fxq1T+gBgwcGOPIXJWDgednt7oUWlW
UqBwYOOat/v8niVg8HmD/OnfKGB4lF7WBjj51t+e0hupSZRKvD6B/WK1eg5tjzNZ0tmrEnUNEpZk
urSm0CuzyAcn6EtPRub6Oagb5TgWXrepH2ovEES9uyQlDMRGONQ/mPPF/5T2LXNSfmna0N4uFVMr
716ouu1XFrC/b1OZabSM8w2H3FHhsK8iSZpMMZ8uzbN2Biq3cLY+Guyh6y1YtJIScyJvk+iKh8/N
+i/E6AhHZARxpuus3GGtbFpZIqrYsczpPi8iMtCxhIeHb0UNSgaLtbTA2V71z40N3x1sGXbFbQNM
p0lkDw92xGelGv9IJ8Mv4A+brL3iH+mnCxVzcMLGya3A6FGNvF5BYKdsNUthQ75BgJlShaGB2thW
uQaotfPHhGeA+z2nbpuGFoyWD1rqkVx2A8C7cRGqLs2BCrmN1MzBdRgLwYHx6jjhUCaqebAMtOa+
XlGenl7lqqYBeX5DjTAlpKRdJFxo0hR2RM5W1VITcELG7A0T89lEqbUuJAON00XDYHsVLKEu4oq5
Xz+ipgeMoeQyX1X6aPqCGyEvU41umlJLWQgzC5Xzu7rhYLH7IG0o6TFgasmHak4RNVSCOeAVetB4
zItII5dyBWIH3LYfd8cjeBwEKnIgeD/rvoBWukv+q3mpHn80OgbWlbGr45keu9KEweIThWb53i87
5E9wsVWox87qqEmAWg7E49Eji0kXYwZQchGmAeGKLIOIQU0CHWyGhVyQ4pWvNVRPDHD2GpYZBeAU
gbeVOQE/uNeCUTltJBbWv4hXcVbOt39u2Aylqom1HvnNRMh0kTSenUrcpSuYA3Ol4LwQ/9RR/zam
hwJy3JhIYZFPkqB15e/Trh+H7K85jP7Qi9ZJ/I2CYy85S0pnQmY9XQlHI3h6jXT+5Phi1Q523juV
RrCOXtpQpn5fFhenhey0+2SbFrvOzXI70jFpdoSP46DsUCqcPMOOxx8DD5JAxk/Zrd0pZ71k2qaG
uw9D+OVs43QRS0fADjqpujrEdm63k8IPqKg+K0sLVXsZpVYzXMrCmuo4c0tb0m1TRSp7+7sr2w1a
kN/SUqjV6YdqB8+v7t6hLRnJPn0Ze8NhY5aTx9eNL7Qk+aWjjIJXIxLLcCTCS/vwJutRl/8/t4Px
ICPfIEWk0Tbw1V59ED/tMGSIsD6vgr6D03At4ktUxMnjJA3KduQkzTvW3uVh7L/2Z9sPkaWUml7a
a3z1qDneSp/hsnQXuaEPOthiGS0FDwKqm6a7op9Os+Z6wMN27kkVzOufL8SjA3slP6CFooFcBiSw
VbxnFs8DOIQk3soFHSbfDz/lCDrpe+eh8f0OajAFQz2TYRvfLVTUMDDBN5/uR6CXCxgkacN9TYwR
gsHDRpx2WBBoa86FabycO/2OmK6NJCsOS1t5Ds2qTy0UXo1oIzt154X2CT2ALnz4z9eZsjzrbGjg
b1dGJ/ebl20R+0tntKQ6b1E3Z32ZpY5jtgXr+AQbVvt+fxXeG7Mn8NnjMHghpJPw82hPlVpmxclX
1Ha5cbcEWPgkSwKRNClK60TNDkflLsbp1QHMseVrFB2o8Jlt+Y9koxWr1ImCNDsVsl4bw6GzmJxu
5Bf/KGYgeGg61LWlRkyfE34qwNm0jWYOC/JeedXX24niGh/QUIdGH9ZjvkuyHAal0f/7a7pKTDjt
JhJa/yRegUKB8xuq5c4TnJGQRSCOyvTxKqLU0JNtrrEGs+Svm/r96mCr9cCGbFTFPD/gTdzE1yKt
/QvAxJzfiiCASrrocBbsixD7+o6r3bNJKzdwC97gDOUpi9yA7vB9Eu8htOx96/kqENKfKAPOEfgq
369RYqfEVGZMsqetZIiYaxMJPYDjg/F0Ku72UQ+vStGJ6354QSsWt8HI3GqSODVPYwO2k5MUZDEf
5bg6wUVriRmOoEVdhb9OYD5X+cdcNiPR3DQvfuk9Ue4ALtzUwp1ZWFSscBLVDVPh4AAI2M9LhIKm
iKsCDf1yNrkSjAtwaIsdmvwz4N2FriTIl1rE0KE60FOETgOCzlekuHqaizrUAKLmBF89MB3IEmLF
rFu8amZOXpK1lQTsXuWsKqQIQsx1qRpl5wqQsxeo2WnufK+eLWeroxD4POAlnTdsNqkl0ccJ3wS7
rBxF51UqViOh1lr15ssFJZ3c7YArSmz4rnDTNtPZoG9FkfEJnU2ovXZNxcbvVXRRiG64hg89Hmc3
VsJ2s2nzP/nHeaGeXFhWNAbpbkykSkxw4F178MlBMtBNGojK/KpBug1OBxg2heJ+NnTpciyv2jt1
ujETfNb5muoDy9NZyyWS8RcJd4/BVKTvdvfDqEutv2mL482+08eMPbJJW00H2Ckwnk2bMHAn1r0b
f261vB2mDnPMzRHEq0sBE4V/zFTmMFYDUk/KyssKH7Rt5YqJtKFLzAAQGXnxA1SHLVI/mntJKWgM
6nPY5iDrkUpElpHO5GYHs1TWxuabcElQv301atGXmY4sHSDQ0gWpPW5YGQR/iakKWl38cGTQOHQF
dcXe9PVCC35TC0MicyRRt6fcDQ4LkQueOIvPRWp2z48LbzXuY/7Gk6l60zPEY64FQhUac21/rpDD
gLOyNKfiNC9PuK826JmpmBewvz3/svLbnt4hmYCJ0GqexsuIG7g87FY0GrtWLq+sN2RDeSdL7eBJ
u1JAcnLUuxJYUJK4xNYDMzWR6ljR3gN6Ke1UK6EkLN4VpbCTzVPtVRACLrgnoOaramHDr4KO09Y4
ON0b2CRQNVwX//yVY3skg7c2XkhwqS7NhOytADb18upWJYRuZSkMW+ozhafGhSuONzZhgNOlLWmb
mtgrjj3tb7+VInAzBrFX+Fb8Ur0DvYSMN39e5XXOXuEqP2gujhxdpYf+Pcq4uiITvz0XRUlu2RGS
FoICEP8lxJxS4DAX8qQDwgWAYUI2E1QuCI3aFtiiEtjudePFWLYpCGEmA5sMamaGmw3w2yW+5R2P
xk4ooEm0BOIyePLb6XWk8/Fpj5+aDITFECsXvOVbnEQX1WGNY/awC0ZCDpDPsUvtgeWLY/GSG4mQ
tDWyWFNgUV5pK8zGFYDR8Iqik2LS+Uerg3WDgCLbLO0UE+cey/dAtzcf/ICdpoxBrUN67Y8PZzVI
Uo74j/miC8G8nXtT0weCrOW3voFI/WS4sA4AWl0Ay3d1XqTM37pVCVEgU9eQG9+qWiEMrdZmThJ3
KURjFfKq2WzDFTm6LAxPa/P7QcNey+Levj4e3NJV4SzOmPouFuJrihN99j7+MIjctkZ7mzykuiG5
4K3GhR9xFYtFUTY4pP307u1xFY6nWzmifOrdsJOWQIvYGJAnMC5Sj4wYB6mkte1U/1vr6s54oezV
2xqLngamJ5Qi3yACh9PIPcjS2S/0OcI+21qB+j2fNJ6Ni3cZyWX0fDjdJkWlbXaNfXPXn++g9KAp
oNo7/i942xMYvCJGIFq9FQQuw8xRgeV/JuBn2Bka8LcWzthsdIHItyAqy8iz4lbgvmdpHGyESje4
8bFeeto3+5JNw90iPzysguGxWjicBkU4TvALLDV19jvrXDZRaMz8xH6NhOq7tGmvBPflvI9noFF3
afbHD8vB0sr0Ja2jZLhBQsIai20XdjHcdpu2LYhYzMU7YKSONkirMVpAR3zdEIpSvboOcHBA1W/R
Y3rsHaAdSVOptPgJ3hNDDHW657NCWsnooCd9xuUVijbREdOmr3MyjEHNh6EtcB1RnRYfUyf+eVcG
ytIjs/Uj8PoLnr9iLjfrXWCRIJrTCGVue19RRVQz/jwdvewDAe04vFGGZYAliDKzxnPb5xkYWC2x
bZxtEvEZ87mkCYa4W8iUfCNFRnOPx+pE2+K44+q5AjetORaAcpnRVztDwrwB5C3IJSzqLR0Uo1xZ
Hagpy66kDgKxASIEoiT35+Po2aNWhtIRVNKZQ8Um9XZ/7jTj25m4Fvd/BA0PtniVnXAihNvs99Gi
f9euJY63TBzKTiLO2EkjW9qKKWH8qodJF2tZ2hzUE0zcNcfUPWcVpFJASUwtFmue1bAwtLjXj7zw
ZFxAPDb3je9tUw7+7ApBuhNU98pLxrn0OsS6/V+J8byzASF812sLjHVvTwiFWoSs2hsQ+TjZS+Xm
cYNBVeJZ9mXxxEXLPBXC00mSI++ZON6FazaNppp/9Xpk1krNl/jc7yYBkkgq2oObMvJ09y9lwaMw
8eCfg0fw4dWwJ3PO8algb8BmLQOrioTBWP6oF6en9/g8nubyUvXyVo61UShAVubUgLzEh/Cej9GX
sUujEjZ7oAscCaVE+mG47Y7mkLtspjgSz4c/O2m207xobWJ/DbRLIwW7GQLFFqngW+OVj+r3ezKr
x30o7XQMAJnCtaAmXs1I4pwMEfSCa7j2QkBBI0op7x2NBD0aCIWJs0ZtawaYfa7tsUSqJptR8UcN
Mqi8tJJPOmqQruOnzoIsnLdjqkvcd9BuSrMvyxLr+OFlsX94QWHCR6LAILjHa492l3XCYiY66EzV
JwAIjP+sGJLxh83rLGJA4IMNG974ADW/wqOHXip/DRrHpJAM2ERZY9KFTA/AfyGv9Y2gAnd1a7xQ
VeTcdhey+d0WH98DeXFCDWbK4vSN8ysOKy4f+wBoohaWXZU9ZzPzvVqj1GxtOKfSq9ATt1erq2L6
TJvdqnF+gHaoptOeHbirRMOFFig1G5WsjmOqr7dawKqcOVP58kJWT3qmpT42+Kh/h4n693EiJvq5
A2Suar6pL1CKLYQwPsNI92ed83VE/7x47KxJdafBB4VCjG6An5pDywD/LKwllGLCn6dQLRRGVwog
sdLQ8jpvwS/Mq+IbegHRO4rMzMLlCGil3e1yTsyAeikehnCKxSroqw5cRUa4qoK0hjoy8LzkZllr
gQonpoAl+ADmp4nYrVV6m6QsMorrNk3f48+eHssuNoascRi5Kq2QqiSHyUQV6ECO/WsfdG3F8b71
0KS8bd4BitgRU1b+yGHIMDpUxtg8lNlT4gsCso1XrZAQkKZWilj21irjIyCVUrbr0ZjtDk9NZexC
XVIkFZmMXmPvtMIFusnEHN8kIeeZXSk2RBuZOm94U5rkBN8xSQqq1WFZUWyCdSdMl8k3FsInTxa5
rljXtU2+Kxv2fHsLG4fXWNj5HFY9iVy1wZhXdOr2hpEtHRAU9tuC3zMaTRdE+2MTWn5TkbyRmUka
pcNa6zWjKWL5OGGQvm2OeKeYw1uYWscIQeBZnCZOwhkyGTaNHP/DgssNC/OqZKrLFTPxNVPYRIq7
13YvMTVqhkNgkgT/WLbebUheyTwH0lyTqdt4Y6w4dSbh948u4W3q9EHwI0aFOqYgN1a3/ulS0GrN
Lja4v3PJ+adG4789nVRM1VRUsMRmXKNDxUAjcdaVcxDA9taNVtQTxk5xQCWVQfQonag3BGcbLJnQ
Y1IVSEUJJ7BqAS2EeOEtNShWWCD9cLi05Wq8sDvnjKiUL6N4WXtK/KI3i/NQPCrt1yVliA0YLgV9
uvQ6uP1uKe3Ms44++RoswbfkoMKvamimJKFZrxlpO69ZQRTIc4pJ8IjIirtQiTnnhz9rMwLJBB88
ZTxtkAlm+9PV763LOPVK/jlNweFWEv8+nQow+NeyfrB6Tyg0iIGX/pdmu1HZmfh0ToggWeelR6X0
nsCN9Jewm99WLnWmbIEGSdbEJdJDQoKYiWhzkSI6T4tqMEB7PeoTBIF9DYc910kNR8xmJHO1Ubxa
+BOjJEsmlelXbYwJ72qGRQgMAG/BqeZc/pa3z04PfK419I9H641tcGb/K17Wnh+BGZ56OwkKEC6E
AxM3ZO7LiOz3wev3mpA6X9EWPqk+SmJd+UXUoK+x0H54FZHv0QAZoO3QZM9JvXiFH4w4zJh1F0AK
GeF/O3ItETLOuBYQZBkGAXwInRb5hqA3hVRzLVKelXRn5yRUMTj+6d1rHnM/L16XKdicgEsMsZWJ
CsbnZ7HWDjzwVuDhBw39RXh+rf+0fK4OO5Hfkvy5ywqn07Y24TRmgfb+2CKeRVL6++AF//sCP7Mq
bf4okB6BUZog13cCObThr85Q6meWqzgwnRvXrYnjTQ3U3FE9nq4NytGH6xukXUCiws5x+5nlqGrz
wulUPr+FuQTcdVPW9GrQ6oxTm0fx34x5/CQheVlsUSKLNf2Ccx6bU6HUPwnPqGeOU7eBCRXUUPQF
wnHgtP/Ral7U47gI/PW2qoCnli3+lDLuLolsjDpThpeJ9wprjuJmTqsbDUFYq6DYOA6Lzb5ctLJn
t6tx0Wn+7s5J6eREilDa39uBYCDB23ZQgvh3sq6wM4tB5y1J+tvg0TFhXyNB9tWGFUX0+0JNQd/W
y9YdKZc7tbYqlHc3dU7YB+tD3Ui1q5g+V2jN+jvQUFdXMkltx3hIb5i8WYziYGcsf0zKs2HIGWu2
EyLCpxRWfqXeLZnKhbzxL0fxsXkU2Z4zXaHsPQ9FV0F3bP8XQXQTqg3GUh1/tENB62z4aP8CUxkw
zV0PrN4zusQIqjuzvUPm34TQDRUfW7bfMleOCmqhedQ1muzNtJc/CuZ3okqzL4kT/boUtkQGk9vo
5hCCBPQkWz6ONDl0yrknJerEAl4McTkTB5hEynFiUGAZIo/iYI0aGMX5AZXUuhcqc9ncJm80Gs8g
3KUlTV6Evn5JTPtxq1Wher9V7ODKCDEbmKOEkEuMTyocasVQWTlR3HRF7LStwlq/i8iqROdimRp2
cqemYHFeErvEbs3Xtcs6vVmPPf8xatYv/knG3vAKzxqhOaEeYaCQdYI3ZfohwWghGLqqRhzbIaDK
ZGzPS51aFmpUfEnLjo0iZzN2wPco24yPo7/6Vx7TVsSioeXMVcXKebw2kW2QliBwaNKD7+x0Cw0I
Pde2h6mADyjsfO8ngluVDW0v/GBvHCm0E7T4XSJjeGrk8kyy6kmhc91q5+v6vcFzkgmkuiORNWex
P9yhJ66IYAR/tqxA98BNMmC/9lFSmsYUWfS9WbtbAWBybL3ZjGbKvRQpqqkWiRTYtLeKWx1yjYYP
ZY/Vxqe8sRNeoknv0fR8DhBT6Ps+m1x4F3EnOxe73JIutFyr9c5YQN05DXBFYn/0Stb6TvWjlA5a
O8PZYawB5zujlpe/XFAFaoEkz3mq9MYCF5dD1Y4FdfsgO/d66zHtPMhi1ytknsLMdNTwpYbavMH/
/SFx4nYRxGg294597BOjPVwGj5KLJtHKreW/qjarIIo2ZpifAOzs//miYKsyYjgPDR7VbNCvSaZl
GjWRDH7Dna3nLllxnYAZ5TJPiR6N/z0SRSYM2gu1nYYhGwaTkQs3cStGIzVqbtT9pdq5dyw3WPF9
VUrVlVWEqkW2e1C1jQ9sT3LmjOYzh5ETpc+epfqo3/6yiock23xulCAbtwYR9zi6j0jlksVF3Kit
Lya8W8fQlaqCkvrm7fcC2NWMZvgmmYR/i892+Uc+fx+cxF3HJj1MknQ/QkY6zDXQqIrartkpg02D
hSsAZpLHLwTNowCtXIJrRqnW3iBsJPvXoq3zkRsLlzC/BI1PrtShDYGU1GMfRtpx66wbN3ZgWi9x
oRZv3NMHkYVhITHBdLFkJIb7UAqIIlPlWT6gMBujudpuNj0k1UNilmKeCmYQ3iHphvpeaGkVQy1H
y+Yjb7LGMzvVqgjHzcxg0JKO94iPRhUqvZTCwQB92VybXcty82IZoO3CWaN/0bPnfqghJGgIfaFf
ngFVzPWyiO9Rv4Yq8D8YXO6J4JAle8Suy/E6nXAHrOwFkobBbYNHCJdxdlBHSYiJVRRYw7N2H/AW
Il92keGyqxQw+U2rdMjfhY7+vvxI2MF6eVUX0CvEW6U/j74pzQ4srfOCXL0zeCSafG2YJ7x0wMEp
tujcZEdy9G65JcRYwJTwQDkemOO3T8cpasnJfnkunTVIIyjGzJhZZ/jHklEHCFjwD3DGc+cTXtVr
o2TBWCyxHO6hRxnWlFjXdl7zF8ZabjCmz7L/z+a8GKSCwJrFmaw2RIV3EaiiLBbsKMO/ZFhpz7cG
EKTY93QnixsXAh6DgHpARJ/wp5MIAkv7YjKz/dgFUKXgBvjPZ42Mu1iEh2xmG5HGqbe0ttY2jyS/
tuzuXKgOHPwm4/ARFAvgMaLefpofJdGUjO+E5uvAt2cY5mt/WegQC3nzBaFOs7Xzpi+ts2kZdHlz
1vAERFm/SDuj9ziZcrmIZVvC6NPusc7onkGUduY3p7Oq2ocAUG9N4OBDAJtzNE9k3l8UxRljIIDQ
JatcD0wd9p/3c7yNhctI2+zZv/h5WyXQs8PCz3ka7o8FAFTqD6VjVsNQhPHb0T+2sVFG6YcCRTPM
hmsBPoOPG2NVmNPzxrWSVfYHvp/zMZyklhcuBrjYJgiYa6Q7cLVVkIndauFT84fAM1/4TELzcJvh
8fZEsA2ESz3KbLAbKCKJ6ACrdXYai0IpiIdrScco/lKo9bec1NjAO/4VOBl7V3Y7foSkrqaCHHGA
2S2PBjVZfSQpwJ3bgMmK/RIB1IrLfr1ODqtnC3IWPxW9vI3Zd0X3kkCuwQsuqQR/KIEuNzB4/Gcm
G29G52XRSDNlDHmTyGkjBN/Df2EX5cf30/IS/fmwWBwu44bJEn6m7gIPkylSi5+35GKNm5O0RCb+
VofjUcPHyIk8QgbpT+CzrklgVzcz9/2UewEUB6ECJG4KFOLVSlvP9PcPmR03FrRlaiBxyQKh6pLi
H8vxOiju7rPHcRBe42zA2yOxsNImBDJz4ESNh6ofluOcEpfXldzBvcIdIqQgxGOxXi89n5wdXiZ3
Kwg8z04BtbFLr35+BC3TP70r+SVmSdsYQLgWfWKj7GOGcIRJagQVM4qYYg5HL15NtX2/0WmVGSFJ
b71BmfCJREONPqUvPnBzVz9poaBboNTBLE7O5y9SdSOpFzv5TxU3aMuAEg84olI/v23W7ARs934l
pbNHGQdrkDTYj4OwYiRFuCOFmjSn30gIGI4f0l0CtqrXW3fcKZd3BhzIfgsRiL46PstL8WFDnlE9
xrAuXmzNqX/haD30Ou4bcEKrkYXf42uEuUHR485/wDh9Nbq7UJ7vPZMM1db+tnmeOJ3tQbA1ZP/M
t3GD+6eXr+a1C+uVgrYJylqnf+ffZwQD2oahkuIDXbc5P4sHDitnd9OYEzNYPqSIv8ikkRjURy1T
ILY1TvfSCNUiQ+pDel8r9pSS7X3oH747BnJGPmh8dhalQhMgKDyeL6txRA3uWvEQzdj+tonITAWK
7heE4Ux14f2olcEYeLYX0Hds32NY7cUjRUd84mZTCTxjdlPO10Pt0IozncO8jqssJo0rZeWCFJJR
3csDloAYSdm/qoTa0+eV1FwtGb60GQIaFsvKFBKyyXXhlGjVRj4GYTnLsRk2f2FV78c2sZaoiT+d
LWIqTsjfW0Q8iiIJtI1Tv7T0Ayyh33fDqz0Ov9KI5YwPILrxvs88oPEd2TCA3COah++NyCfTDNXA
pn73Zx1Ul3BCS7vVtklgzm1jC2o5o2pGx5GAU0yD63WUV9rvptaKTvTFrAEaIpuv7WdmCen7gZrN
kaAdEH5VU2hNdlvh3uaXsj460tRFMeciSD322F2FBykLlICkzp4xr5Tr67NKBr2gwIwdUG9MBqhb
nLwfZBMe3yPkJkaTGFCWhAuXhyXNVgh04hXLXzehmSLiJdX3RChd2vq4v7ZkaWbQ0iyo8UBIkFaQ
wl2IRz5VkAgSfsOgtB41N0tqSmDj/NAmoJ495vW4d75ccN7ECKxn57EYhtqwJdMan5S2troi0SPe
D2Rchbor4xZ66Dpah8Y5r3vhBBdVWphYlINyOiPA15m94RAqovw5T6NFyOPLjF6aYWtaVCYSucxt
1HBSMjgL1wmDRXqvB0a0IlGh8lYZ/32VNwJEAOQ3WNYf91TaTePYCrfZgKcw//ZkySwDWa2nKlJx
L8+j+CCpKPn+eSkEdeffhjWJbUaaqZhn/ttWvjE5Yz7TvK0/Odd4fvYQzMiv5zBp32FCd632T8Zf
lUigiMLduVBGPP6pawfsYvStg2nT5xfRUoTUrAp7LqH2C+AYplOpxQrXNE5ffAfvQZ2ldi5UXjWx
pl17AMaJCxSkaWJ9q6YjBZsp/o9qO62HjPqJmAe5vtQwliHkCaRwXTX1w5q6YQkKgZTUegABT1Hx
XjuKK6Ch+iXGTnkByosr/VVIy5A7y5YuFRh7jnkciuy8ISKAOrFlli+dtAs9Gb24tbBvXtOiRJ65
HUZPXYMioOII+3TmHJz7zUqPaDg7RZBYXpcmn+7JKtKdBfC8g0F3HOFd3qnEIC8pr/5Nf7qx4wXa
r8+eNRzUdoYabJOCnqDoRBEu7hgbzDT//PeCeL4kP7TrgoWrKjvNSlu3AlIcsM24jWFu4SPEIJNk
W8E0ed/YV1Lpy4Hk3f+VlTjdOaDi4/EUt4UyzICcJ0Hk2zImMMAaGqZLrzghXz8rTx8v4F9XvurC
PYZzQ0OEO+OzfoFHZ+JeIIADiA9gKBnDVWBxmvS3eysVo+dayX9gGes42WiQD9DwTErIjPWLH8aY
WYE2MYar678o5Q97hT3ZLdEVEqy5cOAHV3fdwOdmqVvUb7BbYRmV0HW3grw8gxZeW+zQE2SAswBO
zqETAY7jTEBbC5UoGzfnE+zi1QOHHm9PHCT2gUB0l+LCcvwr7P5UjPXuTQIsVhgKe6QTuR7+eQ4L
e8vkWAoQJm77zRO3rxDXYHu/tLRx34I6bpziN/Pr4+IPGqfiei30JUvZHPs/mlsgu4L0cc61Zmfk
55UjphGwmtK2lpPAmEboWLGqB4ZcdVIO2hUxWt1YKfve81vE5TD5CEVMftK/rTn+8dopd6DPALTt
fhc1mvw4pr5sEc1EtN4C4A0CnShBlAAstOMxRomgeHsVYyFs3Z/ojJE0BL3KRMvh1aP07Voy4ph5
zwv00U3yLCPb/4i7UKWvfirMNEO/ILlGsCk3clCrXlg7XRAEA9ggv0BoHLLN8EmnOy2MIPWRRyHl
ZScFLQmD85eosYYGi4rKiIIi/oC4sDlbfol9JqCr9Fby4V9LR/mcddC0i+Pl8P+66ILfIZx8JBgp
4E1eNs/LheohsXIhRUzdIQk873FA78aRyKEqISg1gty4JMOIo4DNGIcQK3avAchR6KEu47ePmZmY
32a5C/ICviMBJeJddhJkyNwDqRKx5SUTCLj5dcNRCnaCtRYUv5ZhOUDeCXuZi/oQAybvXZ5twqvw
X2vjBVsH8IBVAuHoNWwiPzKJmo90PfBVr24l78SBIMYicrAAwaKMLLozefmTWGJsnIcGzBlJun80
tmqiImzSgIqO4AG4uG03xK/9TG0yYznPeJD8wg58U2UJTi+qCajqAOun7hJMhcF2mfL/qV7wFoq9
Kh2kVVGyb6zsqpzaCYria6yPTjW+u42WI+PQsZ6eYX/3IiB7or2dwX94I6k1TUXjPdhVFS5XcOnW
P0mbD+bwIepFXpmUVnB93crHJGdgDlJXNNm82u1YvzuvpzwjRw9osC61It+r/EFyxw/TaKWdaf6q
XfanXNYtYd4wNMVtBybX+ZqCGd+nMFBbhQi+w/6unM/3G1hN8oYRCy1pN0Mbizj7f/9rzk2avK6g
AeLhu8d2l0pIkN0+oegyjHuacEgcnscn7hOQCv+HszrLmG3fFWyxNIj6iW2/JAb50/lj130oLusH
LR9sx+4SUkpl13ckqtBSjrBHazlAVTEz58Lfdkzkdg+gtLleWP8+QjmnUTmEmEmrp0Vp2IhEvE2L
BHPnNd26+HHyvoRnWHU3jA3lgRxI/hoXV9096T493pkZ6InFaHG48nYTHocKlGsrs1ouX81TzpS2
5VWxYLaxVAoOwCqFBIo6cMIPIHWWjmL1jD1pwwr1niLrK89J3eADlVAv1F0vTmZPyic1px/IsMBJ
NHDqb/SeK96m3gZLO1/PD09ZG/9C0i4LOi2GYpcrWnoh6P90oKXjgymawdXGetPjGsXzuxdL4fss
7hgpPD0JBTq6gFuuX1739Fu5aZZFgRmHQXnUBNTt0FB+4mKvdFdWDIZ/S6EbkCKv05JrbJ091+9T
TxuOb4mLP6IdSYLhQAE2OKO+5ccMNf+swTaoTML7G60b4pKDIrG3PICHhcxJtW/p7T85ysOSceS9
uGNvgzdvCoB5WRP7TxdB40FzlLNdO4XvHoipbXIYPm7hcJlCOz+F4tnE+zPeh7EAtA5ossRbVmCZ
xjEnzpSuslx1iSQQkvhiya1fvg6odauebryI0ke/cOTpjZx4CY7TlaCYt7Ob5n5n6cFA1i1O189Y
KDsDsTgnz9baFcCBLtERc5wCZ+HBYYrYdqYWl1G0uSjhnqJTTQRTojz49t2a9XKvy9LrjM6gJ/FV
usa8rein0Flk2ZUvdxqNA8X1lEGafzi/5Vz6wbBZYZuLdRoY3eop1zKe+Rz+9KRPJFk//ZaViZxa
RLj3gSl31M3ye/U+zXiofU39zFSyn3SWq1ioulCXtQkx3SOurZ6bYNGv5HCcfrGjV2Pgie/4qCGV
ARk754ycMZAGEalCjgFaMOP3AB3VtMhaBqB1+AzpkzrK5sfQwuyIlHBRyEXESa3r75T3Fa6DudeW
yq1Cw5iciEz7VjgWvy8mRljT53GHbMG0HA2AnZlx6CMqZYPPAk/qtBkZWvHPxz6Kw96rylU58SG4
eYLMA4dFZFuQcBkbvYn2BhPAsqVXpswBP4fa94KJpFTVKamEEtgxa/vMd2lEA3kizOKiX/97he/E
fcB9v2M4AFaPPh71PJQhpHIHtsULYTTgSxHt3+GWEHo+Qj0L1eWzMd2mWEl66QfKNIxx18Uo7h/7
Ze7pEnntcJj8HdYEkqOAm8cT8zAiuBj4GXof4k+8HmPFIBX4JOW3UAPdNlc8uzxH8KReTT4P3YYh
xWSDCgAWgi9iB8vRBj6D47VOFQL5LmltMq/qMv+o/5o2/vQEi00Uv4WXHV48C1EnCJ9xbGY705f/
+IXMPvSaIyUWrm0rHw9dLvPmn12WDa7u8KMOIJwmVOs0VhkUW9TzG9xTNMBooVsv+CcYD6qkoAEv
ismy3bRYNqeDv5XQw0sW8d8fGFLN8lplvRih2BkacI2r8ebWs2n2H6+8H+/Mu1oBgleO3WriTqym
oIKxTZKwH1yHFxgmqQ8nqKlG80WJ+OWhhgT0oBJVaxeEHmBmqlvDfx1qzQt9JhbyexaTb7Gb3UfX
IGOfKlbrnf7lrxGs8hfdG9ZIt6GeQqVr+rS3nu21dCCct/ibN5GTZ4AKV8uJrBUXZSrm9GU4fWew
CelRsfN6Dwjh5vL7SdeMCeZRQ0ZnUZZn4/BSQeNtxkTjX+6dF4h4PhzBGOmEsH8/MJCB881IT2Fd
R2OgDVrZ20nnHsAyxgW0x6vnnWt3JhGfoIDyjcqgia0Ww7sA1Q7xO7F6jqsAafaDP1J0hunXehti
cthIUv2hwCQbaBy6SsNwAPjcq6VD2pRxcv2PgV+MOlpvS8lpFN8OcYp8IgBE4y+hWd38P4iHLKQO
kf4KyTWjRvx1cR+I3R9L993Gz2MoQKm7+ddJRhvy2rRH300eyi+QTu4ffpBphMlRF5Z/LXoX1DJE
dqxeCYFNlFGYZatfXrLATb6RmWTZDF4YZBgP0nLfDGL++8bbMH7g6+JMyADLFYhWEfqcJmBjpJjF
zEet02B6MSoTONzHwZvRz1MZLCbn/1SBxToVQ407EPEs1nSeN4SNn6BOzFrKhvCogT2HFTxxd2b4
ox7WuP/03/gh4DSxizuCaOkl6W3NIIP3obrxhqXUU3LO61upXj8Gn7too1kkTOm+WDuv37plm9jR
vfqO3Is1I7VlCUiz1Acv0HzNiStgI8iQ7rfcWAxr3wdierpD6xSHPc7JgUVHdFO7jliCQDExCMxA
GWVUPo7Pd8jGhbl2uRdqf5XO7wxOJ9LI+NaJcAhoYW6j8/e+jcPVoH50y1FFsUjPzKrzdF9hbcjF
Ud+W2STmhoD8f3iYVV08Sav8Zgs69JNygk1EnJ9cZFSD46DBVCxCk4a3/7rpfpsxgMgLNQxkVPLU
4HyocKL+0/vGdYNHnoYlR9erOOYpiYaY+rTL+g/ObTwxaRkLy3wvl6Brrq2oXtS9AkQV0JxVqE5T
SkYyQQRfg3stMtCFsDkQJ5DSv9R7d2JSe5qWzpnfYBiSk6vsMr2cUN5wVqJO6GwQ1iz1micuwGBQ
G50oHUGHat7ejhYvrVgMXGhPnk6cWD9AhjNpC5xMvaMbUKFxLiX7yNPBluuTqV5wJWZ2lPlQcwPO
C8enWh1xMQVRprE54So7qaF8aXfWzbG1q65aNDZwPt5sjLOOo4r4Hzu4nDZEYNcq5F5p/D2I/dEe
HiNA9KiQXXhUa0K9cqoQiN2Z6rjZ+d8yu1cNieWXaxDBWyfPKgCI0bjhjaqb1CpnqyAwmCu8KH7Z
tgsmmN0EydEkVgnLWqXoZyUByPC7w2B6YsqD5fYnUiYsyvpzneDvvNUcn5B7+2DCeOeyVsLOI5ql
vGahOj9fYlW+p/QBH1s/36TexVLcEX8OhFVxn9XK8UlbC2tU4ovmec+mP0TVy66a5Ubgemlsu/95
uwMjTZdVf0Ewhdgp5NLqOuUVCKKjqCpjNuVWQfzUT2AN2r5tSZFsUVRnTWdgF+OJDc9K+N2/83Eb
qLCBA5WLxC+isPVyJhb8HrtIgtpakDUzYe8zcBEmRILGOQq1x3y4qAjf5Quyot44R29+5+UvvNq1
WbX4NAIxvGvyNXdKa4wbN3tIfsRlir5k3Kkoougbsy6wbGzPUD4l7vC4T9JLl7jv7ILOyZyqE8Wb
ewbTzmzsnU64iHI2dGovlRZYxU+hDWha4lmoFYuyQljdz88csmjfHxgutQzT+VK9dPF5V8pzQq/g
w7osbo83V0FtG8/cYJQ+mrU4+bJFQniIEZts49ggJxKCc0QIvKZHGl+EsIjUgYMkzzJTt1CbwU31
ubYlWkE1JqTvxTbhhF5EWT4XA2K24SpgGB6us8c9Eg72+cEgemyanP2cWCt9h1EGcJYR0EW8PCYh
K6CLqYbtThCLUvxr0AeU17b7qPMOgMioyjwcLi3LttsV0TP47JSO0OxjIP9C27BhT6DRBDvhqCKt
6aVYEjtgMdst0q8Z6Nl4OCGsctW6B16lRM4YY6a3WVr9zjvXhZyzj350Omp8rYjA7n2ontrHRnRU
FoT1Z9rynwGJBPJKkRTOsFfDOi/DGGpsoc6O6/kwPhfPKy9FJIDcHxjJjlHxckQpxG9WVDoXj7ZZ
2zjpHvJ/c1gwMSALJIHLt2DDMFlz7qntXio51GtVwwGJLpqInYexVE2ZDL4ecLMepHS7cCvZhkwT
T2dgBkdTbuEtDgKovgnG+dZbrwnrZfUshGARGJ7JJnFBvScU5KBPLyvx2Zh85yElAjLLfyW4sXlc
Xv6KyghUBkJ3fTh+VsvbI8TpIwdCoHXfojGgSddyavJYLJGM/MIw40gKz6xXjMT1ob7sUYsBRYPA
Cik0XJ9RbwrQcn2keBNakfcOZLEI351YrVcF/UKJJQQk4ZCKySVcGbQaydfG0rFX4yYiuPxzyPFv
W2I3zxGC4M50bbftC9rSsU60UedjkKvnvOMSWB9q1bDymMCjrV4MLEshQhJAJFrTGUDraJqD+7Fn
UkN5KpnPGtLOscaqCD+IEgnwqj/gkSQTFHfE+StLjBtuD9Hv0nB3m1fzd/0Lz1wX0L4vM/AJwTza
JyPOfOZDoVboEa+hWphs1+VMGdeR/abvGcUjO5ky7PFLBmyLlLh0NcMlAONxYBsa2c7Hv633aIor
RsoaXPi7+RvwQAIU2d6N+kRjjHOkZ8hxBcB17dYTi1c5f0i9ZC6dziIRy7HYXcgs4WnHlSOE2Y1h
9eXDP2cpnEs1T+rmVA8URjMD8e7lvFphiROI17YU3ww4olWtnUL9PXvg5ceGr4huBOro7OQ6Kj49
LUzLRS9+tHiJT/D8c0+N2T9abgN56yv0Bhbw6VNuQZ+ivo9aZncVA0P7L22LebSNBL4VwzSjfmoa
mueFXlBGopCdGwS5VKwZurDKnXhZyzruhErPGlsgHyhnkTcTmBUmewQwaye5X8r/BXSV9DgR7Gq4
knOn1yFQm80dcB8952hE1ryc+KMKM/DnIQ94KZbZ88JX64Gf98kIDP0diAYN5GcPd9MT+iRHJFSO
v2ZFd0CwMWZYmb8EIuJal957krrQoYjsHM0u0bb1Ri1ml6koUqjGHAhEPdR5Np+1SNNLs5LEjxaP
xK1sEIHfa7xJrXkJJrVqCIflSF8wVrWK86Fihx+rlwevV6uownwdm9At5EkAQWy6cbDlxBTt9Zqy
/r0geRced6gAjyaKkd+IufMZ63M/WOWHpDENLbNWsi+sqTHwUA3Yy0PDEyml0sjS3s/edaP3EbTr
SedfpikYWwN5ucYdlozIRuQoOxOvuB1MVLQSJDknoZpcYMcFpGjjZuzVllElqkzxe0C2MEtWfVfv
JSHffkFbq7b3KPpcs8Df71WhQDQ5M8KXUcFcTK7Y2E3bA+V7MpD2qLhxFmSBBmhcm4Rbb9iKCU+K
rQ7pXnlExPJ1boJZjDTDgrXbiY55SNXERjX55HsqNayZyQpshXZGvSXA8yNMeNoCBDkKxJriRPm6
XflhjxwKvqB7N392+geEuRf6VsBx74XnsUHo/zFXV7kT8nAs6II1DAc/IqaeHIunNUJ3U4v8ir7L
0sNCYQffG8FD/n5YQJiGHi0fOErI1eyZXisg3TbJO5XPdcmpp5HO6qOsQe+fDkP1BJzkEbQqFEqq
wmXapUCbfAyPgo54ZH5ClcPU6U9t51tKI2gHTGcsfNB7oQdZLa6S6uuU3NtkXH14eqNQqmFAX0gz
geP0eSo2Oq1Z9myH/lDAv5C2i8GC+JCZ0h8mNrl+dhMHUgpvyeHSvce8Kt11xy6M9VWvLIz5bPza
pJtVQUL2M0eEl5tAH621qghswFVJ64JPpb84HQFMUksuI9cAGgwh2M3+FfkiqatVXsKmhKb06cyL
83Nd2eKPktDMkshWNb6zppS1pf/AplotBVrEru19aL6k1mhFTCepBO/Ebou3e/DvJ5LuzlMRBpTU
dm/Wafwma2yiK1EqamH0s99HQS0g+ehoi72XMSk4jg87tEx6YySThj61CUc7ewPXWZrFzskT2Pu6
AHKS5zSqt3NSKo62Es3Mu1XuupKMvPWPV+BGIBCU1CFjoUEegVLijts78GN1jG1R2oYwQZMuhNFZ
piMTjHCkYu3nHzC5lh6Stg8PCLwu1jfevLf9oUnEtSlRYdX21HAztKmmCL7bp/3goMPOp5Kay2uJ
oScJALD/Ji9ItEtMi0+8lRz31v5yE/O6S6D12u46EtqRxwIka8gD1p+6NYStqFmm3lTjiwaAcvIT
OLAe8R13KGKsimclX6MpLPLWze0aULoXkB7aUUvEa5N/iQkkK9PJ0Z0dN//fgcmYKNWh2liLPZDA
S9TcvoHPiLet6n72pJN8Th5YU+Qc8k6uQX2AFZL2kIyp69nFVGxWGWBSOy6HBKAru6aHI5Etb8+H
/FQoui0pK9zLUF4hM86b0QxqkTsiIBLaVZJ/k1AcQ49yCReVIrnLBJdfvA7++maOXXbcHl+A7ZA/
g21irejxGX1JY6SNnyRco7qAAwbdxMjvMcXM955++pqLGHkQcTwsjBmZM2OCKpIHvDBBjlDOBX0G
mFLeo12no+W4ciYTHN0EvJ4utRL/CdbvA3iGW/rIFjtufKDUoxSO6TWo5wX0ALrxhHftgDPWNNel
88NOR4GGWVaLMOoxguR99Xz/FAvLQJ9tMRV4gWCeBoHjITg8kqjnVrOa9IC4OdPyMDA1l1m5C1KS
2es6Pvy8UC4hK+UtvDyaD5XwtpScumP3mJjtDeWYDkVY4HSOMzWRmrj4NPLt1lp2B9PxVjE7BRVR
skt2EpZvUTS6fCEAQVGXKiQ1iASElHWKM6IJdbQt1xIKHyJNH96DtdNJtgAfxXIM+U+o5VaLpk3N
QAM3geAcpd3Nry1WHBVbCmwvNbP0a9mOT2lfKS+cd3qNiX+MReQylBv3lAsNHSfoHDLOtkw6H30+
jZ4IR8Vi2Q3vd+gdl95KUp31rdrLy9Le4m6AufBdxtoud+BHseIJkL0jIb3wOM4qHQVIyoJNhlh6
BlMfiOuSGxxuV6DpRsDxgz07EtQWD8qQ26g2dvDOi+6uyYRVlHmzLEBnXF7c3xlAfpTKapcK5cy/
NrHUQi0MkABr5w/F9CBxxV6j/pWa/bUwsljTswDf0zHiGS1IGL8mxx5PS/YAsBRkZMe24S0E/Vdp
jOkzcy8fldoeQOkh9vwvAqyRgvyY2mF0hPBSKYdu8u+Za2kux2McFK6VMEXuy7DJk3WglZKctU5L
bccC5TqjMSx7qTVLI50pWX4QpXhOgQub8t/EAxKFlfYvi3+8VlahMvHlM1Dp4FXBWbXltOu3k1Au
i8tf+3KGQryhJnJDdfmBZNdqsh6Y0YJ3KuiTBFELBXC3KCWsap96W+YLl0EtLTuJZ7DRyK3+NW//
rrpkBeqjOJFZVaIxT0dSnGhBUvuQJ4bxl0JtoHc1rjuQd939vltd249zklOJ/Cqw+XtNk78zQylk
sCCj+fnGsB2KEZzIgsS8va3P5eq0hC4F1wirDXapo2lo61cEyyrgRNwto3E78ojkjZOdIqM9ZSB0
V3YsRNbIc6xaJW/o7WGeFUntRV52AZOviDxj2zpkeek4tlU0sW7mDrwYIVKQYveLEVnx12wofw4w
1qhqCmmgr1cnY5Zulc+1QKUx0FQ6nQ2pGl6q2/aynfzlQddrYp2nDe637Q0mvV98Q8zKl9Ce/2VM
36dHMEUY5gXC6vdKxiGt6CJ80ePWvIt39YWAk2c6eqfS+O6mtSaEAVv0HAFLA/kEEydzq4LyJzsv
85rDBKkLgoi67T+MrNU755GSJvr/H7QsvMC5kBcxX7EDpUy1htekxT3zCnbRgC1lZOMAfW2IwpMq
nbXsFdK1j/8JjXODc+Nf5QSKApx2Ed6npMD9F50rqGPKUl5ZY2ku+zphzH2eCjqMvoZCVSGbQzTm
vXf443fiwv7aFt/Wo+QhEdBcLp22gFi0NNbWlUy27IXHAUhxJ8KFc1BlrqIHe/V1RDdgRHcDE+Oo
p0SeSzAUnxj8iFJg/grL9mRl5pHvCpfYnO2gNinwWDm8WgaZ+SfLchhCqELmCScUI5X/8vGylOjA
hj0gAdwqNnMDgpz2zcmG+9ZPIfenfPDenmHYFhYbYj+0xmm33Lj1APH9+B0WyG8PKg5rmf34NOV7
GVHGtSN8kOKTtDudf+5gMMhqupytY192IH+QSnTGoP2zOKHwC9lzzXa26Vfm08TBDHy1FAQW2zE2
tZHuyMIpwgXtirRMduyv7q74FBgyLCJvWd0HgMJnIoyx9Uqg6XNz9OW4uXjoFmT2YX1ziLkDSsM4
g09IZzYmITuVLaboIncUxMZnBUT1by8U0ATXFMO1TFQPB1bQyhZBYm41MAqjJxajRwMLd5+fr5EQ
yCipwAMOEeSsYk1C/npGyXh1/PhxsRlia7H2s9L96SSR5+NzW0Dtss+hQcfkKRzakfPiRFVcCpsG
HHDxbUP+/vsQpaygGL6xhExgeaMhS01wSnOJq4esUcY748Vc87ECFQIy5/Fc9E153lEfgTEaJDRT
lzYkCEVqEc1zoG+2Tch/zU5+1bLewfM1Qh0JaH7XxrtoyiQzNvQHySR9YisCsSfB/hSphNJzdUiB
Z8+YRrzL8MEFHtv2wtdnOF2TevRbvWPNc4+aljzQBwhcnFRFNCl2hVILKsL23W1velpV3IPfeFlo
5oOUOhZ46XTHi2/T4HyIFxsbcXUGbt/leMt8P44Fe5qSYhwGj4YiO96A6S3QBVjM5/QQtHDbK5Nb
vm1psexSLM7VN+T3RKmkSBBPLb9kA8UQbF22TtCyNQdS01Upko8mhbmYZv44kwrpp4toMaQxtGSY
OE8FLKsayBpApjkAwboh/TygP60ciXENk7eN2PvDi6+7DtTi5Nc8Km7+zhjTqgsPgsYS4ST9kCmg
NKMoGq7gAoD+uo+3EJ97C07Z7oX5QvZzDsyvh42iYCD6Rx93/b889AqXT6EFzbsjfj/S3lXIaagD
BW6d1pGj2EMx+L1wxiK80KY7S8uY+dYGvbh7BT3GwlhC2Dg4px26YtMiyFwXDugmjhby/yn8Aldx
slQgvW2KKGibfpThBscyRlU5CAG8RZ7MwC6drlL6nRUy6jrWeQMS9yzJzBRtP8HmzpEtTi0zreCf
YvzKSyKhLLBjtrhKZefuwy3QuRK0g7NEgfba8iS2K/1GEAWhhNk+cwzssKYh0aLxp7QldarAkckM
TNHe3znNv4EXxsbI9yvD+8gP5+AIWynHNoQQvJzJveeGfPCT0fvh6iLQ9jLavv16QyrIntaKONFC
N/ZR5Xw1JrgiS4L2nLNb8ruDHpPPRuIvbVd0WajrCVOMG250vbRJKRGCI2ZcH5JPgtF0pmssqyGA
0P+eMmLPbeAUmuJlSoy04nNf04VFZ3jRKxh/Y7LEHpmu7MscVKPM2zN/cZxfMwuaxMe4S15PXS6M
ufTvIZm3xmRsAIh9wzDd04PD3lOm5HYx5/PZwSZSoZJQhjLHM+2HnzWz61Yihjv9A5zqvAZMpmvL
HOmSHW2AwvYfaxPnNcuAYSgozcDXknJfCqq0DcjeiQZV28rz1EgcbRK53gAl7la4Iy05KayfnSxl
s2yJrGnTEQpV1nAXob8odT/wif2iRam6GKX3HsrmYCszHu4QZYwFU8btt+kqj9hDv62uoGcqkNuN
+AM7azHGLeDLYn7dCcgZB/DqYnbvh2CDU96eSufCpFiouxjCUIhIhWcs5IufzasCTTpw0R2n9YZU
4tngDeVn4FQAMH+jqxZXQVJiyToGPUx6XhJAOoYqOH2PsQyPABawMNMCchtY1ecTMlo7c9efI6E7
w7OqUOIn9RgChtH4wLZo0FEfRIrpf23/qG44NbHXL7WWkYS1OVwI0Sr9YHd4kXKW8fM8nWD5lybT
nN82dRIVxWMb97YlNaG912L8vr637UkQJoeXhjPglBcWRRG3+Uo6V4eRT8CpryKGujzhpPUl9yAl
ApEQE7rJ1PeOFXUg5WjmhPAWaDdDpnb3giFbhCZHQI0HL3kCLrnjBGs3JytlofyMyTe4yxRvuort
a1p6/IFaQ26NFOZ3uhH8mzVDvmpfS4CsaY9qTz6tfIlovaOocyp3WDSuczDYxpbf4PtK9u1m8KQX
/kEY2Hzpmd+JHqzwxHV+of76kT7aLRj+YAfg3r8vuDBM7GESyWA/BRuflg+V+b51wE48ay4nXE5M
hohkLOjC4XNzCxYS16p7FZCPK/wIE0hCfrrzkK3Ff6ArX7f58Qzu7lSLkv5+k9JatPuJ8wELec8/
7eu7jMKjK7Sj3YM6kCXsUMJsYt61Id7PyNe+lY1KLcenlAvG16gyazRP9btN8qcw4cYUtzBdL1jY
eQV49Lk5s2Ff+fvr4p6ELbAvxSgGcBLB/ja+9FfQI9bkSPozwmn1M4p/WgDUx2bRHC53x2i+FAfK
tO0L1E9loo2AB0adC2kG9OJfyMdvQhUQXZmV3rlxorSULvuUdAbjPCj7P0buWXj7C7QA4+AfYC7L
Ym6ylM6SsxqcxJgCQj6QnSTCKmRF21qL8eek7RM1Vqp2grC/cNGh7c7O26NsOPeoUdtEm15zkDY2
jIk2O4YjpvK4tbQcp/m9nb4rkpOyCHtSkwTObwzP/5u3Y2Xxupv9eClfya2KNw7RZRaKeAZ3rtg2
JKthThPo8v/BubIZ9WpIZyK0lMeDllLLYUnsxtrWVdybVXPBr0MSPrhczDr2Y0lzSuc67QVgOMzt
qfCJzaH0zF25f9nVEE8H/WAPRBCwVY/FwTbM3tHXKcjnegBtwaDrG7hNz+XNkKQPk3cbewcYAydo
+rsy4HYpLeKnHlpcCR3ei3Cs0V7gVvhCClahann/svU1yQpvO4vjNYs1BWijcd+ayTHvsH2+BhFF
ChNwEYKI0Qfgn9Abv+xh13vPPfaMflZNd/qkGyLD3cGxz7mvsw7aVMevd4xAokeOAQkuD/PZeA1V
i1Sd18/F5Xmp3cz/6BykeqmiAKACRAkRXNuh/QuDS7wDR9KN/LYGHwsWQ14Zx1Q4SCKwl+zmMp0b
1KV2SKrWIzwWoRKp/EULUtnst3fACBINZiNM13eIRwSTHKr5ZuC2fXyLZYtvqEfb/yze8Dl94o83
LVatc3z51DE57nM9TO2C/vyMwE1gvPB6T+F4GgpqTwedtQvPmZiGT6VAyeoac+6fLguBW6f4li6J
oQG399Pg3ystH3B5gnM3k/lGEkkAvyCboJQNgAYmNXS5Va3/lVfZCL9sbgGxVAbk4TFbbG406pGC
BXnzPlUICPJ6pswtgMOVh+Oyz0mFQT7a6H48B5kuUbedCBxwDIA1PPYmWROk1uNEWW+4S/KWmsFR
NjTtgHsAMPj/uc+e3jbcKU/vIA0JCBMcyc8QhTRsspFC/pBFhzYMi9dTPAYrY6Ug90xUAC4p4nUA
MQqQsWSXlyPVIZGbH66lmiAFGqV/TNtqvU2y9hqxA6zobYwnRG90oC2rNTtozgH2O5Ad00urnYEw
PCDbxuMTngn5Mc4K8w/vNkbe2EJD0cqdp6f6TBnpW6X56+zQm3kc2J/YoIAUIT1CkVmPY2Ybs+ty
DB1Fj5D48YPOMQIhHXsi9LVEm+gF+p//Twp0UBDNn6S/20PlulL70G9pYiL/KHm4At0JEw/u0Hdi
P+GS7TgmrdTN8ya3ezoH9NsWqGpXfweOaRUWj8gwxP8PfsBFTOcfZR8IzlpK11GuJgjkxi57bd5y
u+u4ziDIRK+nVWWNYVMvWAM0zYxo39ogwtqt/j7LoGuDPE24+RmMX3Sf3rqnoLweNs6x06ZuM2AF
E8EAx31LjnR0SP5LRmsYPAbmUnoG4nIaLklJqn6iuHIO2YXZvJECy1ti/4F3j2bx77Esoh1JQ/Ul
DVWdAoQdChSC8c7k4OqprIA0NOx2PfsOwJNq9ZkmM0UOGpsr09KMRFzRyNvz5kMdPlH1XOoi509t
7TzNS7NZBRCj6SbLi4DIC7ig5pTf2qqwECdthZCQ3FLvpna/gL60PK0xVi98UpLmUBP98eCePEC1
W6unkaNlSSZpkmUnRyI4dyi0He85wTucKBj5xX5y3oiguH9j0Qq7HnUUxW22CgWaLqTrvsoYfOL6
Vz+vH7NgaRPjtD7v27g9UfuWktDICZ3tSLtp1E+PDv51Z47o5qm8aonyjCSHzoWjLLv7YfASsJ+n
7AbILsjx6VKdDmtSJtqwtF/B77xOzl0Jmu6tjeAr6yRhhABGsCgB4LZWzjxXj4iPI0jPWBpeJn3F
xzI3QrlK2llLz1N0DMrfuOHJ73cSAKBXBhjjD5ii2y9+42Y4K/XFyGH+0vSGv7lxyhVzWGtaO06/
yvScrV9oUKHoPA/lLEMFyjSLktXzjvaourw9s2UE52TsNQMDLIETgysyImhpbSJhVrry970KR56e
3mvygBFqaIU7nkjlNwZ6knKORyN3SPs78k6T8jxEackUwRaMqxrvp6ONYEI/lSS3I7TSePIc7PXH
AB/JXLgOvbxofLlE/nna4y4LGLM0tdpnXbFcFZdrQQlD17yha6HIRaYtvfLUCE8OS71kykn9JM2k
bOZDH+0/URi586LxFrHw+xgFrwRANzTkfcD+74N4fGANRq2/y7wFrlaJut0EHYRiXZw0Pg2wsA6n
PxkG1IwceZ5bd8LIhgyPfFOSMowBD9uVhh6QU8a6WCNoXe6HGp+0Yovs4praXF/r0UC2j4Ll1r8P
Qh4b4gFpa11ScktMfA4Uz6Ulo8Ze74HN+R96QbuC+Z9fSs0sSBZp3tHr1S0e7Jogh4vUSK9p+w4U
hFP4rc2GPDfUrfR5N4PGxQVu+UmiNuDTwBodBj8jOcYuO6QDJNELHx4aI+1i5nN1t28Lo+7Fdkrl
/Brb4rHcC+dtRjExWmV0m+pYrW7ykTDvN95WAISyyjouw3tIYEtg8rwSCZIs+2AkEdzGmKRUBl6b
5DeEwyw2WVOkQJTCC1ZV9HPGHeCRSzCmzX3VjdHs78Ib3mAgep3Y78dy5NlzqKYMV2HkjvQzoAUl
v2Ki6hHdgawkz+1CmxMSqEvn+c5wk3Y9YPG349v/ofe0rLglyyDF1hUAKlJvhg9ujNcz9EbIdBHG
8A7ARgc4y1/gPtlPAyHK8VkUk101e36QGEoN5Eo6ucQztIAJfL1OhfYlusgLqEk1aQtOSALWEVLv
TNH3Z3byZHWQCTn8BuaN2lOZ1aEDrGu52LQU5DLDyNvwtkX5awm3ebM1GtG0fFdPU/qxkK43oXM5
Xy5XhXmT2ZgRy1S2MZwcMo9xGgAdko+opTPwx2LLGceeBJdHw2X4WseefgXDExCQx/AWwEQHH2sS
otJwyw2KdD7NlFBoGMEiIDVxtWteB9htf79L4PcFj/G/QZIIDC2KdLPgvjd/6UCqlLpz2NsRnu8J
w0tL9ru4dqtHYw/dCycdnK4hnNcLjjG1vhqKdJjj3/UnCzynnVqPLboUbudmayLLX1A1hIXAdQFz
e74ga+chhux947niDNcLYYRP2FWjSUeCrrhfAiFrgBJ1KqNeAtCe1ybmA0kpUAFiu144Zduzx5ct
jGCb3oeN06b45t+1mfhwKGgsKXB5xaNWu+FrRgq5egj1ivxA5vGVgQUZTAE4THscsJ1vpe6ZMazC
7Bgod+Sy5oScr6jy/u0I4+ZAB+786UNk4YBPHOU//otpoU13UULKQzp6xMc6VjNNEl4RafYaRH1G
AqFdgRdNQXl9rtOEkutYoI9qlqK+MCOrXDvAvI0rw0/FQrqvF+E+3yMqBC5VolvwSoTQ4lOHJtSw
X8AS4Yzp9XlkNJtIZ5UUsQGdmsUKeKJvwlB+v+uOsLDNDeyBpuVERAevz5lwalsP8VxZ7MHdsGBK
tGxDAQlJTW4IKOrmRu80sW2wlQCdLPGbmbg0Er/PF4XnOs5MeBISMG+1FKMuEYXCleaWZTKDxH+Q
enk5JxIk8jGK5YZEH7I5pzNtyYfa2VVXN5tsKYaxXxhTU0lU8nzrzzsMA/Yrou4hL0ZiZxso+T0A
XvTi4d0yp4omNDTmbEH7BJfUpNUDk8dV132TCyLljbCYMrdyyPd2UvBV/DRItgkv18DASXv7ZH6L
DBz5DBgnJHO0lhIQQT1F+2VNbT2X6qJpkMRFxkCRCrdRxTK+jsMM56nUcqhaXjoWwTQwwjugSv35
zksp8clrvUsj/AAyLftee8ziUaMePFX8nj1WM5Wao5lYrrPVZysh4mda/+o3IWZGl+FknK9Bxi1S
z+E7eTc/FNT5UL5AdPxi4PIcUYfpKu6txTBL5i9Qas5xaoHbmkGphFtK4GG4N01OhLjyNMz5ngiz
0AcRp0oK9Qe1BeI/Q4+mP93yFodFkmtf7VFDJW+bI54M/VmmEbahqww0qp/ODBZBS7BdRcbo+VAI
pSJs/5cN1z9yIXiyoxiGIiz0gD4w2czxYpK2h+7haO84pJavXPmWargDyWy14oYRomWWgN8t9gOo
GS14miM4n8JXC/th7Qj+ENmr/CFgBU2F8o3gO1vxfO5D+BPBgZfe7AHDygmQUqp4jCvBFm1nVIN2
sG7c+E5+ffhusyFRIEqQle+q1vBYifRoAewEC6DxlFp2esSLoELJ0GZBKweICIKEXVpADPYQBlmL
qRmudmdI8rxFGwahCFvCVvwAppRKyexFzQmLFF3jO62fE+XlbURHoPdBS6DuRdIC1G175C4kqp7C
Yr+mZ0TR4rDdg7D3P3hytRHVYrDYWtQF2SB0bOnW2nAgVlm5cXVbuy+9JE4F/GCEhjPY8nsiyrKH
/rWVcws6VzkA4Z2ZYw/Fe6Aw0rTrJoyzBcoTBlcqbWyjEk3pwtfKpykzejPZu3Ss62k61QXcrBFx
wYUgkcFrb94xo0hF81TYqkrfmL+tRePItLjANNv4XQ0ZJHizqumiFc+hHkKuYzmS424OAbeHuusJ
K0YLnkxNTo88Ryt36DJODiRtCMebHLU8w6u6K3bShZlvE7lZC2ZtM/XAWlhuEJzX/HayicOAeXBd
wTQ4Mbsdu+HKe7ZaJnF+iJ7Ps5grrBJ2cN3rENDTvyQQJe8D+/EQouHw8MpnYLM5k1DsuaTPL15/
XFiJHfCN0uaDm+3h9M+iDYfBO/JAnQouzj8euOcs3RP9/sPNtbB9UWSjkS8oeWypBJHBNUcTprSC
YlefsnSpDbRTWzPfW3XHWmn9vUAFnPUWOdThAy1zQsAPqwmin4U6lsQ3AUhP3IhCdPpvYHDyILLV
65M5n9mPie7sGCzZTaCnhmOHzudBLOezu1X6VbEYXcuRTtvxTx3R4JKZ59RBIbJ7ECUnoNVNYLaf
6wK0Ngh7dzusVYjXOihe8KvSPCq+bNBO81AujFbluzQE7ANFeZBfVdH6zL45n+0lud505qHmAn7i
/pFrn1cB7qcF0EvlAqZxN7IQqWiOJvhJyHgjrR7wN/q926pALCXwjLRLsaUdtbiXlAYSkhE9vSr6
K6Yfkr0Gv2DKkTA7g/0HBoWbZIuDOp7Vo/a3YVZZ58FVVrXKu7QjZFibjnER9SIABG2TFFOT6pML
njigSDLsY9d4q4yiXPe9igldKHFVBsxuu2nPxWcMIR4qg4UutKHuN0Ze3t5Nut9YDghUP5HuHuwK
1EaOpXxb9ay9FAWE9ZjTByPJU9ZXZSe1uRqNuzJ8bfBCzqDSeSEd/rdSImC7noO018Ph06q4XU7T
Q2JknHEzUa/nKEnxR/C55GtztjVq/IwFRcEjC5Jx4TIGa/Ph25AFXH8vaLXaTPHdLJglGQBGQw3a
0xU7+mpMIKBY/BdnPW4n7T4GrTAeA3xjgnCMNWDBwlk5bVe9LWUzBAqZWltZb2qYlHiv+L1nFL4r
LDicw4fSJzjZR196m6o27iu0bpGvKCS/ny7zT/LwAg2kyrONtZw80DZpEHFA3TLV9xeSj6DasLqA
3MXYyDNbNHiq/mfLfx+uBx7mWxk8XNy4/koTC7P249Q0OxkNZQ56aI4wD85skXf6Y7FQykxFZtNd
VORw6BKUkJ5glgvXmjVKs/tP2w7h24qm8/y/GLsG/3wVij8ravKm0rsGwiNyEhQ5SRSCqgL5eycm
+gXF+cCik0ZwQxeQ5vGYt2yahD8xMbyDrkIlQd+6+d0qY09TtbrCSso1H9bYM4PHcwi1pN2sEhUI
u/KiQVorY4p8VrFllI56nVfoJsJOZid2zN299xV+OyGiTmz6kuwo9hbQbriXNOim21w2WaQmtXmC
3mO1nBz+bLoPydV/frLryGITDSeEtU/x1/1bvOfZIfNW/9N/KLK/H0aS3oIRUQVwe9nnTg2hesJl
Ppuh9dOdvHerg5k5bIw1TWoUth8d5b9P9GZw06iYKSRZMeDt8DGg4pQVkDW+xY+7cDQioM+yME55
gikiHDXfwOUGRxfXvjHFCcRrYpgcHsLVDYZljbWUK/5JdjvGtZHKlDQzvMrvTnKuLKCmC4iCh58d
kru3eNKcp0lAN3JSF4CNXQ2Mnz7G1szQHDbWsZnkpEsfSlgGiAio657aEkZtEbrROnzXAIvksBzV
h/AXqX6FKhazZpS2MQrLtGX15bpA8IAhMauFPq5rhB1okkaCq59nPfXdUFv1lvHnRU0Wxw+omjeE
AjNaXTlGjE8NSZWUr/scQvgI3gHanlQKbfbRBcfZb4e6iToG4Rks0p1iBdUDoei8JTWIdnUPzghG
R9NAJ7CeWcnfgMQsn3HDyQmXDcO4fQDg3ZD+Pt0ic1I22YHrfgiyyEv3UIlHqiL61TlQZfGI7A7z
1Tb1l3jDa5CDztVtrQaBWKhRIzE/SAzed6JvmjDRYw3vJ95ZQauz+FgIGiTfza172I/LmaW211gb
YqJnSF4ekRpmeIB8xNiAZFTOV4JDTqaRG3sNtQ9rLyOKhNQTDW78vw/IWUJIwsD/aJkzzU8hOtVv
NsG4tGiqI7sRj1TtLZFfkYSmHOiJlUTm7ikOLshoxyEUke1F6XW7TJ97rnhfDP7SxqGwYhNQR7lQ
dldJHl34fHynklkGccNdVHVhRXPRhhlcocHf+XyZn+Wg3nRZF6Aqo3ujVPTGIBba36hnvWa51Sb3
q0y8CBibiS9TSwij5OhEDumHV+4gbKwToSTatO3G9TR0eflIxsd1dpNQMEqnkke2EMaP9r3/iqfw
cx6uw1rPJRo3ckI9ZQ+Cb87cSWPKUENBLl0zav5rJQLJWb7V2z+OgfgXetgaDS8kLVp+Ou7qTcXd
bpGaK8mjUi0JWWojmh0JjfdOw5lc20xmWvDTNlj0VAX7SZhgUtxD+b09OvcQxyPLwgwW44zjNr8v
yB641vNPbqyL+hTDWbK7rZ78zfV7ICjFL0c7WEbcxCyljVUKVLnqosJpCN0AoPlQ4h89RGHuqQnh
GvacSbgkzYqcdHgsAdLvt+Hw4c7XEWuNw1p87mSNLYhan9E0QcBt7JDorV4w2dC6ENUfRxo0omm9
qva30/XRxk69dPzoxFfn1LNZ5KK3h5UYqWLwmQ0SRxyET5BOEXLWbOpkR7IQtEgB/Y4C4UcdmrZK
njjAI8NEHYI17F17xb0s7gYWdHoF6ec24PFBo4kD0doYYQ30+Tt92Rf804EkemTeCl8fYhUExcVm
6V/YNkfuxVuDLfGG9v8B90dK6svLxaM+ADHaVergF9W3+pqnZX1uMmLEjyMW1db8T0xzpD+xCMRG
12xYMECHjA/jJxyf1LXd/Zwur37pewWKin9thlfg9BgX0gxB9nBwNIuESWBTxiHZk4v+ndOPrDkq
ArfdfC2K8TINughp29hG1wiz9xcQ+dBuJWK8YR7kwKddvp3KKuwFotHe155IKgAXJBM3LDmVvevZ
NKkVVu/HphIJkCpt27RM4XBvS6bepqoXuuKsTN9IrJt3LS0d33exLwT6oOyUiWxBkjOJ6JuGdT+U
nBkvaeSkYZPgtP6u4lySDct/vqUohHAJWsUxopLC8ERRopKS65qJuHBS0Q89SKfaXJW+Ed7lCKiV
TPk+TalokteTMq/2gCsa303XFKgO0DoFxuRSDVdAxL0esfx/1gxdQyRLDV7XmYE0os3gyYTqxEvn
FJaDpncw1/uwgNvFQqUykqFOqjBY9LEAXE/XpDsBE1cgXzAxnCRavlu5pD9EJ9BOpLZYVrB9c6kA
/V/dtRWIohhaNkIWj5yCQup2nv6+R0rJvMYyH6EDLv0AsXG9VUhhBAPcxPd2ZTRsLojuQTPAHfPO
QBtTjZVCp3VlpvN6uLrgivYFFV2pMtGJsNImiXHDkvrZsOfkNb6TgD5qy87j3gIcF+AtuOnr20p9
H4koewCdfxwh3DXSXbMjESjntnqEvFsN7iesPeaBJDGZqUGXG6I7LAWHzxFv4ZDzCJdg9Y0Za2d/
pZuzac0BfuBOmx4/DtdKkcgCGcZuddVx8UC4MAy05kGjLapuIWeOFNFdSYWHfd4vKh9wm6k1apWm
lZUdcbPOjQ9KWU9BA7HO+0PjJxN40SoEKTiS6soyoKn22/doVDd/KiEjmFABHZ88URRpa3PlgFV6
snZaFCcXYjINeVs8+V+CJnrNAFzMDM2tYWnW0QdKUFF4wDsMP0FDu31JUC28slPYlMkCqOfyFjjk
nG93tYAO8zJz2zDd5MJu3eWiRfDy38Ry65VUJMlIv7LUI7AfTXTdgxJz5+Ps1mrK+A8eq5szD8ak
wOYuF8ABTx813o0ESfWxBAm6jJJAD9M2+byiT8tKbVCVwbcpuSo1tERZZNtcDF+NwwtatncT4IN4
G4h0YdwTUhMEiKNDI6AsSyBr/xbo+k6kzSVJ7M8NISPCawyUeJmtDUyVUENeF1r15SUpuE51CrwW
QWDHGaGSVeoN3NqFbaLFtJerQe7kxEw9HWnqteSmcDBzsXafmty0Tm/Wf9njOD58DBxEl9AaILxT
dgBnEYxL2UZxw40SpHq8skns3XSEspz9xyBC2L2ZQOejWRDKfqKJji8ppOSgMX2rcf1u+GagioDy
mkcYOYubFcCISlAugnaZeVeHFCUtsO9mTMJaE6d11PeXdcncCzrxJ3LvQOFEdwYqnZbRUvmQSAWh
0S72mUrzMkLk8hltD1cAUaMmlQd5pPlX5151BAGfq2xG7B622UrA7qqqMaB03iKXb0UPXzPMYwRc
RBYKexkddk7RkjARM0blrCIUdS7oaQHZR7rmhsgfckZUZMyi8L0DQjPigysJFeYIWa+MYPj3UxC5
jQCLBVckrViIJrRU/lh9Ba8D3E3CPbeeHfaL5gtrkSMFcJ0VQ2Kvn/B/i1+RnicZFuVcB7esgPti
PVLB2elUGiRLUMQApv+zbA15htD/FP9tMyOfPXBR7OXYLlPt1PZ8QMsVGej+K7v7spzXsxBec6lP
KXYgPdri+BdO99pa88ZhJ9+acW/3Xon8sMMtfT6yLSxBH9UKNwpsUrVxU9CmfEY6bkJgPw4Ye5FN
1i0XRH/n6CLkqYvofkWPj1JT1bYnhTWLtRQa2aJyU7ZV21DfBa+x18yYoIgTzWI7wR4yL7V7zkq7
HWEMyQEtUTdUALhSP3dBmX0v399cbpiAKqdvumipGOTFoKsrZC1ItK+tkilBDipSh5JYEOeRm4Q+
0UiUWgwPY5ZJeIHUOE49ydKZCnH2jN5hWnpK8HvbE4lS/oK6JZtTB3kyqFdEOiavDqHtV35RmC9T
YnLL07Xsr18SffdfM2NX+IijjpFpUxz2gcb0HXBivJ/uC2kXvSrje5kO7epozyA4llGkuPNDkfh0
YqhDhFew/O6aXDQ1M30lLNrDDLx30yfOX3yyZzDhVE6t/yfkWo910ZUPwO7ruBa4gqt4Hnt+jxiV
+pmfhk71zMXA8cdQ6cWLY11TLxCyyRL3eDZdqHONnEdK17JxUIqqlmplqgHqeQR9ZB7I99v87ru5
uqLwFsHxb55n28llaHKK0JX6kAfe6OpBbjm9qhfmO2lnm2aVm8e0nvj+y6nyZ9eLpMuLZS5uUK2u
dZKpB9WS5X9kgSBDF7ZxVNaxi7McJURCNQSHqc74kXLqBOj+e+PtYKSYVoWqoPSiKjiMw+gN48dC
1MmMmHxauf0zEuv6B/nFY0HLNR3JRx5bzX1DBRGWNElvgU2yCCoZWLr8Iwe3rG19Lo119hYypOPL
PfNf4EYiRVn4VmByenEAvyxBEvdAUGV3WdymFz5r4CSvwM0DUrWGpWddJ8tTrlcPw6QUWygLa6I8
1gnPqeofvcKTTFex+UQGANv3p4F4ZhqN0ae1Zn41P7r13qXCic4SN+AqWC+SiMFh8PYfJrnD/S67
OkIqwoqSiMKqn0keGunyT2Gt97k0WS6iUBF9N/3eg+w0vKyn3w2Ggwo3UedpL2Ai+yybaJ095vDE
+p0UrnIRmmtfU++5eV8FRtCZ77Cr4TKwmZCvGV28A3qKL+8lS4mnJAYGaAaR4GAZWhuVWitd6Off
dKb3jf8QzqKtS4naYimkVLJbgXZTjOHoCZea1N4HFadeNOOZGvUUyz1Efg+BGZjcv2JvTorNlZzP
QpGi+Ij9joKVOztwvJNYo+5RIAJMyDMWKCsYEtnEr8d+k3K3bUX9bbvUYOXQawaqaT/M+h+YmFkl
umVUPRgXDHOiy4anSiE7Z+aXtat+KdfLq16zrOhGWLlSwNDILq9niOH6s4EjJsmAHQZIH7J+FYtE
BTGSfqdqJSF5q92mb51dLMNBkEi8DXRu8TyLykwqVhl8+K7qzD2i2wvrANMTDRnKiHNhuL3/9UlH
rA/JCrcCSC2FRKNno0OTHgt4htnGwr+o2XtGv+q4gb2tbaAge7iH4O8k/PaKpdNLuRUOyzUzE57a
7LIVPluWwIwolhdldhjczm34hna7g9qokuR4R0ZZBWfKX0YAN9oQzgLHIKSap9qX+N4LJ6Vas7+6
zkF89VqYFejaOudBjtNtoM6FHwa5CdY2P3ZIXOj90GjJ2t4Yg/4pFF23YXfQ/o2oenB0SfzPtVLD
NVAwEHdl0FKRB6HQFqzo6yrxIuzLIOmnpiGZIVythZ6Q3wROLDmhh1cXqiDu6Ntiddro1a0QHKgT
14n6lxVJh+O4LGNuW/MKqbjjzRtSsv9rLBKtvmjkfFmqldrk6vZNrPvwan5dF2NwxfqjH895GpwU
YZEtnxpKy5+10vRsQfAWwCfTB60avU8iUE/LZzSv+q7VrkTKOzZXjFitkEzyxfGScYaKu3hWfFcW
3j7JDyfpGrdRSfFOlfkXJwv25KZPHpGcytxNfvFxf+Q92wxMxMCqUhZV71zqbqZlNTOjqrepodJ8
N6Znm1JbrbQeYKWbbjbKYS0ex4q3zt5rFoctdGvCp0vrXhiODpsdRVJ47tPwGi7ArP8WGzkqEYuI
+2OvkzuEqXkB642B/W2Lx+4YiEt86EbrSIn6TYdPohkqLDiMjNYBLc+P4EKqWY82BM5ekYEYq6Hb
CAMcH3VhZb+E+hpavvOhxe7lDDufV0m+ZZHcNpokVFVFo/G5sqOKWWZwiMegKSQDCBKbcCiR4ktz
bocBcG9qal9b7MSAMayd7K1VXM3Nf3XBc1NaVkDsLsYJZxKcU69V2mavsBZMidnwGCdI9hahQj5D
T1xWpx/DIRQYx3TTmO4HyYkjxqIbIXut1PYxqbza8thZm/F64XYcNcbY/amnmJ0oukHvMCqxexmT
LgVTqBLqUMZUWp08RWetVWoDuLk699mElt84zcuPO+Ca9IW5axjDqNVfqZI044xhx2gF04TI6FdK
UHH28v+TclCFdgIA0lCmhReY7SbsF9m8M72TO+Gf9HVEvSqXEC7NUZ7IdqcL+cuzlh0F5uZXzcrR
KVEbAS2bmZIHhLldLw4Ppet4/qzjKRJehQRsIwXTr+RUJlLEXlnTwDa8r/Qe4riX+PNugUMrwoEi
q78D3c0HzO8vMQecC2BUVsY/kFasS3hZGcIOkqh7Lq2cUG+7i3WvcyyWgQ4EJMojoBKXWmgpg/SS
suVuYrAdm+hOqYWcAoHWCs0SwF5S/L9xP+N2kqXxadPDsMEtXM34k+46MUVamWeHfxxbjL4kWb3n
vMGKzunhyKou4xY83R5KLV34mD8cHjCzPWqR++3sfVwOcrvJbhuYy3IRJY07g4S/wNdbiFVrTRfm
jCnIIGVoFupLqzxh5aAToldzPr5ZCC5A4PLMarS3Lmway2P2Kz2bbjr1KscjGUdC0FtRQVDkQpKk
0SPtK2yiO1/+jzqBKldn9FZ8putetTQySFESIQBIV88q4Jwf2yXNzw3ddlsnpM0DotwdDTSn2WRE
mHvLiikXnpemcXg35FCaWL2pbZrzPFuYWKZCL6eNqA22+Cb104/iqH1RKaWI2ML6MQ8I88bUSwR+
ZvrYXwDlif1ZLHQYsNk63fsGfl3NJpiN23g3tnGTk0lPJVHmkv1te6Br8dDJEV7vD+gda7kaTD+f
TY17JSL0SwTSavnFabvIXmT/qHp6LU1vBPFcneqZ66Ria83ZEGj5gPs4Nqbvb8PdtKuHzg1WL+4u
SVxn12pOu3rydWoYoJuSxitAGL3UINeqV+xqyse5ROfjJg259v8qOTA70Ji/LS7DWe7XXsJazx8f
mjclUhRmgYJWBmGN5VJJSdDjLGKFZ2E8jkQfSdW8S2UZqh6+pfFT2u7OfvC/AWRPzJMid+19zaLX
VzRZ5wvUYyP4v2XprW/p7DRGVUqAEBMIcb9iu1OiNE3t28thyJScomjyKig+aYSjTKUIokEhHW94
OI2tS2WX3FD0BRlNiSvhLxS8Xvqy471MCkEECJYGozLMFr+8CIU7OmHsnCiWrZP/6E2JDJ5+qt2C
u1reOpK/g6ka6p/W7oLoOz5n8q6J4eQIS4AU4vY1G0H3igCp0JrDxrUfMhXprAAfhS5IBdPPizv1
eg9ICduPF+40PTcvXnvH3MRyjmI4FLSrPLnSW6/e3aGe0y/m93ATpIzDCh44mWeBkqrot3ojVvmr
wNfCrHQ8YXraxNbWAVjhUitTFaLfmrhDEFdJij/bU9mbK1uyLkGfd4Sg9qbPwfnStMmFuXP8tMlb
3374Bq7YVwiq8s9iHK877DECbarmiVjxcYSZERXOhDdHNLk1xyHq47Kj6Rwylu6N2f4U/GjrY6Bv
4t6jfilSgnnnT1k/QbVE2vGk81wRTGeAo4fHDVknPF9MzwC9tyL1bEsqunwKKUYIozsJQvEYcCn2
GvFUruQit96PLb4mvDs1kaiwOnr8gls3DyH9YfoRmq7bVJFEfVve8Y73BGQ0E7xNcehpvDCGhIVI
/scgWanquydSGze73hy9YFk8AwW71F17AnC6bvlu89IVFbvzpUc+cqiTaO81c/WoR1XDe8SUV1b9
qdalVwwzEPyERjHDSQ2qAmcWZszGi3Cg45FSTuLik2FWd4Zk/vDm8PgEFEoY/4Ow4jMBbiTglbTg
gEURyJwZVjzr0JafKZhvHG9AQSaJc4qymJiO2wQECdRfTO4PXuPO/uHXT/8MwkCt+pr4XWImAKWs
Pe3RY/2ga+V+9gBSi477aVpQKBxGPiY6GxBgBthTdc4V6oBX22PVqNgy6tGPORy4G1KTCn4r3Ssc
I5ubrfDw71y2B8ClbSvjzOr5Sz/JX1EZiA+C7oSlVoTyucduqcQpTuG4cSMxatNUF1xivki/6Y7H
+jRPviO9WSrvq6Xr2JV5nRnuZzn0qfRGSBdY0pOs6ZMxa6hnsmSSd0q4lkwbLYr2v0B75302T9qK
Lv4IoZ4YNAPQvOx2A7yK+r7kASoi54HpEZvF1UF61dUrgJmwufTczoDiqj1HfSys1F8HIR7Papag
wvm11xLVAmtBn2NdCcgpMCiTtp5UgqzbTv8CwkOdNnYw8MCLZ8LC+uzu3l6+IpZ8YuwC6/UGA7ho
fJefV1TOsSgVmzEz1hq5b2lXcbEp6bCyGRhs8O8dLMAutERgrV0uzwLGvQRvS0MIEvD2F413senp
FWERmUZaSwJCHdELtAIC1Fmw7G4ekArQ54IZbehdcY/XriTEFlTeA7e0UicacEEv7Ok9HCF14qB/
SDz2S6E6+x+ILZmCo79eZFZyqtTWKgUvQuWVLspfX9MjFlkvJAyph+bxSvo3F5JGJ8GSw1yUriKa
qmtUBIi5MZ0ZRXgwvVoDEp3dVwHnE1ZGSu2OdJIjefDyYWgUNqEJtYHczOoeZcbCa97GIggj82jx
LvGRefoxYi8cCZOxRY/7VsP3Es2IKyf3r8IqDkCkuvAtPXOAopHnIUPHp3SBx5DyP6MdzH7LPGfk
Y9+qPAJSq9vVoj+o2nj8PAKWG8S3poMUhbqJU+tgmDCBYi4EUVFUU9bMOEqZpBkeuFYLrtQYOfHZ
jMtvBxJ+X98FQZgrGGSQvHLvtuMJXNWSnGTnYGaVoBYFwAB+DAMTb5NFbLhx36GipKiFmTKVFiFv
ij7yZR63rtZTgb9/x66rcL65/N50aiT1cZL2EdVU5zQdtAEG7b224F05V3d6pxR7j0f8OIHt9Hj5
ZICOfAq/8zsSHQHbA4XwxCk0KlM+rk4aSRaTQUGXzUZK3DHTeIhQkMwFrIrzqH5v5xOKGtFiH75u
WoTfVXCdXc4yF/SQYRVumQ+yuqT6S8Qn0QwAqDzQoyn1OffHQyzLGHPO4+IyzGz0LLTYhrltjFRZ
sDZTOSLqHRLAJh9k4kWM7DbaiRxkZga9rxm0sNaqhZXdBqOR2GT8w9GXSGQo/0ioUOQ707rUqoyp
SBv8V4smxBO4EfmCS0FQ/+lABN1skTTRoTyaWRvwRBJ4lrXb2wFQmLexu3zSVmF+bfN2Nv245t1G
ms8qK8Ebiw5T+AfIcUeK5o04nr3m1nrI0ZD61j6DmLThrGF+X1QwN9E0sDSG/Jv6bN/JhdHlmhPL
TAwxV9a92NzuTN3tBJJPhVqpYHQD33u12stslNrKR2oXGyI57o6a5hTOrzGliNuhDETQZ2O1Q3N0
04OAWFlNwEq/BJNH6hRiBWFT1ytuCg2MGjvSujrdwXX6ldhZoFOFlopFuxgleXuk/vzVcKfI54Gm
aFSEoKsnOYftrpsFxPW3waybdlBMBAGjK8lmQZvIugrxqRg4dBATDcwD4DnJ4YyYy808ch1/YWKP
F4RV4cptJG9oG8U695JScwe9SjdzQ83PMWveMV5rIsi3Lt+/x1CraZqhiSMMcNaa5v5SUelEmJzB
f+gZh8gVDwnwZprDr8GnUHbbvi3MIDZRXFQe1oeezN89n+WXx1dPXz9Y//OOxCbQn5b3lTIpHcK5
m7XLAsUnifOqZX/UaiO6JeBUbG2hXEhGR2DN5pyvKCEmEDWNfXL77cNaMy9nn+KvmPnroCQ+eROd
nK2FHNcud3kw5HhCbhkOEE8jMJehOhX5S5LOy+KwlGVaCziISc/AmaRyUh52Lit0htLdFALMyD3H
6AwI/FaD/Y+RYNc4TQUi9YD9TwNVf8e+g4hjkBo7gdsjE4mVaLVloYy/xYMkAvHFxeFkpiKSOv2g
fgHFHiq/r9XS6S0Oo5PocHJPB6F9M4b0RwX8VMVlYrh/5w2L7QzrQojEGSD5ChAgEUg7JVFFEZyA
IdhN3W1XORfovG7OHKkYP2DQnhZSv4f/ezRtOGOg4M3Xi8f7NRzwtwmxqw/5eH545HDdAgxur4e1
H3gwNsmnYoSE0v7yjXKLcIskX24cTMCK1jaC2wIUYcDe+dHv1yHUZPmIlScshbliSQgAQ7ZFP1kh
P9sz5p8fuEA6jMLjTCyvs/eTCgtjQ28mPVpjGsyvABXr4Wdb7Sj3X+BeOVODjb7urv087NNRgkKl
/AglUIgLdbfWETCW3HgAbyVtUOEL55CLkFSwGvrL93LVMkJpDXDtPy/qL2a5ccv8fnNVkxJcLFQH
pMP1GvBZXvUXKiYyUvJ2YGABFkw5hJeO8v9pa+WLoqKm1EPrgrHQN7N7WIvScCcOJ6n8GMszhYnc
OtPhsRTnq5A40N3VyFYJ4xSOdO5t9GO0kE2bQh648sdL+5opjg3fpzF2QCfEWM/iWeel2006S175
B4DJ1RaYcUvMbQXA5JX33B4EZYjkA3cOLQCP2umYDnHDKlFNVUaLkalZzo0rw1/jC2abHjjgniA/
o2tQllejqppCGCqnUC+yUpX9xM6zFTRrOCu+O4AR8uz/6e+gWGq4aRhymCUqRRTwZMBKPF2ef6ps
KcQzWY8NZg0/4vecsBhynVfAQomRJttFy5wt1L9iWntjkF2aB2fBLmIxiyxlvJgGADoJFhHOjCZ5
UixkLcvaffYMmlCgZhdWgaSYpMhyQhdNWg04dms6wVE5tVdPL+SZrVvRX6bchaDY7gYOWY6WAg5b
PUddaCXzCU3QdrJqonsAxRbHtH+wO5BtxhdMSDNYT1MtalUnUS4LtkvgWcMx8DrOvB9/GW6ZBnFx
hJOgvoDtAzIr+JAz5bVgqFit1oroBYQ9D6I2BAlsZAJRW/TP4ThHzVte9UBaR8//gXpJQ0MsZNBo
J10TNrAE0dlsylMI8w/7yZcF4lF0zWdfQ5qMKDzZyZPHAW4z9D8Bs6J3BgOmNlymASK2ME0GWgbN
KBgDiSsSnDGcX4Uwn8vbHliT1cjodmqHOeXQvskslI9Jh59uVVIgEDlvJLSdct1prMdoZJImwdFV
bYPeTXw6umZzP++FNipBfTf7dBv6xf/voHXxXnQHggGwHdL0H3qcEXGV9HV7xaiYF7bdt8lwGpFr
UBwmlzLLdiaUmOwc4MCnFxElBJsYM77Fvu9HoS3djEqoau40HUGKpFZRYmCdxNaKwnbaooSlGc3d
LYhEITyYQJrrOU28jwrXuccREQHbY1xFj7nIvVj5qFiAyv15MnJRequO6ikJ9MMxVeRshbQ4VXQs
+mxVL7WO89Qf61cCyKSEmhemN6yUTmbBTlqEe6i1dUpVSfRQkp5XQgp7SitGleP1xAMu9tx5eutq
JYE3ZFPEnDULbnJLVVQdbkSX5TySuPcEY7zHFke9uEHzX1RNkNUwsODXOIRVLSnTN+Q6waWcuouB
qRQdYaeUDdjPwZumip1PUjNHoV8sRsPRNogDwhb3i0Ppk6u6ZgUHV0Xsn2MwbByra9XDe+n8FIL8
BAVZ7lbl5teAoEm5sEq46y+HI6J/PWncaZXjLC3CwEsYFTytFJOyzDG8LM4pqb4dsnqMvulYSTj1
zElnJ/gfeK6/ygJJy1iLbUlf5amXtcsLxxuqqEm3LOfT7cPsuuTJn1RKidE22diIi7fJ8Q1Kh7WM
CMLfJ9W/QcmnQn5piNrzrbZSRhuyYh/N2SWKbgCYwfqLjYKZnPzerxnXenVojUlUjBuPcmKNOpXr
R0PKS2dQhI8K0pkdUZ97uHFUTl/kuC1o+cnVDrYCmWC4ci/29wC7K/2shHf2grEe6Ci9BpNOHkhy
RhkMAvtzpMXsSsCeinzXahpD/zJ72n9CyE0PsLbd3uRQbqYDsMymb2UabIcHstX+Q+FNfy4HMmX2
T22v7stcyqVOqET9e2t3hy9dqJ8hIEXkyB+CS3a40nFtsZvaBZVJU+2NVFgDFNl2obLkjCOfFwf3
ThYgWjbzC7Gzmug9feKrDZpwoKaWVUgeLTR0hpTPB2k7Fxh7h8vc21GwCsUfjtGaedmNw2q8nX/l
x4c7BJlRhUKjnrLruWZa7MfYDmHNnvxpaXJQ1zgAPbmGcrp1p09y52hDu6fdLeWpf89e3kgpYiXA
FN1RqWVsPkkSGI1dQmIKGLBw82hddwLjYLlCw6FV1mXch6Ys0fQ9TS7Hlf8wxUVJnr4negvFhSAe
K4PfewhAZH22i4PLYx6KFTwYTSO2oUHlLZut9ztSYcRvGY4ov80GJIxdVHN6il61Yd5SLk4O1KbY
vr+rqO0e95q+NKF4HVEB57UTMd1hZhUFuNQnyLf+cCdqObp1yJ0z/fg1hAA07qcPIxZxEI8Vuabw
5am43TKqPcdQq9xJ2nC3rAb7dWYdAH+UO930Hymcb2AONiY/dC8Giv4iy6Wcuzr/BTxwYOG4Y56S
pSEIUDA1tKsiEl7UwOP+E1oH2o8SCrJNB2u5ts3meVZoySpl9dGpwlZ3Jjy+lmpGYGero+VVlXhX
qftNlDxWhqE6jAXC14swVGq8ehq1SknQubxjYkimZACDeLSG6FmdZ3S6rR0smuLVkHgMtW+ZqC/N
WXxL6hmWWqZ2jJtuaioK5rEL5w89EUAdZMU8GHafR0ym/43CizsLUMd+1yWwsxgcaBAdU6uzQ+jv
WULDxEAOQwh+oLTJKDzly9+qd7iSKeGRsDl4XT1FKKrL2KAhGf/qUeiLrIoRpfol+pOMoB6ErmYt
u1cVaIRI3159T8cyJZxs273XiukqRRAMyL5nvLsjftyiq/Ioefntlx7Ll37QBNI2MsIq/vQu/Mj3
04z5EtPi3xI6C2+QXqJXBf2w7GD2viJqQ8UTd0tsK0A2bHtfxoeErRUe4xtADBNuQx/jG26rDeg3
AkAv+agSwKZyUTtF6DcCyzegLiPeWizbRygDocMT/iPl6T0OWhUhm4pVcnqbfX8cz3Le6/WEeaqB
TitzKbYNDSnUUxfcwMhpTbYKmLjOLgwpqimi0OwHV0v+EABr1v26otFyrlqQdl32b5sWJlYslv+S
wPAAUpU5muF8CkFWV7wWsvFIwHyD7pKR8W7trEiJKRVzzvQd8eHLm9WnU/ctO8LERpDHKdjgR4LD
odcysOdxDR3cFYKtRTYLKFMzvXSqajzpcIoMF3jeHewY9aDIaLnSE0mQ0z99koMMzPRHMlRD6hDm
h5etFYPK2BrWjY3geTyIBCrNmBV5rby6Bv8DISoCeIHSlPoK1hWGXaotoEypStP6sfKHfFc9DsQW
Bi8G7vglOjQ3dF9wrWLqgbNf5eFGjzs3p7jxqknPEtljepIMLYLdLY/Lfmj+9xhTMyK5dXuSp+/j
y3GFRGj4YOF3v7zGY0vbYc4YH4WHNKyTnzrv63PfwmyD2FOYEqzpvUmTICWb4eG4bzkj4A3MKWlE
Xep0ZqGpbfwzOdDLtxsqVdC8SC2KjmehZ/EBw3KWFtG9nNMs8SK7dkW6ys6xgcEI+PPI0uYFDH51
I3bNCGz9iEC39JVNFWyDXpHgBEhh8ghh1buGbIxsagVSj4OsUHSz7mciaPvm6iNedvzya++J2bKb
8jYxKAFMjeBkgyuqyogGMDUvGcRfJ3f0zz83wtWDfcD8h6zaDMxQXLkos7brgwA3eKz9DmmlCbp0
vzmgyJQ9waWEC5jj2AQL2YvE1ZT+ej0CUt2SFpb31Zmzjmm4adqbgu0xj8LWrgCEJXr0Lm+J9BVS
DMdm0OrQbApDPFtjsD5yuq2oWMOc7x+FrbXn42sAaMcw3FhZf4UmLZJfKzQCh05YHBs13m4gqceQ
c4ELw2kCtGyFGRdFgS+s8AVkAR2Q4Chk4XE0k8+7R1kVt3fZoWlqnsuzGwnUSRApvJB7eXnQFdmu
tYd8RyzxqURuwd+aBKfYEZ1MbYxyw/ovQdMUNZrfMmBt8a09YJuRVfNrYtV9H2hwmMKmQBshJJNm
ofA6wDmAZ5X4diUWszAGciYg8S10PAMSDekGvSpIWEuqCCiXlSfCgjJ+XNiXnqKvrabKSGbylkZM
0TT1LbbS5PHm3JguzDs6t6yOpNWht2Qjqd8SKvcpH7sxS9kM3KuPzZw4RedeXVS/bEKItrKY7h1G
XPx0q2J7CjtWwad9286Ulj3rjB7fmtf23sFf/bXPPmP1eozMwoegiR40krXtZaBmPExFicvZaJmt
kG9rICSK0wU874j2JTI/4r2+PpzlY6bE0iz9KYHJ8JuW1gABiHc4/8UrfoTXhvLnNMqcejodjAas
G+c8CRgXQ4Xy7Gt4TRdFlXWGMKBi0U/giDEO79xjw5f9Tn81r2EQDHEmp9/djbZJ6gfgzUGgymrU
GmuwdLC94soUfsTqa1KqnHJlLxHQpsdmXStGi3gkGbiD9Bbbg625HfLxQJnD6Tf8bZKZNO5hhRaE
M1uyRW+WLmqOZ3jNcakhW/nuERKflY7wETMTAQhFrD1aVh2c8gMxrp3NC8bkie3rULB/38xVxA42
MI9i8uHmmBcyNWZxwABFRY0KhBapv+gvXTa7qsM50pKh8FrJcl+aXCV10K9XjpigBF7SSdA9AynA
kAWG8s6ARDyDeeqnnECESKo/9UZ4MJdD3Y0iIaZWSA8SS/RxRMcUcx3pDrklfHPKRW2cXUqkmetR
3fAr2O5fopcgLrRZ3cYqystye6LYV1hjADyP0hCJwC0P7trdpd4u1AVqF1N4KA3yDaZmqR7rZqS7
wH1QLwt8p/jxVPr7Wpkoe169U6ssfZ4BgsFp54fAb+qerq+E4QkJvgIs7yB6wK4UUXvM6lmZSGVz
hmUogkeM3DlFEIo053SOkNGcG2FnSgTgVqxD2gmIo18fFUalNMCRt0ohIdPxCqurZQlWii9zdDVB
n/SOf0R4EA7Sx0W8vsPmhswmO7hNkKb/tNjA5ZS/DkE72IPO8PQX0BKbsEmXVf0nNYp0IfwnXvtx
ut2/D28u79HI0heyrz1tHxEcTqKQzJ+V/fmHKpx7hmV+mNLdyUGEtNP9Zc69OhSAnlL5dBozNWTb
CkdiFl2BwyekWTFP80dBSRY/+GQYpm9nUXBZ+zWhSLQkj8+3rNk4wsy3lkmRxKE8oOgzOueZusdS
CQCx283Pa8SsIt01L5DMx2k1/n3R6nc+vQsACIMjIxWBdV2vkFUyontPLfCrF72+E/cKRckGaNfB
JI3WfxvNN4Jsd5us+k0hndMd1H8VRH8vofxc7GdWyu03kxuFaCqVumNf58mz/XWkCizEwv3pbNVT
2IWdxyE7GYcB+uaWpYzN1I14ismlH/tPt3rE3smkb/RTbNSNpNhbJEzjRn3PbWLE4pB/aKe2CsON
46suuxL0vKSSCBmt0qP2qGVN2BS1s3eumb+Cgj/bA7SiIS0ghzLDsbzhmX4JEBh67vXsLgRJAQqp
IkeyiHLQ1/gwbPRlm8iEeBd4hbLd3h0GooAYh02aklVBtTubyXcMqKyX0mM3dLneFr13WU43Phmg
YEms42MG2ERwu7inytM+BhlplVehCq3k7i/kFvPdyPklAiFBMTdmZFkB/ihirQube04XFRvGla8V
DEYcvYA+k1y7e2d4UhrlPW0akXTV4SOJHgjKuEwmzGkFpCGMnEZJbFV3dVoborc84AYtBNEpgydD
tNQ7IT/99qRB3gnRfH58Z57Ky3R8U2Zn7PcESIWcWmHOlb4LjA7vVSmTIBX0qEjQ96FWCXqZs5i+
Cs3w9It5/gNY9q35RyE/HNsthiFBJQYliV+85WlZohwu70Q8NSAkMD3z4cs4NRerjrNNtF6iof9c
S/AooX9IhXYRTBMm76B1n1x2bljcEVR1bwEJmClj5ZqUbebJx4uNvs9uuZI3nQnv3VtkQG1pHDmS
UgktcNS+lejF+gF182e1wcmgLOqbz6YhuAgK36UL9dCyMTJUWdLYmMyFmTw/1AQ6ysytfanxKA5n
S7xowMJALs15xoAFY+stg2uL+UXQKRrrYeC2Gu62iLoNW0+sLPmwfAAPtLRSwjEijGgox8EeUZvz
g5FrXwxTS6bQwJMcxw2836Va+ELTf6QWi0Gx9C5uirxgql6iphYmQxEw4CaAXYXr3YoxKKGoiDMs
Ko/cKe1pdpjHHJLtj1UloofssXFAjOTHU9lsW9jinC7c9SZuipnfHkXA5jGyXbRGbAcRhZWWfZAW
86eH6PElPfryp4ySQqv2z1aThtXdZExN32AEeBF01SsLU0pcBgOI6x4E7QoF1bJRu3DD1QtH6AGz
+VjDL5ZqY0CdYqeUyfKdiVv1dpsGlxuWP20eYJY9Irg/MfEvs3zSrA2yKF4jCqcT2EjG70DsvQc/
0KDWhqLAg2DnR5tDsGfxb/7UnATFWq+ueJHXyam4TAXRnRb7BzlmO6H154IH1FcZ/SZ78eQ3Xnmv
6R6f/4hJW/cyEwnlxLCFx2KBQxBKhK6VIWIENiXbUfkdDcRFFK3M+4lt2RrFi8FtfmRqZ85ExsD9
eR+n760Q2tk+9ylrdsQhF/kIAgNgKVL0id5fchEnGzqeno/dSpI9fP0vGu+aduVvvfWh0zDIJicd
OdE9AWTQ1hTHSAtHUEo0BHdTrttE1FW1pNyOJhXDr39kfjTgjRguHxioNFUUMmlxK0aa/LW5Asgm
13psGCMquC0Q3bbbEMX2qemRB1hzvmMByMjcu1h5F1ZjuGpoFuHPMV9JT0r4kJLKKWaFO4cvHHVz
vnJrLy9NZHpI1/HvPUGu0oW0/C408N1y208H8mNg0uxOX3Zg9r/1Um20bmZDhkrrBVbdgXLnzlKL
49Yqa8krphvQZQLrih40VHBjgvPxMCvtw8EIR0hzVNLymBHtwhKYzq5ul4og47gfiiIpvlBZmPsj
WQgtf3w93HiItj/mxbIaJs2egZT4WSJn9wqnayLvrG38fpVs5WFesSvx4oeoYeEPqzKoQcdpmd2j
IjoMgHsRz71R9CEBh6KX5zZgccxH7GrhlrhGKEDBUj9tYdK4fvuf8cnXYY7eCJdbG91RF9+jOHfc
mxvAqwigIwO+GSwgBC2rAQ27M7Z9T2TT24MBXEDql6lfx3HeBWFd+yaht5PuaqtY/VxjLi7AmkOK
vJPuJcmX3wTXF5+WGooKK4fO+UenDmEvIDuGTUDxVbWgzwG6XPHZ9A++NoB/xSlpTS4YQ9qqF69k
8oboNnb2Uv30xSOi5Z1htmvF7u6diI24DND92GwQ/wkwH6/QlGGH/dsuyZ+yEf5uboEXOI5s6mf0
EYnoeK0rcVxZqK5B5CHbxbLoQD3j+s9iVMQ+sCaQKZg2i2WG2kCbQif0rRw7pmRDfk3HjyhTL63h
fZMjRjgysflFYFoYJUDUk/SCe91Oq1FQhgat6Hk+nSzOGCrAwT+k+ksF/l/faeS02SrE6f6Kn8GA
ACSQij5gpi7mPH05CZmpl9Esn9r6CNd2qrlO8AsyIOjXKH3fzamNj+JGllIY7cIstsFHRzI7bVXB
8MS/Ng4U+Z0rlSn7dwqgAGpBQ3FeXps6jmtSlUsZD5YlgTySd9RDPnTFl2Des9PL2gw7e7gm4cKH
yCH94a1rCo25HVLIAUJZepEmy+qkAQWp13hXbtypofv0+//5whTM0jSKqNaSjIY7xmqI9YACoq9J
g3GU17IPjXUx9sPeCPqDpZ7Ap9zqzLW/B2FUif75Kph277lBg8EJiGLUYq9uaigjNK6FyHmepfx0
c2Aqox2vZVnXCp4R0n+gQm2gl9rfolQstLq6uYaiNdm6EFg6uM6Yf2E76gSLzddBpzqavIzIx0bH
owKD0bwsukNMIE6NoQDPcWHjahBz9VpKCz8SrvXNqqhBMBlRlwCiLjs9pWgc4NUKqMbJzf15Upug
9l3Hp754Xn2Rw9U6qm4eQK2AHLzKIzw4ZWRFhzm+6EkZ3NHRV4yxE4y+YFb2xHpFiDNjmhyZZz/d
YIoSFiRNNXfTjrPKIRro2OAXUAuqzj8vwRR3NcV3UXsLmkc7i+FIig11whQqSZy1rG44zBRqvRKb
90pjozNLolC5F9yBlZVCERT3KGi5WgPYjbk41o9FhQMS/khe8QtR9qQ5VyTGqv7zgdzGrwJoJI4+
p6H8/8wWX3XuVpGwSwgzlKRAfr6c6lBpL3uQE8BeDIGuDvAFFZY14jU1lgUUEzvBt1EGe0dcasEX
AnYazwbEdH5wpZLHx7IMhV1JuEdDlUxs/E7SBu0aixEi709OZSZ/gWaRM8VSHL13znf9hxjNORxX
UFc+S1I2IecgceaTa9zOLz7QLBEJ4Acgk4XX3Vw8iYapsftrjd1ADPMXZoK74ePiGyLlXszsrsKS
AGYe3+GV4/Fji3Ls+m5nvh9K/mGtDKQ04HO/scz09Xzto9b4TnQlqsZuEQLp9+3KfxP1CObsxhCK
nxB3KxQBkVCs6J02Xd4mZm7XEYvO7Smj4t7t0rioRXg/uHzrjfQY4KQEK4V9TsU3IHSGNvbx73C8
pz3OMIjJ3LZyOEnI2RZY84j19HY2yUJ6Jh9FsgZXfJ2O/VT1bS9+HOm4wyqihhw6eHVVjx/eWGkV
Oz7iiiT9+G9BZQ1w/07gE2Fh4nYQ+havlHCNJ+YwGzFyZujpvw31W2UXNVD+faPA3KBgxehgEmgw
3IrM1OmXtvG/671WBiIXhqoHS4SKmi6WcWwrcfVtoQKt0nOccR1NQqwWzyTOOgn3elf8FVsDJMOq
FTNo17ty5cnJIwsf5M2X0/KGlHTjm5FCMRwz190WqTWLfk3hauzElxx89txfNYsQNoVOghev8iyA
62wkHfUsCU4Uvf8DuB2v2/XU5maueEWsZnikBXk+lVEw2W1NbcO0cbJAt0ZITnc/NlOrmJA5CqAm
qXJKpPPA+qGMrFjUw2/OZ/iKMuRdgAkAHHQ41AYvwPEbx8lST58mWZ4xLlZfZSjkUDMp6CklA7pr
WCKRFidNLBmioHuiyomFqxinZpY/7kGRpsiX1YZW7DJyCmSbCw209DlirGOnlEbpQ51/43B7PQZY
5aV2kxMouxNvj4zANMW4cK9XP7rJ/Ay4plIZJG4SVQna3Oav3rU1JtOX5e5n7r4B51PpjEeo/NX+
FVCtajk+A+H/7wL1jkm0ps3xfCzWpDR1ltmP4NQqjqzx9PcV6bjLaepjdj3ZdveiMLkKWcXkG2Lv
L5CN91ISDGlxt7bj5cCE/O0BmLZIXiqlLL/SUt5wvNSIGjBkPUgyUGBtxJUVbWavlkLwM+4zoc6S
IoYaKu/hJ3MxT9s3e6MVkT2Ik+0HkxZYpIuowRqimvg2CgJs/vt/G/ofaijsXqbs/CCC0czlYPbp
hD8SExtion+7/2eZcPm/iYzCNOtB4yHb5HeKL5PFZe/m0+YQlL4v0Q9bqO6A9xk0gAC1sa4u7znw
vpfTTFG4hdd5vDp8xuvqdPq7G2+Kq09Vr+6BXr+U/O6ltgLupVtBAh6iBVItlJhJxRG1hCuARIfE
1wIh4czXJ39h0zyw0TtVaObbk+3yW8bZlWw+ml0M1XZxFMw/Qg9VYUdrxLU6a22DGLvaXtdHbQNH
n8OFq8bukeVARlSAhFxcj1FknaLHvNzDzlCoqOFunfQ17+nraku3/UD/6U26WcixjWyczPhsMkgm
hMhDufc1nKTKnaGNVzeKTST/xclCse1r/EqtassQ/d405g4pUxS3hJuKLgdWjyI8hU5giMWKn/VX
vs/sau1235qQ7TCzPwxQ8ut1WZRszADw9Q7uISLGbbdoFxi0jQyu/RX8gy5reF0yJZEYt+e/rN1e
hXqPYCqBtqgBjGDuy3g+hEO5q9a6pUc2Oxhpn3S/3MblQsh9FHKI7xJG1OBgKKEiv71r8xKmbOXW
tR/PJj15xupTfjEYBATY29BO+f4HH8AWeAF91yepwzO20UJzoglwhbT3L7sq9cBE7lRXO8wYpPl+
SSQ+apB9mRDoFVyf+h3NelT5UA9M/UmquUaCQ5xAuw2miW5H4uVsONyIdrFitIzkvef8WnVwIB4c
nhSxOHH0nU4HtgQ76As9gRLGyeCxbSbK3aIAKpoNKY7BpDzfHuzsl/0APEzZoRU9SkNDhErUonNJ
RU6wTfCgx+jwynzPuAcNjJSAVN4WPOqQ9moDLvHSq71TvsxBIpR2XWXpmTH036gsckxh9mhLNAgd
zTGzFclq6YSB3E+j0jsQf2mDcYGFKIugg4WkcMxHVHWGQ35RJjMdkedpnS1g0wSDRGwJQV206Mh4
6uG517+ah4YD1lnOuRLtMyzFek/mpHQvBMUoXtSlHDxnA+HhkgyuawgbZIuJeas+BrPCslQA1p+U
S+Zyqu+2YLrYgGucdB5kKlT/aGe40I3oOUGZGy85FOM6ziHDeO10qVg23yrkgQ2iPDE5mTM/WSce
6XZ1hLg5LFdgouD2gX/F72I7RqYzK/yHIKsK9syacX/cedp3ZCw3To9ojwVRxg7fd4SJRQDai/ZG
KAg3yIv2S3XXSHDjNGG1KpVS0SBjRPu4uy6oW1Oq6xRe14EI9VzCq5iFrNl2ahG4T9b0G9EB+BeZ
0jc6WO7OWnvDWDLcao9Jjxq6RRcSZuB5f3MqPgQQ2wmIvrVpBxO0xJFausVKsl7W2VSuablbuOPH
9H/kXVGPGRRix9ZYyHcb1+LHB+pPFwMW2r9WBmGnwOhg9rgKK3MLl/0SBkHl2K/bo8eTt/qVklNv
diuZkyV/srpA0bv5OwiSlri8Kl6KNdJGXSVT5L/l/jzlpjSazNXkL1eMsH5N5fsuQ5/w2Er2Vacr
NjrQVNwbF6Pw/oowqxIC0qHTj0txbU34p3dfGuN1a6dSZamzL4qTO5swqfkkrqyGZ8IVdeNjDD+4
ZgzOGjeINPnqrg++SLWY1rfjUIhEk63VLDj4txzJUsIMBimT4AyKWe8Klf4OQaqSEKMyRsRKd1jd
e5xvNPkBzV4j+HUf9V6uBcsiCmM3Ck3a2W8a4Fe+EkVua6n6g+qNE/R6DeblGL2uJ86V8CWrLD8I
e6NgWZ+VCmJaLePPmrhC5wR9MvrQYXNcOIVWp9zEGpOcORxZ7vJEDjoTKZFuOkXr9Xp3nupIg3J4
ZQhvReV/FsS7Zfdsso8kTL4o6h2HG7QieiZBLkU2QB4iihouIW/PfiwMdYahLAuisHM0+SbbG5Bc
AsGR1po8Iqmq5TFs50X8n/oAk9726hGFAyIkzcoKw21YobDykwxSqRdWZv7nd0UG1HF5Ab49XgrA
EUeHVBUsNXF/q1QI+pIqsl9jfd1cMvnJleQt42UZwffHrCxCcqDU80pSPea4r4fHH1ElF6FnKo/Y
TiWulBIFfx7aDNoQQ0gjYCG4E1LVGgeKHFlRZOVPGV/jHf46iPkfKXOOpM+j3xHyPNzhbSJrEaA+
bCQA8329Fsv6KD5O+B+wEwCsJ1/Rp4CDi376dKzNVzz1aZdBntdGjOEDTJnSsFbuw9+BT/+2Pho/
pgyX2ErMJ/GeTDW69nNmwxbgf9qVQ8Hn1HR/Pk+r7AYkNDg9bxNVG7wG0mo3cCQ5+aIB0FDzd70U
s8VkRyNFnAMqI1Pxj7SfAIrQ51nlb9L6yh84Q4oyQgYNffZLjR7ppcNmWG+obvJNHhh4WQ425fmC
vA2cRz1X7/0NY+Vmvh2gfnyJkZKJj7D/Rqwq0OFsV0YBMZr6bDz1sHIDRbA22NQYBuUhgQNVj4vw
U+VnijydHgSGbNmj8Z8NFtmwVIGkihthDBHMfSqLDrRq4mboWjxDqGg6kDgIBxXL7qjBBQlsjCyF
uYIiKz5fCADHe7gSBNwzQN80SYxNkVEYVD7/DTCJmaWz5vZHD8YffmHTFPRjPrKYz1jdya96qNli
lwooGSl+alqojfBNdOdfpxouFtFSRLsqfP9/eQPhhNTzBIRa23toVBzphh5WgZ0SlrRRrb+CQ0gv
aVuHahtOdsOKIGKX/Q1yPMUegdjrTXfvBXNgY/HR+uFC8voJKADPbLIuAo3uJMAJXm7mr2eWvBUF
onPKoBKen9sWsaBBzKvqeo9gWwVNY2vU0lj7JQsZ2mwlgIxvCZpCab57iBb83Al8CXP2iHAhBskF
gx+Kl4kEijzgBkPvC9R6+VGAcGM579mAY3DnHCrhK022XDUrdsH6/+WVkJ5jObSRj5ToexqLivpE
sxLK1BKLuYU1XCrbipCVZNxbs8uoCZLQzMy/6Vq3+P1lYujbYTU4CH6vO2vDssVNjkg2egUVMROE
YGVBZcZedZSrjYo/nplPl0xXC86HI1O2L/RIRrBRlXQKpun89t/YNwPHI4uMdC0BGcqX8BlMZEBk
qABIvxOqJ8Sg8DAiyb1opU5bYj9Kww3Fm7ot4JA9lIpGGLF57uSMuUE3NL+q4vfX4tPmRVaiGDj6
1Mw6durmo52+YZuuZh9hU8cjwMupgEf59FgWitMHedmRD5SU5VV4sXAefT/xHvr5EgcRIPJDQuwv
nbw0h4ZXwVNp3GWOEgiH29uGzzPMWg5jzSsMZiXf+ncRY97CdnWer7JZk7KRvyj8XwQ6shrosTqa
F8IHgjFP0meYhclPShz7wujxRV88TGKwoixJmSSCEwZf7+QjjiiogTHS+3MokEbotEHmnBVCb5YH
f2dJ9MFHycCcQieiPLW7KEjpMfL9XGvszqBXHD020kqH3nAjptAXsBT4U+d/DgjdQwH8a+PlxTia
7pnMp4v9eiFXj8jd7cb4CcrCEw3g91UvigE1FGYlcCh4TSXe2hqBc5Oc3hJoKAfeXQhMyD18U/1R
R1WUIXVv2mgNQvjZPQ/A3LiciRu1kRXUqPamsNn/mC+tC0PgZznxWvtrHLRU7cqTIOGCHP+cTJF+
ApAk5Hyhh6qig8iUHirmMRnpxyVhbu/IsPAtKEZePqUWPEKIZaI93U7KyFNyt4ilXtPQwg3JqMgR
MyGm+eXCk35fywNuy1eLzkS7r8jSxgFW1BYjHMx7KYq84GhKNd5v+rVOpwRvqa8+jn8DLVs/RePd
vDMuCnBGrQabTAGa3JDmmnM6IDCGUZdwS5bSqRZ4r4iyNHfQk8vfJP0dMnvrsqCUAI7y9xgObokr
I1KtDH0QuVH72xqobeKlHu4m7QiOGSI7a7ezGeuQt2Azaenfl/55ugL5dp+TAmVOJzGZ2Ng5xDW6
Sqsaqu1Y1Iq2rsHelalLjpSpaFbLszXApSCLIWhngR3p6oDY2Zz7mQjtKBubWQwlIfYWiOUvfRoc
yxy7ge5j1MdQQHynqdTdMCd/DNidR7kyKLEsAu88Lzu2vg2rEVYUb/srqYR75qF5Kvm8yT2IjXS+
b49QLopevyY5lgaXtdz0rcaU9hlVnOmaNqrV7g1vwG61WGfgyQlJTGGoJ3o/zvx6cGmkZS5srK2C
BrCud/0DL8H7ioDvRR0EeMojDZY2CMwRK/aCU9ACDkTUatsaSZTrE+mS8XlUqi64SZ02xXBpWh2f
nOo7kHP1IywyCbSArYGw4pdwc+0ANWjZrBVqo72yPXlPZzPa743H0d4MCrFy4ZFZjaM2DOxFGtFA
kMEEjwA54ZUdfzXGrSAAIm/rfNt7P0Oj00Z/gALCTDyIUTLVqJTceEYSSgeeEyUTrVOV2cyN+UyP
0pQlfGMaJP+iKgJ7/+jLTH4Lit17YGVOgA/yx5tF2bFmReJ0fh/sOiM9WBMYjeOQauC+9ClIW0ai
aI8Clqp0ENMLYGQAD7Iiyku0W04uJr8Kb/Gl3ecOooWeSGdlVJtHjq2Q9WuuxAJy+cJtxfKw7eJ1
/8JtYBNLbvolFazpmBgvaAcmxKwqMIuprB30TDDfMjfPK6W6RKyo7YjR5B+BtDX8iltP6WPKmrEd
Oqs44p9jw4TffoFuiX7y9ZqfMiaqGIcyKnJCNBWN8aTWPQWG6/j8r/og+6ET/r2UoEhwtMgpuKAa
7DaN6BnvAJ82PYqnYSL3uRV6sg+ow+0z7sfhhGlQpPxkS+3mcJIJBa7HCdhJLv1guvbKspLyI5/j
jg6H4SpQCmt2LNoUJFXVt3gjB7YrFJ+xscvE34W8W4LV+T5/8JjEd8yLF6niHdtCU7Qw/NeY10K2
JMbMvjL85xDWjLifWB/tMQPnMW8FG8uaOACwhIDRH8jZMzh5V454w87ipfqcgLQItTYRZme2jjlV
60+HUAyZ8TLQKiKFm1qt25a/PFgDKSQVt9+zmAit/mXN3xwRTYT3yE9c1RjFpO6tnZAiSWEImtvy
iuyPiTjM3O9J8mxhng1TMyXRWs+YGgFalBSt8UcS54YeDukVa2Msjy0nL/LJ9gIbosAR3zMm1kvJ
P4mXD3RBby9iHOyU2IS/OFagUYlmN2oIPuJU1OP1Ysr0ELVdOFIY5jFXwOkR4msDnbLQqigl+6Tx
mcJ/GnuoGCavNcOpuBjFQIyJ0v3lfJnyVq+7/fFxfsQ843yDjP+P//U7Z4Ki5gG/7JXDBWJlJJ6W
PXSqDrfMkBiYmnkwvpIWnQWyjElnqd9nnlei5zQ+0vITkIMG5GkMmeZIMGdmErjJAi04s2K7ggY+
M9KEysontHpIpPUCP33NpuHbHQZI0361VAuvXhOabYTk5GrIqgpu2qz4Npy1ROoDfHlVuGlvBoP7
+OrBFt1e0w2Ph+DKrq3Wa9N5XD9DycQixDtWtO7vkjUWAZB0Nm9CRSe53cZViwtaroBCN+9wFQna
26HiZ01vuQ2Qin8ctNsPVPGP9/VedEYNnz5XiWfK74KGHBzacxFEa3505mhZUQoAdVbmwxv3r6xc
HFTWZXbfFlpIwk0a2tab01BdeS8s/b7LHSKNDSHZCeXanoSLEZTRwqi/QY18qPAkqI/PT6lDfmxj
UIQykTHC0ZyF4f2oZBB6OfBk99uxdPLhNgs4Pt6GBB00zy9GJ5zq131Y9+UD+CUaJlSVuHLbK4qN
TA1yExAD3iEGzna+8chBXxDM7A62oe+Vy4869fVDOzZQdELfEm3Wcz2NuyoiAcAtpYSXa+sED2CW
rMrchvY6lt1H8Am01H/2UFC2tq+c6u/THXuC4+iTLbCtBO8zjxAG0MHo4NUBZg3kQC839smJ6H+3
J2LaevAVuB1cmWwxi9AyV8ljA1e+m1XhobIz/UYajRyTHK/tmPHUiYlBzAB3LQWkb0k9bkNLKP22
4czJ04V8QVY7RH6riFJWLz/vyoISRjBdK+EuVmUxst8wIDdifzgy+hfcPSOGMy9zW6atXuC3nmqk
AooH6lKuFP9qvOq6HJol3zE9afiAK0ryo8FjsKSIk7qfoRnYL3jpJRcpnpqccDxCvI7nmNqU2kXU
qs+srsT2LHQmbGMF5fGVPoEaX+Sb9iqW5aJHE6w3LN6Oc7R1ygPgrk+nf64aYW9NcKT5gJUK1o5i
zP9qubmhh2aIbKPiwLfAuMq7dGSKXdAHuDaEs0hY+C7H0iphvmNsDeM2phstjsyQALS6+RKMc2nB
JAzRK3uEs6dk0tz7XEeHjG4/8MxxTXsdH1XmJUC8qfjYPSjALwQDd0/eDy+mA4dL1L8l7Bl1BeMg
9S+UHRFMbasd8ZW76tiGwVLxyxUZcTQgjInvlpxwMYHVYKbm1zcRddI/T25IKq42VHV1QHpWYaqg
ykiaSKecuzZwdUnXCUz7wbC0WaO6jzNUqw+z9btZ0WXdXYoWjSJ+0y/93r4wQkUf7C3o6Bhtht/8
GQQ1dXMvu9S/2YOHOllTYOQuEXEmL5mBEgMFYRei4CqeIRln+TwYWDk3vZ6WHvQsawgtZb2xczob
w/b4eOYE0kBk6Mwvjf+iyACtGk4JDRZowu3gOYPZM/JRraUX8V9G+5KJVToZeenqpNGsqB2T7Zik
iXzkQjhmo88kgLX7cm0o45krRwl5XIDQgnUqb+CoiwAoUBlId17KeJvNabz1GKGOZgE6q6xMfZ20
miBFCIYyb4WS8SiE2BOMiOQ9mzCTM037o40Z0ULff8vLGyjusGHFubxRm/xluVSwAjNYTji4gkbk
zjroVMSIzcIMrvpacCjPwWlB34KMQu8Q2WSAubHtpWt0z9hDO99TH3jRDgV21tc15E0GLyRaH84+
ZObJv5khMLXs7jufzczsNWMmyqqtdaXQS+GGnTNzZwuUGkvDVuKPBZbG1akWtA+bqV+QOMF0sux8
+WSiRqwvHpuSpmGLXHv8w8eSy1Gcy9gESpjh51TRTnuIPfQOHRKqw+EqtYC1kpvY/FtQlEvVWK/g
AcVdrN8nCPcDChH2JyvWsgoucF6Cjrff7NWr/cqZqgqpeAa7ZKgMsfGJAZrvw1D8VmOtdNXHOzZj
dJmvdmVzetR2T/bSuMuTf+SnX9fMnV35wot8aAC/sHgOCwviT6Hhg9XVlq2p7ZOBv4pOJB3RcXND
xzqz8iw9eHZvuS7+U8gKdKiwkLJv6Dqh75M2a08hhwBny4vg4QSblCYk2FhVsZvOWRtV+ihla9mP
NzLiBgmZv49FUggk9BnaeNACFF0u0aKp4m3V1s5xVDum6lci4cS1h74GtTPoFhStyI/3wFVWD7sX
guuVD29uK21D6Wsw3JG1muPYEdiQYDIXGQRd/WO5mth2fDeUATc6DsJ9UVIkTCet7WSIMEilOsA4
Zg3MHMXpaYaZHzk8LYVyAk+9hZIMgK8ZyxwK0Ptht6w4VQKBmT/5YxzQco34wC/VkCr4kjfwEetR
1+mbgI59SltFHZom7I3sj0zs3OCA9h05su/PMSlr1kBVbNxZ5oKNu0RNgdRA5OQVy6DTR6SJQzDY
YcBUf7ssrZT/PJ8Tig8uuzQD2q7lGmKJcifiFgGyan8hf80EbDTDI410ZmGg2VsqAm6+Qe2QP7Z2
fKbd8qkGdeG3Z8nyx8Kc6As9tA2lo5dWYCDpMpcwE9/5Kq03idT0xd9Ar/OlKDQ9iIV4vnNCXC/G
psn1zIYNIAgchZKqjsTzux/rH6sL9TM5S6+JNUPYaBAefqvmZmPQFdlwZwmmWpmWimo7Cc5qy7VS
OV+ngTzuIZ87KrMvDqaXZgVMjiBAmyYJoWyY+ysJWGNIe40MxhbciBxCti6Stc/Kw6EpwgVhBA9M
KafuFBJ6g6j7hCD66a8Q9YRMDMFugIZ/s6pY1JEHaykE9rF/2sUwRqZ27BfnLvuJzVhb5j74Flcm
MkInOlo7Iy6GrjlhINGgpUQg6KkLZcoJDUkWt7YoufPLr6T7TBplyypUmUtIgXQ+Aura7W11sV5r
N+dafAhGErQ94NkHG6oGsXg0kYv++QCo6GXEWgTtpkGgTpD03K6JYCz5ifAncC0dMfK9vH1qKiHD
zTWpLa5DT03MBRb4qRyvyJE2UNfejLNlb8X3xi1WNe9LVGKBLN4lEYMfl+rrJXcfMYES588TwF8U
Sz/CtDoyQQ3ONUXXcFoWDlotScHMvwtbaEoN/JO4rxyzp80OG6lqmLvi4uJrTpSujsCSJU3aZh9w
RuS6N0utWybVqXeLqFzp0HwcrTx3cRc+0oh8vZuTqFDHfCkHSOasUTJLoWJUpai+Q/BaSHJIno/A
3d8sE8n+05hM/2p3kIetOjXroFyZ8SFMTrjxYCvinUoMz/KkjrYzenFKzgJ9idOgvRyzUY/0/0YL
Wz5SBLexhrApNU4Q+EszC7omJT/f+SoTN0XjWVgPvQ3fjGb9sx2KcFhg9V1+F3Zysh37uYXj+IgJ
pAU4V0lZw2HYtELKvfsVNkagxgYGvST15OsegSY+ye5oErvXV7PWQQdrnoFEW0I462S5QqbZJTcA
WRM4jiO/M7GY6+/rtjgogfZ2AhPFklYSiP/dkIBIQR9nuBTsIOFXToUHiomvwZdwJQd21P6+mQI6
05foROug3/qggN9Kr3KdtF9nrygevTr2FrwDJwN04OAWxFfVb6zU/UCv836uqusYDo+hboPuFuSq
RxgVDsq4Ix6NAcyxfVtS2b1S4OdN6yREdlNLf/S4fWYtF+BZ9YMrCEzNXWNu0Tg9yFkAdDrqiBpP
QEvwyl10XnBqjaIXEtyKvhCLmpmm7HHaWCwuPVb5d6nScCmHI4J4hJO8iLZqAViQD4dHpdxssNOn
2E0cynfFGRXqvm+xHvZvOfGgPFmRATw3z+DU+DohcRjOj83qw/dgOGTiKv2/7pIU0PGl8TSTwTVn
OG6+04lr3+9khDr1UiHDWPY7YFAEQJAJjbfuBQ4KKAn5jE/ECdrbqwx4VGDBki7mpLW/Y1/rWACO
erVRDWwlht90XeKhaXuQxlfA46iG9miIY9iIPNgBTqnV9njhsCcrm3dXeGUubpUun9Q4V1WUs/Yd
ep3LKml2zeipp6VstTlPvqCAf7zsAqr+lHMFOjA14BaWQtDETPh6a9zMmbXwUNdLAe2TlpnGLamN
hadP65XroLYH+g8WV7yB/G6zscsTzIXGM8NfGfU2SHn1XaiwfuCAJjnmBuaK1MlP7t/y/mOFYaFx
yaxHWBJnJBbeNUfZREcp0KaNwsN8LKFb3o4X5xGWYieaozoBv/9D7pF6xPCcIJzT7OjbZlrOqTRP
K1oqCZjU8nNmEnCyMjV8GksFYcogLcdKcBVZ39O85apc62E/yYhRwHs33arMv8jyblOunzyf9DUh
mpBef+fluZNs8HQ+TYP6ShKCgwF17W2MAnhdsamN0qrDEC9A1VnBPPvFPQ4lxWop6x//xW+gOw/F
F5cW7XLUdtFtlMpFbWkkavD5H7Xj3dN/t1OCcTT1VaKrYDe4Ht1eveFRT05rDoXWlo0ovb5NhucL
fPWKyvLker4FaMnR3gOC3D4iX5RdnS2H42nYnHiVbbunvq+zIUxyUhPBWecwFZYS8ipF7KqRYxqU
/1jkTEYxGyj28gVfJPvcPcGEZyRNHaqqyaqFR8AQHC59LDNd4HFwbmE4fQD9SW9PjrpfknXOgunN
ZdqfrsD9Z3EzQDG0+fI+QjJD9Swnv54aFoluBhbC2kQ5lIqhtPC5ETmW1sC79puqvoQT7Utoxjpv
cAJHggG+o6iMH7H+vOD/0zj9f0z258unl3JINucmeegEMq7DLB1ayb8uAA2hfiJf29pXtb+w9i4d
sRliIn6bGYqH50ThLBCIOtUEVfUkuNfCofppXGgojXaM7tMb/51bSdv7TdgIpykvrxz4Kai/ahTr
XeEEZhq0DSBmGkdNscnujRVvg7RzVnVsCINR31bsmSj2bwgW9yQQ+9HWkKAW5PJZSXtIgOuyEarQ
mfq+0hX23csqxxwb5lEB5FewiitkD2/Qpu4bSFrF/XZLgB8dBxdXnhgNuoWY6UQEf5O6B2RRGf+g
4yJLB92B9Iom1OL33iX8tJ0yRtt0Sa6lGNyF5uy6gB98n99Y4pc0ndz9MC2g0P4G0vim8sVIsH6G
rHcIOUseYDsfbYHD3oET7TdwlVRcsxDZRNwQN1Ci/ZNqKfHlk8E62Lms9LuL8GOc8915JxXThLWA
7vI8BnUHOWXqsrRNRUGDILjm1xnRFmCxL1EJfTM53/LzERylDLPd0AD9uZR9C/IkNZdbgp8tR5K6
EbKCQLAKdOWYuouFsCM08XrVkPupf/3IXICxcu+C87ySKZzDt4Qy/DCvRRkhInNuUDtWeb2AuHIf
fU9mS4sUM3W6JJUqgk9ad0Sd9i//P0+xbLmMqCJ9Jel0yTQYJSQZFxa8f1QtyLIjBB3oLX9r8cZb
t5zdEcBJ9cvWEuIUH0CiZZYERNvCPvvj9x6fYDPlm1ZGnSCyM1hLzQOSO3iWQ2HRitbav5iehhHR
lyXIwmse9f6rzfzqu6qsbME++JriHYPF2txeTETYcXu1VpFIjmqKg0aBseNMMpyK68nZ5QHtGrgQ
Tn2DgmpcrAjNAxtrDecu/GB8DtrEIdFMO3Bm3Tes+x37no+D7ryZ0xa/tRHNnSNJqBq1iAYTav4S
5zwOyLEchGAP6PXuT+d2Rr2FkApYegBGekYloCevrJRhpGIZQ7rKR9yssZg4ON+V7ZlRS8GxhpEL
uVX9ImgjMaqYik0yaWI4hBDtPcttpUVWxWZkp4uB2Bjg7EiVVGEodzNHUuyckfMZd9BabzVA45Dl
GNXB5v5kO0AWxUIG0j1H40ymuqzrTffbsq65Lt5v+6U8XdMbXa4Qr1YoolROjXtA4qo7jhA9zhoj
z6ghYL9Fx2efalG0Fp74UcbS+fQJhZysUo1izioH5N3S2GO7VvT0nq1fQuAUjidEPSnKjrjSKZft
niQSPuGPefz//8FeDAhJ5RhTjY63nBPj1xYgmxXpLSsCduDtYFiPhd9TN+fAkfyT+cQzXeiLOrCS
WWkD2PGw4NlU93kLmB8ssG6RNMRxvt/8P4Ndyze6lkxCGPUTGxP5BPatzTE9vb4IKMKz0RlOv+FS
0S8EHl7yx7e2qaDT2Xxi9jyauYAmybCNqapvze/8EYFQ2HNKWDjMr7NlvV4JgYf7hTmPmqZOWFXA
DCRIt+OebehOKtMUDlg2GiXWAiQ/68XZwBWiRGgPLknWBsncKKfWatTdpAaitLSfqAFMmhtVvDp2
wdoTBEgK8wSwFcpeBUMCFizvTsurC469v/CafrVeBC6ich9S9wqCOSs30py1iKe6G8Up/GLSFRAj
VM7REM9RiAsnyPPIByWvlOSRZxmv2X5PGYlG/iDMNjT+zTiDf/EesFnqMTxLZUZH4mZiY+EInoLZ
nDOqGweU22YaVb20gIUnC4HONVuJ078x8T3HOSyvK8GdjIHSu39k+WQxnwN1EycfmJd4Z8Bpk3ux
E6BmyiidlcJncxlFB1VzEs99EjzeLJB5sNyY14hEWtxlOHOyY1WZcbumDImSfV3tbZ4loLyDtIMS
qFjq/cxDPP7pnkn66lrrEUTz5vXGa1hhnYVAa3caf9ApFzcJ2lJJmEgq/BJGv0bPBLpH4QHM9gXX
02t+rQ3v8n5z5K2flhAJggAqdEfUDeBYy4MA0Q1VnGRKl3L8KCENX5/EvDYjsX+1L5H9PDfC/Wyj
amRdiYBfkgdyVyTFbx9lOwqk/EXRMzWLxngkde2YXvdm7Ai2EWS0ql8S29Xrva7ytSSchO2fNoE7
bsMBqu+L/vv7XPJoX80Hik/gLAFLcFrYhINwZNTFdUGq3XeY+zb9RDVJWspZ47zze599Qr2vGOYu
C3CQcWUoQ1KU8HPW9zwzmPhpxx8N2FPlAO06Abb1gnYU5NSILR7fe1W0F17abS+faZAUrjJS90Lx
FZ9xgCXv/HQIumtkU+nFuLI8ofE5QtKp1Tjo3ttD3fp1DdFCvY88iabo1OSwy7fY6jww8fMBW1++
gpisN8+aYe2f4n3qJpFDUpBPvFTkkKl2LEuH6WgOUfrlWhh+cQbaTbOrsUf8ewlqGXu0HDKElBCo
AWEhppCb917e21S27S5xbBQFvH/8rlU30VD8WyZq0F6w+VxaRgg0JG+TzcFTiutxdfOufcr57Dq1
67kHtWq99As0JfcWUmJ9TvdcOe47dS6nC8qYR83DnG+jMZI0nYguBGfpzR3m01wCfe6PqZXK92m9
T/dolF4q3rg1jjka8M4ZA0fm3WIzTnSPFWF5G/CPTftDIodWmu28kLO382Qr7hIGdv4JkGTk9Lbp
G2uBDJOCm66qyOHI8LPlVlwZaEKwGFLtfNNuXENEnQ03cmvf/00G0i6vwz7wOAO0w4X9xCTbrwSs
qBRojpZmCVcYv46IIti3WH0hI2kBVWEWNIMCvV8MxtA3Axy+HCLb9llfIOvK5SuT23q8APNvBbUR
eQjkL25kN/pro6NdzMuAjoSrSNY62fRmOsoTKLCjf4oLkN/RVt4df+eec5FQmpBaZYSipR2divdj
WOiZM4ld6vDFbmeGLwX0uxcJKVXA/4sSnOdLbuc8/9Fu2RXLIs9BOPpwfDFXl5k37Uz2OYSzbjb7
KgNymr/tiMp+YiaVK/Srns3fK0mJIAQ+tbO8RJWuRU8Woewms7Ec+QZqwKEITEkIPghD2hLAj7jt
sXtUJS/vs3TZ+z0Nt/MsHe/FU69OQm2zSAQIrfvOpuOk9/6a0V0mEJoE2vLMwj+NdweY3GMrci6f
2pfUQDEUYhu+CdADDOPSoy9AxUjmEKZq019lj3jI6PnWvmXWoCaaeHjoF2YAfsUuvLmUKKiN+Uza
XHtdfoz0nM7tU0rrUexzFavSphRpG4ZnYTXlkbDRdUrYNSQtEb11bpGBWH0+Rl6yLSK8hTiUI1nZ
LJS9vI8zTv8caJODBuu56NdL2PPazkWLLiwZFgqLRk9FGinHixSRBtoryOWJ9h0j5KoPUFsZ0rmi
fDjzpQF56l9Pb3ZQOP9wI5/mivQtdAAHKlbR3i/031dRxJ2Kkc/7jtsWZclkHFKjrKVs3bI14GZu
0r2J4FVoPPy6dDP3yArEBYyzrN3ei7/ckzbjyF0ZP4foZ1rJGj5g+HrZQk25dn3Kyf276jt1MkJt
BFX4Yan574RtDudE6XpVNZPiMn/jWe8NnNn7BUWG73QYEtcfPXGELCA86LfLCSauIJ4X2AliQoBe
2mKdL+VAq+RAGqpNVji51ejLgadcOmWI9zQxbRxXS2YFFoZ3c5v9JmkDCC0ZRRPaB0m9Cm1bKknd
AFZheNUsPEbfkioKgR2/J/FycrVKFohf8qK/k+UtpcynAw+LKvYvXRAi/pB4kM+q8MTcCMgC+Ye4
zwaoEIPfCRWJYFcngznIsgr02PCnvJUiNxN8KaGOTm9TGTg/nufEKi2lQDJfW4ZAVfwIHT1MgDTJ
rPF9rgsWnUjr3PWvf+9XTUSw4pmye65jpjkunkpbVBqQM/pR++G8xiMqD+InO4adrPrXYCAmDtKu
+k1GLDDlEMBtvyNgz7av9TrBSSSzsSi9IU6LOWrE6rhhE4ZS6pcrNnLuA5/qDYc7+IEDfyUNHVbe
SBaWbj5k3L4m1uRT+1TE+o/Jh7xhkQr5p2U7AOWzzvicLV3s+BVjI5bNrwxswJhI04IvM3QsyNCw
CHy9eRU7reE+cVTkA4rb2CA/5Z3jeJgYd6GjefdG85IT0qh+HEPfDQB6OceshbP4RxwfHYRTla/3
nb7DOkWM4s8DkrluUdblgN7q1Ujz8F97BXwuqK/MsQxkOQw1dlG7j9QaxXpKlS7QXG3E7G7n0B7d
a8gFBdJJfug+MNV6vprC6lzOrwQQkuPw0/blh6Zrcv0iFPnBTYHBveSM7ndSBzUc7JNwFnQ1UfKO
7/sV/u6hgAkVsHYcQlAOUFECNGeSvwZf+iXdlux6M78D2qsqERgTjDOPOxynkQNThn0QYsLPkM5i
w8eX6gG9xqZO2Ql8UGU+EkGRVUDXStBNlKgB/0oWTharrCYvMOtPegX3kCFSkfidlJ3xZccJyJjF
5+95JdHUUcQRzDX4xz55DTZxG1uifZuJHko4wi+sllpWfoXzszKKALxHkIwuUcNM6Hk1j1ECFjlK
pmwfi2oe7CCjXkBgZEttHmz89btlOXdtUxGdcbNEKb9vMeLstnoK50V5aPcsq2g7mTaA4iZt35c3
jxvwP7ue2WBa/kqVMEArQjMnms6JIKWLYabFbSdTP+jjX8xctZNsvZHFDrkU36cM3qXdvT7Fq2Nu
IZmg83bwWxJYRvJDyQ94rFxZR3kcWjdz6DxXatfVRKiDG8v/tgnywjKeV1Kzs7Mxd8cD/80FMqds
dfxGvLEaKwxMhu0EUf0ng05G/YAW+Q1TD8XteqHz3HlYsCKn3nXz1i5IqqCULkb3ZDxOHLHRqLqH
ZUEmIHBc8KB6v1ZIdk57KOX3bx44hA+7PFtB9ubiDpgw60pQcq+muZLET2m3vHaRRzl5YpuFvcnY
zo3yanX3ALqKmsTCf5Mpmx0a1VE3LHfnLhkvYOph2PzM5SEYqP+6HzE4PGLfRVDH973wpGu1El6e
nLb5VpmRURDRUVwvF7rf7FCmCEYyKmSWiRNcyziajdV+dPkU0YncKyQNRr8oFHtvkqCRRmrHk1lX
lPwvwzYW/NGqo1Ey+cdgqVvXKqBFZVlaVxZODmTrd2jnAXLkf6tFPmncUv3QC6PILr9UR5iFjnw6
XLniDn/xUxOKBYQKjLRh05Ky51Y2w3KcmFvpOHOY7HXQw5K7+NMz4ut9fWrGuJITQ+PwGaxB+ULz
BnO9vt7S4fj3+SEJnATWtYeC/fzXQNby8FV61hFad6jlwUTUg8yCX97+W06MzDpBy3Z2fFtu9/s1
HGTbwo5MVj9X4DiHxrl90tfr2vtq8NehcTtOpJjTBwfo1RPjJwBWdtMPo2tT/EjMHZR6qkjcK+J1
bQjIZm+lNclECBaZ9FDHgn/RpsR9w7H2XQ/fE34o7eWJ9fsqZfIJV67xX+46qXgCgTkIS4P3fYWA
7g6p0mJfjGpUXojd+USTmwgj4L3NNXMdLonVxXygwn2ELHLNv70KduwqoLLMni85ZXyu5Sc3SIv2
b/p7bBYxoQdvxmL3K4klBmOW8tDPWjEivR4j8/tNyBlCl4V4B7a/xsGtQFFUh7mX6sZ0Jef+VRNU
eydP8DX4DICNhwdNiMlnQuB6OIFvb+wKSFsOZub3F18E8ZfNgD5EeMz3zQ2RVk9U9NiG5QvLlcnA
QDaFD6RzX2uPMGD/pG6HQp5LaGO4j5gnExBDcAeH4W/uOGlEUUICBbMKXGFk2nkrN1y4KHFaQL6o
G04Bx7jeHWbigGsliogJsJLyMPkEE+3YFWlKT1NTMK94skvvBMt8DNUi1qsGQn1xJ7hZgrQ0O1eN
dNQZpvHk1qHiyBL3IBLuJ7ETthhnTNAdrb65dVWggMyOn5iZJND6p3N/YrLmSLjMdiBkYmEQk84m
3XzGQNg9N7k4VXiWkbH5OrzIT5s4weNtqodpOTuaBsuh+bOKDRwzWBVfgawE17B6WtUUyHh86oRA
u9yKl8aoN7lUYQHiSHOOFNDkL5auT7ZqFZ8DWESVYcYt+5kMlr3FpdwsFsHKldrBXb37ke8dlXe7
LGDIHklubtQnBHgDzOTx/pQ6hEq6wOjKaJiZGWCY0l9doPlNy05YYBJUViu3BHMt1eSQMSa8bVIh
Zc4vaJJtNR5Eheis1S9eCFOQ5SIP2/F2LeAa6bT84TXe6j9ltJqVYH9L7/yHneXuADFgpt+MddFI
jOSHgUlu9qE/EB2XJj1zG+bGFcRUYTB9ZLAhLgNrMkSGMoBC7vjP8LinUTwwNAX6xnpoA14X5vok
TIBQ17JzQFlQADeKiknpmjXfPzmD4eD4P494HE2rbYnQuVAzho16XsKElrCTRUvlbB0mx7ECvvyw
1nXDzkurKNABI8SgG5Ac7DKrxPanLdxVefeiVA2Z9CjKXSgeDNd5WJv9LlTqUFA34caIp3i/ehQ7
q7S0N4wTXBJ6uQ4GLXfzaV+sc3S0HZr5wSIn+jO8gZiQ6y8xIb7yDDEOLY4Gzs8yK/kWvwS2SZGb
1CD6L+FFXs1hTTi+ezaAsAUlG4jGH7m1SCmpEJ+VvWxTwXn7zxYMTlJLkeC+b584FsaGEUtBegQK
wvtndIrkXI/mDR1mAaPVa0mHAc3cKUlKsXWsm07/5wpLk3iB/Hcm6tboFOCCFHmwUWLF5sixh0U3
mwpl9hwzTsDZhhlqFqTLqv82Q+CPvMfhy7lj8M6g6iN1IRhqjRA6alxsKxbg7DFeg0Qj4yElZGgD
6xBo1cKuajEwrq+x+34rukd0nhDMV6ZYWl/MuzsWHsQDP9Fm9Oeo1hWI1nNwTs9XDSTXK0Ee79YO
zZkz5ETZj3JbgTVhoI5CZ3sB6WmI7JBD9KFgOS5ZnwGqDvGvx2WENimSz0qZMCifMZY+sA3gwp7s
QoImVORV3Wpoq+Eau/FA+xXBW/XamgeZr0w5pBZ6angHM9L6/B6jEFclqcVzUVA8KBvrsbDl1hyb
NTl4uM+4jQAOs3hPORz/IG6e0wg0djRZ92V00qFB86V/lWdzsKpuUsldqdU6YnZlrJougTIV4hcV
1rc1RqEOcY4t8LP8skgfoZ3NCntHbqKMZe0+w2tOuy7l5Sh79IZ42FhCXTchL/M4OpANQ824dnhy
X9MrDjpWoS6l+prFVGzceR7CpKy/2bmaCh5we+4XkHQ5LTxQggYlLDnFZaF/cdq2KbD4jgfsxmdq
H3BLOpTERpLdoGu1f+p9Y2cuqod5s30UvJEjXl1wMdD+XZ2GXKUFjn8Q2sw0sSuQ9fUXWDpYocmq
fYLEZhyK3xpIQ1cK/wAe4/2KmwMQsUxYYnsRy9ixr16N2AP5LZ8MCQ3aT3iUyvBXSTzgrY76w7j3
8hEZUjsA6L/hCXMYXi5fu1CEB+mUe1+AUQz9Q3rAuy8o8czSqfMtIW+LMBPTZO1t9g0YMEL1yc3D
/k1kAlQffeqjdP8q2TCkLfpF+g77r6nCtrKk/pIInhj2JefCNohJp4zfkBFXi9lYQqLO58dhWeCS
sebmDkwLkqDf5MoFZdrHfOKzKYH+v+JE5OdbffD/ClY01BrcqDelL6ezCvDLA8GTSDNQ78EZZqoc
Ov+fj0LkxBXkulI3xXXET8wUPfsEzo1vrogzYNIqUWtbG3cSMoZlmzAqH7Qe/vKa3/0034FVO7FA
9QhqzGCVwN8cs5aQAM5XKsYCRHNitJaySDAwQlLVMuHFZIiQGw4T1iRR/umYWJn0NGVsIy71bzti
GhQdXg6XfO0JHTDR8ClIGNxj3O4auorRWpmRIsJaUwirsK7WfTvFf22Z6AQ5iFts1jWVgOs3w+OL
9/rArepIY6aHRTU0BxjPBggTLj/OXdzVsmftFQDWwN4tsnQXEjBPi65605vs9b9ITuimuDzuuA1S
HhFi9eh9aXVoaVUAT013xXPCc/qkQkFtCpkjxcdGOnWqAuowWJXWVM5RhfY/NlQUaNJc4dAvBRol
UcBpzGO3fHZYuGq2hnE/woIzj7ZJTBmH8exQC3f5lHBUFiI1jW2dRrdIewuSTDFAPVfxKHlhjTxp
Go8yoeD6kuiGPRWyfei8w08cxEeh5FTxXPbRn3+bGjgP84bpabw5fgk9iX/Q54EqAnENRqhqWyig
Kz3Y1kkYz5/yMjYamMnnVuO5j/ghZB1ByRGHG+HKbul0dH18gp2Lp2f3uKgpzScYVvE4anOxbhlO
4vApuh3qbd+NMn6do1/NXjuKCMF/wsYiUnI46KTa7DYeHziE7wyjJcMGH/5Ew0hHhAiD4218JKA0
femXbhzQ5L49CHwygti9CJUezCwNqZTRrQI13Bhu1MkGHX6LtpuvFCmNwU4f5otG1o2LAZY7V5vo
JqUkCD8bnlDoI34xi7A184RT0+zWTecL/IS5D1pFyrj63IdAEPvmTRUuyKNH6xEZElHdS7TkCtmX
82TiTyHqeW0PFZEGAYQsR0WKYbdqaFiGaB+P0Dtx3LEPE4oQbYQ/YKd6YcE5IfscM+TN03Q/gfP5
GVv85uFAsAryY9a9lDRDIdcSrOjw32+Jh8Jw4yy1XLMtal4/+Lp/mVEK6aF627Uv0qnlIYwnNE95
3+j+PSjHCjnuRBd/B0Oi3L9YCVB2LcEXG/S8ewiRGyxBT5yqBqnku4CEU0y6semdbb/FPuuzvKGf
V5qFPy/bUXjHKaEE02b8b+63K+v7UkbKMDszN0C2rwiL7E2vx3/yeV+2xuZpU9jxFf7JPatDmU3G
HYcKKA9IQbPOuLr3BlDHK2+o7ERvRsgqAd7SsFhnwS+Wtv2xNAH8LxTP0Gf1FDreYQe4hjmQxHQp
S2kk3Ub/VoDL25C3hG+1yG/m5mYqtMHulYziLZfIZ0UvJbtwz4q7m+1lM14ZBNZAbQvMeIBoIEq8
v8qN4fg/wY7DIJFNev8IXxWqIy23T1APgQf17tz5naQZ3MR3W2cqZ2Rf/PiqL0cKOxpHZWHy3jy1
W/KGpsxsVoXXnj31iMgA6jJIeNFS91kzLlriq6xmN+YMqVGbyJbNR9BUjFds/trgXtiMzhDiWMm1
W5WWMkmblelEp+6OBYVHqA9gFdlvCTK4pniGf1NYASMbBaTKCMBwLBPl0Qe6HPH8OkzlCs/JrBXi
9LaVrNSWLuou1Yci0DZ0E8TSZ98U9s6F29zk1XNIwYBj4mJ2StgyiHUhA/Wbv6VUlc3rSohrNI0T
NwIRZrK/yIBpKxIcI3NpD+m1zghhaf/cUgtCMtUSv8cErDqsCwBz5XV79/VLBq81eg1apRY/Tcb8
k+jP4W7kp8kZUO9JCakUkwP/jQzWQ2LGYxvE7wHgbLJphvAgAY3CwKW1XGEAPS14y1aKWpPFnJBq
Fd1YY8/4trgovZN11wqIOa6pPPrcXpd36o8eCDnRkw5sc3LpAeXIBykR3ZNUIULGPyL0tpkAGSha
RFQdkAgr4bDEg6Ih5dz6e/SF375/lc4BcLNgNZ0+TOJMNNEX6fcfKMOhSRCOJN+Pc2hWIabhnVKx
AaVXYiCH1vxsEhzppWrMlUHDt6FmDulsGDg9t6ZErvtxo2wVeKK5U6di6aN2wD9KeADitHDN/9lS
2agBgfscKR5Rmyy1Td0cJO7TKhV3Y7eDDsvo7SJGM5QyhG1hwgm7vC0AmHFM1o+hifpkMLEkcejg
h/KDNMFHkSta/LWek4ORzQepOG1q3rhRybrmsCZWrnAjyX/dKY4UdqEpFBvxV7iqn03ow/POpX8e
hhwO7o5LjbwkeFVMGxWQizhkYH5SUODnljGgMQ2HzCH6SxMkMA5pYCjJcDuJ2MD9CnLgo8XwRrNh
feWrPlqsw9IOSsq9PIMsEX/pmxNYiVFn8S6jcKbOzCa5R0w/EFK/DZB6HQ7L6ivZQ6JA5Ashjb0V
VDpZzf0l6nYKYAy8hKPQ/LGRAxVHbZNod9HxxbmhCHKi22kkULJZ2goiF9VcbrMCQ03UKbjfDCKY
Yvwf6reGBdPVCpN5vnuNT+//hcS0lfF7o5Gq9lo9Ezv+pVGFOfYMHuLRAcyGdWVEPuWxlpo3grdm
f63gmjExbA8ymfjZrPteaUKB8OVZgzwCvck5HU+YJ47/mvgr0gySb08Kyv0aDCgNvkiXMsc4PwSL
e0iFXLyKs+nSCCXDuPOKbiZshH2kvJ3v1+YBEuh5VX7im/TWSsZU40kktLyKb5Emd+DH0E4p1HF+
fo/uydMPctMjtoSjTKHKjEURfbRS93eML8lUcLvgzT6bG0Wlgt3r6Y/r0Alm+MpxSj1RHG10dbij
tnNDeFVRUv2YDRjtGYx1QE1kIznEIegDqBR20K2U1rTrWc5JoqDnAxXmq+YN5vceC7Re50MGgf3z
tvKggvn4t1nBI/J2O7xHDqLEGKQBrMFHSMtKjEN3Cj6tLmqriXnwCgRPB6gtM2ApfCs2QA7EfiBY
C5KGEZ0F2zdNVf3/I9f+ho8sWKclwR3WZWVmrnCx3jMz2Gi5AFNZeMSsptQAE68DjBMGXnhctsIs
gX8S/GTWQn0mvCZlFDycz0+AuNOd6nHleMFH3fT/uT+5ZbCjDGYqjygEfchwsRTeHTFXW/Ha83ce
0UUfVAWG2CL6BpNQHp6FaFIxdnBu/YOJ/yi1hwzovaKCKqILjtEyon+kwtmFLac3XWwPLftCJVfZ
nQPD6pzn49bCjdHiHPrDLpFU70lMS0/fbHk0yPzMGFT8ufgLcl3p60wxMLdtcgrosLf1rVZ73WVq
JBKJA3EMUivpDaKmpOWKurXs8BPwojrfYN+uKeamVMKhBpyq/bHDDDT/bygZ1i/SX+dchdEMGaU1
kNn+RFxX/Zt5lxSq5WlijjNmjnAcCveztZvUU+ldes2OjXGv0lv073yCdfARBA2x4eUw/ZTzUwv8
cHUwhaxJ/ZHOkZo2Nby6I6RlFODLsADl+X4RB5GxVquDOUER+REgzkPUxdEHtQYFJK6SCC7nkcLH
ZB+dfRI9c2mF3qnD0Y48TAAPZ+UBlG1NkYYOEk4cqhgQAqNsspjkxpp1+Xzb/VxZAhvZAer2pld/
re0MMJ4HO95Kw6Zf6xmCrw9r1FLk92GqhmtfnYZ0GdUSS0Cm6lkSNvG1QaayMkJOJaFD2YyxC931
lGzfXhKvfiPahD7NqXFLHqJK2S1AYZp0T7NH1y+I4Q8HrwPhItzqChvAQbhFuo4rqth5uHDOlyI8
Pguz/RZApgxhcSKPWdqr2SrsNWtUgIrEViPIMzt2dFGjiNuxd7gnCFvG8++aT+R9Gtb1P/mekr95
51RnzYB5/EIWTcONQQWoQEvZUXUWDWmpkavN9RQJA/V4l+Cd/OSol7fr9AlW1v442NcsLg2UKi+o
XPefbdTxmYPmaR4WyA6ws0LPkbe8kDpSAD3xwW8tqyLClfRL2wLtqWZhY+kc8hSZRHge9X2KQidS
VOZ1FjWoFDmV664wDLDnaBosBZfgbyMrOsyYavJ//negqkRkVw7eatOqiNbC0vcHaSn3UractuIG
5MuWI2BsEXPgntkpR3UW3xjFl+qnojOF2f4ib1NpjpiSaQrsOCUo1oZamHoGvlNWfGgXF68Jwqpc
VgEkKgDmhGKYSQMjhYCljMoeLFtDy6bQmiGAGRiUndWE7z+2Rjd3SZsk/QhvHgQeCbcfkCt5a/Cv
yq2zoSIEh7VjcMKtRgtP0oEJfrmr2B2wZ4x8yBl9SfZD6jUAfMOBEfOof+nfz89PWIaH+00UBJR6
iEETqbBz148qQSzXu/rELn47veRBxw9EZ88IHYgopBOfO747kL69hTbQRVk8Gz/gNmTmpj+Ij3qg
32GhB7kmKBAms14+wnLUypnKXOvLHB5Xd9uAbm4h+Ep6gbyow7Sz2xzMX/CNNOv9YcMD3QROG6Hv
GQoRtBZxHDmZEQ5V1YNvAhG05Av0d0YOn4YhK/YBndg+/awKBpmym8eGPM2D8/YOc/KtyUEQthnX
jols5q2z70uNQZS7yP95UTGfnBzqw/BZ0RZu5vEtynHNSYm12D2OphrucwVXv78hLF0a4X7A6zF/
xoIyAoyXhO421PdSk725UU3JlxMGyMxtf99n1ddv2stYfz1C+V3ttKWIHzVRtmmABNdgFTl78dad
n4wT4xWpVvkRIyV/Yjq0aMIz/qjtEBiALz+x+K7QbHmN1t8fkYq3/dvzjK+bpTLzL2LA7URcWwsK
cD5y3CAwfTJrvz1loksls6mUK4wHNInQSpj4s+2btbxZh/x+9m7FlS27SxKu4MGRtQV9xNglq6R2
40Sw6G5IAX8gwYTJ96bJtZRsU+IuWtZdYsS8lPW9CAkyWEuT6mlkLYBM+tNN1TjaRi51Pb59ugIC
fUUfB6nZtNGvsZVVupQDudEAaHlF5HVLjoatF8ejby+dQTJslikwAKyKcBtn9LWGbi0SXSpWOoWQ
zsiual1VVXlukErhKYcqYG4XBxZG4Dvm6xFpQx2AFzDXQWAUtPPWSA5wP/z/2OjmyOx6i8r1SrVQ
OSO/DsFKBdtyDmSROnMUQWn5RdKN3X7OYNE1fi17GhGEnnAZZSBv0Yet11W3CI+PZRwWszxJ1ZJu
Y+pZ/ViX2CvKlubSU4m/JD4zvL7SOvXlQfLaJ2fVCtP67/3/9rikkxWDDLjTB7XbvlHx3x3HhU9S
y5JO/I/yJ/TviOX5KWCFVLbnBebXUi0YQRKGT2ncjrQ+ufSKa/OmbEAzAlzfTXhIe/apFLV7X0uM
lIAPBhj3bFU+C4MKJk6ldv8l5uckl0lPGFsfUIbOAfy6U6RZO3uDGzhjqqENUidSJ5TcKGfIXApM
MwidQgjaLqStmbiY3Pvbf18/k44ulz7+g3FsLkg9982IP5HBHEuYlMmNTVZPv55BQoOeIFN3sn9g
1mQa64y6gJvinghA3w1U5k1Xkyp2Ak0H8rd37sWwNxbcH/b9QIWLD0ccfc7IMAugPW9ghJbCzwDU
89ov8NfXNNQm3zbx1AAlJ0Su5v3ufn0bDQURAcrO4ybEwjmSgZ69J+20QQ8sgbXllqjmw7Md8jHd
VhXtfKe2lAAK1RKuUB/moaL1zYbVpqrV8YRqz0Npb3X2FbUneCZYuglqqxLDN2OdvMat8OVsam7J
zMVElFNsFd8k72hQwVcGW58FjzgmDB3mJNAUzZq6Ik3YRK/08AgXyrN7J+RylODfmfwMlADmxmLT
WaooHcY22ZgG85rSbSwkWLj0wwjJkEFHyoST0DrhR7YJU1fuNHzqIBNqQoB7GZe5UVWQVYOlr21e
hi1IeXpQsAkjwSIKMRzR5ocJUoeKB9Bnlxj4Lo4EQMh0C9Q50yst/NbsiiiSz/LV5ohO/R8WVSp+
ewhWc+NNyVvmKAYxmvYiBh5iikpIAxLFQxqF/D4bN+67Pht6atpR2Nyy2IS1NQ20Shj/2aZA0ODX
xOlaAoOL/q2Z1UIZ4l27MJUDCSpe0rD78ZjRq1s3B+tdx1TraeIhKfn02Iy/ui/Axog3d+qv5lWY
bDeb5YUn2PRfazt9VpkgQ5ThSsgMOvv97nzaVggbVH8jeGZEoQSAGvHp3RUs4x9Pd68E8P7q3CJo
44E9VUkRyMRqV31yhBeYxL3b5Cu+vKmALLpyEJC70FU36QUDZXYU6hNu4Ae9QYhErm/JAV2GAtWe
56THZb6W30B7M0tLbHSZkgHcsV208+8wEaaUTB6iBlPTUffOYaTjGcLHEuJN7Lp8BfbLBBmzDhqe
b0s/HrCzQcePpBJ70rOhmbXFDqnolnQnLY7V6yOFnFY8DPw2kbW1qlZ9uaHeDaQXDsequ/cdysbM
1XlzVFJdmJacf+Pnoxe3LGrRQfuy2Sz4g5ZAjV5+yviPYuiVg7fANxvH9PqL9wbcV7HistZQG3uF
JGTKclbU2Bz/ns39t+nOka9QnaFSpSDJRgaf6yomKAtrhJN8KuDJJdH9s5tfb/DM4r1FyVaOOm8t
NafNujOZwDQQuuGEG/DV83R7TWt0k1Ieh6NkZeX7HH1muWrr+TDdOsnahm1LQ2McsTMSP4t1lNFk
6xC82lf6Op2WFo+0lMdv4dkZPgRLv8WSqfw7/EMF/PnMhnaHNwnI4Xx4IHVyKndQjjYNoI4ZqWx5
y+vykdXvtifvBj4YAM/GAoWEHOz3apAksYXIa5jIIVvdonZ6hPCEWmnhgxkn5QJAvKwIePbdhfvi
TsMHSxPVqYKpQ6zANgS8AyAPW6r0QEgD7iYtXbwuqUSTeuLUSdK/1OZ3W56MA772H8tSmtFP14Lp
wew9tRs0glBNnILTb5ZXzhyVFQky+veQwZtp8lPEwJYrCixNykneklLClsC11vSNf9umFAOujOHd
4dPSb0qoEfdmRsxi6VsF5UL+6vBfQKS1CRhk09Au2CWX3kwooOu5CuBhJsMn2EFLLDgBRGxkW0uW
B5/whk2NyyssQeyQewesLp1F6glj6IPIY6Jv8KkC4iKPI2+XsnLyPwM4mjZ4YYdEEj6igrifKhRd
RY3FLSaeornmYsQ3BSrc23Fv+bXfZtQacT5aObpniGB5A5fHlQHhMjPnNu8+fm9DwmJnzKbFO6VM
ZVuLkw6pART6Olui1Oj4fkJrOsy5WGmGLlInhhZXy/43Clw3kAvO3cWJCPHqtNXwTl9XkKFlVRMt
J2naOx/IDalPvSZOgGsrmTNGBDBdkIyn66PEh1kCA6ZL213r3mVxTTfDvqseeByHW3VO3+BN/UQT
TwuF/uNkRzYXcM6i9HYQf5PtCTjU1lIrm2l6P/Tk4v7k9NhO7UConDTILQCBK/EpbfuUdjweORfv
H6zR0I2zfCMGzDA2lzp1osVsuVpsX6uR9/BGmE6IPnkbyLjo1zpvWctuKpgo63zC/w7kNXRau25M
SQ6v/ArbgEdnNj3wKHPfh8/NSi8VrxCpcJZibIP+jh74ZJkSL7gGCEnuIWoUXjBCOyhZ+KlhhYAp
/BYVwAQg+hIVvBGsz68lTNpVe4B8b4U25/XF7nkfNTimgGcLUccSpEjkDV1SJAMskxSkfzAhKD1D
AzTvGmxlOrwzvdcp4feVGklFRyJH0qkHJRpVCXxtHDZA0//4oCW09rkux2NabIly/lN8mqgJUTyA
nGQi4lmLdaLAqCP9vwbhYVidvSCtNkGxorFH6uZh2Tw+eUPo9sQyB5/B1my53SsSw9C8vAWYmw2c
VyMjNhE1YhE0+1ahVzrZp4F0/SREiNvFkMhJcvYqCe+Sb+mHlKELA5eGVQTb07kcFEPYqEJIA7wl
csR906KTO1LbHHFU2xnhzbXvW61Qd2xcadf5qlmALNwaYSAkjfCIlPyxavMyzlKsGsMe37Gr0JbV
OY2nvV5pgFaJJ6dS/Hzn8PJ+SY6eH/5SksM21VHNDROZqC6QEVE4JhRr8ErxPhTQ8g3r1lp68NrE
7a4mpURnkQXppsRFnTcTUp+5xHgqwZzKTVJY7kkXPg620YE6NEQLLnknXIuJcvyZWcMR/x/O0V2h
bVTOajsfGv4iHrygJN3f2UlRJN68RUAcEI34Bx/AnXk4isfGmItvXTAC8t0Yfmiwd6DkNYVjRTBe
wIFrHZQ3+q0AQU0gs1sDNHa4X8N4o+YQbRCUiiwuBN6ud39GzUQ26o0qoFeqf7+UX1EQgQLosvGa
38+ZishuCuMwnXWcs5gWsTHBrsrGrj28G7D8lQxWhrq2x83gqZ0wZoHoC3b0a7/usqVwc8BnzZmk
gcfAJikfjdMe0mJo9xF8KeNGjjq0FsS7Ur4cstUQCqsqxN2njwdasYD/CqpR2+Efzy/61YbPH+P/
IHhJ3m+QKDkrNZbTbhG0tsute4fTQ+euycaZOBY3usifp4b8mxVU5FfvKBvYS7dazojAQC0e9nPh
//d5FfzNpocMOQRnLSd4jryaUbPLjpY3k8+Tq/CfTvjnkoGzygDkn9ieHnrJqQhTokSQ31rOPoeW
RUquZ0JkAC2DbbGPo4OiVwgqVC19SbQPpFjQ/Rdjn7pUiigklm0La+F23jK0kl8u3lg+wXaoLebh
5MqzA4emgfHqru2ouwTOgC9VpAxqe7pE5unoMbfLRbZ1LZg9E2HbjG0dblElTS/2nea5R0s+krLc
FzCshvkwcG2FPckYxwX575RZZVrd5p93R0wQh+ImqyJ+xsUe89tUtknfXtWpuXvVLSGBgrbqTcTD
VHjrCZ7EsyCi1nTnsHZ0BkuuZ+ziMzPFdYd3a0MZWudKGktnJAsYPalxM5GbfJpB6x27d9JVk1fq
aI0/vbw7YmKENym+YQSlJPwdsQ7SsZwawvYw5E9M4qw9nzTrOnhrF3Gw0NI4+HCMF9hA7UOJniYG
boMMEfCgedsZmDla8HrOa1EicnsgYwvd6XK3cECc0kTPewEiy2W6CH+wY1lZNE5zLUPdFgHMnwCc
nwao0LRw+SzrzyN1AsL4c2jep4X+opuXeKhjPssQ6zOSFre+KGKoSs8hfGFNM3rykshMN8GOEytf
yUaOnO+Mvgs7dR5CG6XdTbMitLSB5MRabqPpsA29Z8UhPId87QBI+iNUuefzdUvXBaSLit1DCGtl
mooGy4PF20mjJl7nqonvF+FRCIctwxGMiDxgyS9LlioEiF8UD5RZt4XMTEgbaxbb2KNFCLyo3qeU
ZkzAPp0xhhIsZZoGfhzK3zsN7fybJsfml/E0FhoJDMUtiUG4rfwerj6Rxp927yKlj+zV4gKWiEfA
tvhWks7rnE5FLHpD6vHuVbudOJYXlbZlhEPw+r9b+EckY4rU/2jAApottTI8l1pB67NKwet/Yngo
gBC/Sg/mEJ6+EdvWzun3o7fmacE0+MhAqHxtQyp5lumX2tm0kYt1h0v/Ak5Gn7DSJ6h7a4T4UCX5
UnaFP2BFa+qfvRlfs4N8cJ1e8j5EbLglFyR93jk4s8fWf/XIj8eeX7/O60NP8BvZIOeWNCA4AffT
RcZsBLI3X1taPZVQcc34fb30XjV2N4KZtsGlhCAOZZL8X3er9lSfsb0GjfPhSv3Z3V+6YxKqHdwD
iOPE8/o4vV3KGhfJFlFe4CoxJkC/bDqUwErp/EpLhIYMZUJGCL+H5rPsinnVH6UhI1THhf4mT+xy
DsLkV2fuWXY+Qt41FJa0LMYWZjnlWRRYErImxvUhd4ynmhtVBI6AsTSPdipkjnl5LmedP0nkScZS
d5xWATsALGdIjWHS4JQpJldj6jKgeFQ+rXfHbPSd1lxhOrLPRYpRvLCZzpg3ipLd2ktMxqxbhy9N
ZSBL+Ly9xt+HsibUz7om52ryENDBXzAzP7D6wkZsBfy2FcGanA8kUZsHsZn318LDJ/b2A49vmDrU
K6VHRnwiewrk8nBS0mJbcJzFeYIw7x4oy8Rk7xgcIh+C9VGs6u5zNMqy2erK3Dsc/6Go8k6O+cbK
6g3w52x9p0iEbjWxdamHgnKfi0HbTL4fZDFLwPjziKifsLJWlQvzLmDDKew8jsM+Cy9vuwJjSkRg
JNhtpbmK9J1+1zmfn4Nnw0hNSyj5aJFn1ieNgu74Z3DP+Ows4F5+APgIDwJBzgpgt++WNTgVhv+1
Lw/PSHLsPgwmuaBXM/JinPYAo7OImyd+ttjGf1wcHDfhiiNGsN+C5Rj3HeUjZDYALeEZpZJu3rb2
XkW5WwA7+EJJ9wtDn/GQcAcSmNphD6lfrWgKDZwCNTc8eHW8ZbKEcmkvxqqokm6p/Hjuq9O7I02a
U3aPo7AVa3B6sSot7YudmAD17RqToLE3FiaxgRYvKBvf5NB9MQaUQjioahfMrOPp6X/owFTwZFAL
wBhbhT1DO+8Xu+H5zz/OTmabYc+S90IUxlio5fbYT/RrWS0yBDdjANa7uHapV+suc6kfb5l9Ebii
JgOK/z+ubJ5+5bIhEaTstzs7Jy2XpOQ6llDRmoJOrywm15CYEXPanlfwNbs7qdA3NDHSq7eG9dN6
0ZXz5OPOpKUH//oAscO053ZutiiHa3fNIqBk2zJzh+/9Jog9QIH8Ulh3ocT3t6RnIg8Lt+VUxDb3
isSJd9pB4CRrZj24VGrYzfzh9r7VlSCazd4sJjdUpLTUZ2pYWRJ0EGjQF3I/mR465t6lWYLMIzVC
P7tZ3qJREkF+vK1neQE31IteIkWmGyk1DIZEI5Hyu7lTniZ3xwbUWuu4GaiTFtrchvXPvlbPR8zh
aASE4Di522k4x8A0nQ2UIAuQtn6e0fRkKpSzvjAzRKruLDE3pqc0XhNSsJ85vAmWxz+7zYqa7A/g
zhMMkz3Zoh3fl+ieDrYbyKrvA7QngrnO0jFXdiCWhFvX9zdV9JTol9OTyWiLVEzgpkJY0MeVf9Gr
6djiRWTDkNmCETYADOlpcHn4Os89fx9bktaLcjD+p6GDG4aJAcReRXw+djMwYWwRUPk7/AjWAqN9
2N4Jk85N+ppprMFRXZTc5o4Vk0OJSlOqQ9sfhvaC0nma9lJHAD8YJqyD91jDlcaTQgUHE98jeY6Z
MkT9jjiMT7icT2EVId7dilblbV4bQ4fW6saU/SlQjRLA2GLH5UA4SUXU9iAaB4vjWJ9Q0wjGNn3A
WGQKQX2j+nOI7FWa2RYrQlMOdyLUEKEvaTLI1ZqJ3UOoo38BK0xitC8DFg8I0aYJWTDa7irrLCtY
w1dPUMRvNmLCrZoEadE3J6TbuQ1MX2OzxujyDWrgm3xw96HDXm276LfJ0h31zVN/EKjPUJFbp1rQ
rgzhLp0dA53iaMcIdzfSyah6GreCjy8+e5UMuvoejXdioLlg23hcTI/8vEkcdxOuqH2Pu1t7RjUj
rl6LHcUJ+6RL05FR+1xBXiLvdRfBmeHE1pvM9lha03mHVIw3ocXMjBwjKhDKC2kgBx7su/F5U3Nl
Rv8eGCSBZynOJhyW8AsEO8UxsOQuRYWk8vmptDORjrjVHvucvQ4hYbIIiDqaKV3PJ95+j70mbLMS
XPPdx6hnY7hv5+tSRrdMLQVyOXTZMUy6LpEEEEvpZuE+uG8NYj02/m77yqYkTJGZGEHTCcWIdgxp
lhbsbO5BOXtcxVFHwsihhq3T5VU/HfMnJhvUirzbF/mrUOupNJirbEyDh6ZPXYb4bSVqueO9yOrV
8m0TqOnCw3u4fH/meE89x15+x3TJbrj/r9zC/LEHqfhvnl35ZJ0pk9O2TRoqOTqy7C0VWKpaQmE9
OH6xlT+tb5jMK8aXOILtSfkgHD2gpy6PsbYGBtrvRs2ZXF/YP1BNPn5rP8ybjYop6E22HeGGcLEi
Ev6bXAO/9irwhHg3n21jDYa0Ya5pSgt2aKykhTbKaD49rjkUJheOzJIr6CP6SUzvLfVYjQG5sP43
ruknlapRDZjehmuESgC8irz0hys9U06552na/VDD9jHCEs2njWp/MS7wXU3k7al4xLQB6cg+/p5A
0Dog44A66akDQiEXEEgMoYpz0agEHU4LgRoj5Zx9Y+dFq20x841OD3OACBY3Y30V8Sg0FU6borZT
y/ys52XayniGzeEgTkkFDOp15P/8cz/JKwGAxjfEBe2RXa8L5rHTA/rM296UDOK9VAVoJxdY3XCq
KSyNh7Krnivl89TuN/KFls7ucBTTUbM2af8X2fnNOeHJXNhnmCGWCG5SH7QGj7A+UwVksMY7bxTi
tIYQZTI/AskmRbyjN4DGyG8yW2W5PAPhoOmFI+yWbf37TKQsgabYc3nhwskZheXuB4OKH8hhlzvA
603CIlZgpDsMRvl+EPzDbkOkLJL+d+Pi+oBrqzt7oCK2LcP7x551DMJxR5drdTppRpihAPpw01KJ
3TXOFAeqVnLDqfgA3Kv962/EuLVgW18x/JKXWCCbLAQAQeKBEh0d1ulJL02+m00bPHjiiy+CyvPM
KRa1xH8RKRsX7Yi+ejmYkkJlVKf3Dxtz9mhtFhivFPXhX4YbF+U5ooBtFrRxfmPCHjk/XHHqgYRv
f5YHhBd+YlLJpnygTP4W3AXq9HPcSen87jdEfAN9yaaJbNWUBQHZehviHvrZyKmE34JdaQmdzEdS
UgQJ7+1P40ZAwQGkK6sFkZgTylfxb+y5Q+Ow4SE3n6MR1xCqaOnRbW0IssoNVw92xj/WXI7FLfKk
66HBQrWgDI6zXIdbo+agidUkr6rjTVVh9PdfYnmrHfwe6dD1tsXlMBdBKZ7ilXrwmE+p+YdLhE9/
vU4Sk1wk5/KzJ+dfTPQjxrtqtg+PcffEL9EH38simT4Itdk0qkGT/NraEA/pCG/kYsq3wxzBjWrg
GF3om/XMkblppAdcuXyqhRTeAYAr3oPmyhVxClZGSzjKHgfRUaUwrBXH1D6hq1ubL0MBGxQCV9R9
ho/WREEZtMOB+85s6rcL7hgk/gGYV0nGFTwE9v+1Yi7kPMHXlF2b3dw7qyQW86YZE5f4+UXMOJ8O
74hY/XVCthNB2XEDwYJNPyBcDH32qsOWxvKDRoGHOkqMZepdcmlznAU7sgP461tbwaDlZvgZdL3v
Fk3mumS3Be1WThTBxveEuzgK0mi+aUNZJB+SwG3hChAON+v16MWDSTultlnHwqPJI3Sqi+LgXmLZ
ib3VXRJUlMszXnwL5lhVpQ/A2RIqus5LOZ7qEOnPCP63SLO6MBIIUbp75HNxilqCE1ZlpXnwHG8J
Qs7mGla7Pvn+vzs4Gb4+xYvVGi8S6FaUhOgX33wiNsuQE9CXuL6Go+WYQUZYeGEWSa4UAypfH16j
P149tEyi29AyDgYosvWUTIgaiN/gOA08WJ1KTuJZfVOGPFlKR9BBA4WmOPkPY4oqYUMBcQXzMlA3
PSda4mAv6MQcBjHB8czSvTME3rRYO7FNjjfSYoCb1tty9MIC7Z6krvf1cv3pdtRa4zaIXKQf4CPc
tIqpDWJXV5NSYpzhK+7xAinT46DhRXY71B7U0Sz/eGPafrOsgCPlUKtkxx7CRanKsZ0LC3+cQiaF
8FZ42bbadVPDhtyrvuEN0EKwAG1UKFegGViaIcf8zQ1Grk8MK5ypMgTHq2JdSeUuiML+8AWyHvIl
r+QKyMXiVdJPgTb5cW2QZG5bAHxP9qvSbMKP4oDiAAL/5fWuTdwGwL0aq6fbGnuPVGZx4qJrfhPT
qBYrucEHOZw3Ckpst5/5/2hTBbJNQ2MMLU1KNH+JQcE2UoJvHHh8JnyJA+wjYuLkqUgRzlgPQ1LA
ZTE1YIgqzHFo1k1dnqhRwUr8dU6f8nAZzbanjyI0Dk9OYrhjWnk1LrI8ewSQVJ6JdndmCO0mhl1F
IF77BRMb5AKpmvfVIn8SGrzSm9vE/n4UZiFqDeh3Msn2f8/jr5E5DKeaPc0slWgABbCzd8L0p6yg
UNmj5HcN6YjmZG30vlEY8LaouwzKUb58MQ3Y1J2DHxjAPHQH7gc15e5yioCFFWgoLsPYwBkLw18u
9CcAcfYUr8DqQpLvUmpbEpQnRto9Q2IzGHuxg9SM7CrT7mKk2nujLwTiJXsjNzNGK1jy0/6sg69Q
8wCyKi1uCagJ/WgOO/2c/Fbb9Hd5ngn+m5Ahh/5IXfKEvhE51MWJF4yUxQqCSCzyZFva6kKU6fdl
nuMHN48NKtckgqffUK3uDrGfKbcj55WfHqQQmLgp8k+/7hnhkKwAWj8bpeLS2LmYqz661dewVw2g
SoN57A5rQ9G00wd1UE0/Eq89ZfkYA3V0z8iVFBbopOH05h6O4EDDTxz2e1lJ4nabb3ovbhOuAhHX
fbsfEClM7O2rPE4sAXJlpcgDp+Xy9WzcTdhvvimIs/pp5kz/qFmYFhjtno8p4Q2FAZKXR/eDIxXJ
GHtK0AKrjDPHRg5MeL5F9uyqHKJvfpvdyTSx37r5LXClL0qpzrycmbN9bUEY1sjdk7QThFV7Yrlg
NQhGP2M5u0tS9v9hg+A20MRJ8kUUPqAcFPzhbS/cIXpQdqG/mW54BZ/BqVuzmXyP3Agz2G9biosX
IL1nUdyogdD7a1qTl5z6xBWW4DrK99SVoz7TzjFCo98B2KKFMQmKuNPykoojQICdcz8t7CB43siy
2siY1QAlP6JeSwbtgixv/zmk49WR1DmFQHZBMGjgv/sdW/tT2V0ms2dewrW4qF5sDrPWC+hDHD1N
GGI7dGVKnj/LQuIuSBI9T7pT2Oj7bdcaX3Klo4+ib6+beo6XiIBE5Lca2bEpwCxME5uBkyIdBaoI
LCG4NzPDnbrVrdAZIm9CMjI2YAOqRuZIk4xIMc8WkIdPWqNtfpi8Hx6yHyTzaYK7UpWcVQF16q0+
0yX0ngHi3IsN1CMhk9x1cQ3Di4VrfYM92Fh84Xf82Yru2NRkKbqnfw0Tv7AnMlQR9sjg0O6BOaXB
mQRYNpjfPNtZ1JD7mS7PX1x7n3VgyiIQPl0BcJbQKsgI+XGYcY9xIcLV8TNGDyS719RTEJfq8fGG
ixwQ2qymrjz73YZvPNxNBohg3+l1iCHm8HSE/WCAxAXLC4iYTBDKV6Q8tXUY/JDoAEmxb0ZwN3rI
7AgVar7khyRJ8R1acW45w0/e+8tJ3nXWPEDhSZ5sM4hc+kOEekp7ntaZU2Ah8dxUMa2fAaANzKRv
8Di6JCiBMhI8hVys5l8WCU+soC8GL0gmEwlefYwdknW80F3HsDVIPW73vFzqTrtlvrelpzMQuc0m
xWvBQDgDK4xFceun265TuY5ejeymAXheS2Hk1OYbZOxRyABTH61QD+g4xBj3w8JQCT2L+m8nH5ml
ITFcp+2IVP1sMNA2lVySQQQt3uw+Zl16J60/Zi2OaiD54f+LAKEuh1DPhfg28D+eYsqAmn+Js8kl
0ox7GgScz/SRKKHsxzMNGP5B3+McXGPzmcJ5hSd0VeIk4EV+wSHQjf2/Icj+DP/5eQloaTjONBVE
Nc20I2CPKtD4MurRgB7Fl5HquEI6qBSs+2s4TvHIrMs0+715hBzoJkUxYLiXovGSWTig7fc5IWiV
imZU9B15Si+bcGcWyjAKaU+yam5M1vF94P1R86Jye2M3STQXMrGfeDtKAu/jjhz+nq4yhj/fjsg6
QqEXgYLPzau9HzIJ8WGBx6JWgpVL5V32btAbmDRAeVsbi5MnyZdqxwauFo5EantalkwAvXhvi6rX
Hly3cJ1w1JWfcnulI7y+vjiOqhYf3uGikFdkMw0CCXQGVdO883X4Qr72KYqX7jnInTH/gas5j15C
Nok1Cr6pahWqKJYghtTo2sB9VVqDpymYpAF8MtZJ7Go9Lg7pFfJg31wluhLE65y0IIFZJbdS/+6E
W8HBvmIs8ZZEEYZDFgQiy6tdgRliEI03ifIVIK5gdBoDYCiMKRAfEyBsFfXHAR5lIFKbF57mtbtG
MqxFDuPfQaEu4/ITIiDEKNjMiRdmovpy1O/MXRAIozeg1QeH/cLhX/EW+G8rPlGL421WuCCTLGf+
c3C7UbWjKme+DhTUm0f3cuegpOug3NryR7Gv376EpQt8oiQMjzbNTQMTeJHipiO48TVOcRqnF5ud
sQ/S9bJY6LtuZKhBnk88ltkJPm8CPZRV1sOUtESDXOTzSyL/CZsDjxP3ApEbJScUfjmcg0WfPrkB
qiXHpLJ2U6904Qc96QISGV8CoTIv4XWrWRfQJu7D1WdsmMfNDkmabFSDRir6hRx1ksw02iwuWyTX
X7v+CpvGXlBXaB3iM3fabiMe2wFCxsjVMPVvw4aUjN+P2IE3KoBXrro5mrdMalRKInfuWBXjy5v+
N/TLRDx1FIBiDekv8Pg+Sp5uF0tSvHlFgF98PlpoJtXPYE+RkGz6PhzGyCrt4284yRAdl8Ygcubb
Fjp9cudahVDdVM3sTCDmPFHNp5g/2AlRYTQLiS5Sq9wyrXMtxSPm5jYzkicSfCnOBkF3vXdmNu40
dhZL2FUmTqxnfchn/zgm403nFskWyZon6OcXm/1F6mQ8nqSKm1v7yjRUgc1fxXxmDNoyE4dj0PxX
Xp6nP2zmux/xQO5TH0A8t0qjbCLYxP9BEnr4ki/nuSuhiPbVhHcbKStm8dPOMH9fZg5LY5CKBGK7
ILi23Q5x3zAsZq+1WNTqEsqkcrlv+oA+fC19ENc9DdCwXAWFjPT5WcNLdNSA7Bj0IWPd4AdK0R/H
JhdmHg+ubECQc9U4zcZhT4Psq8EQ24T7gqAOiz9AaPcHTzvf8ZA5voJmQdUNLf6W7XVANbEzRaob
2eyd21GUkfDffa+WYf/Ze/e//v0F/ry15HJ4fFfzoYegPhxsEzOzQmeKIYPpg8Es+/tfkKpfpEM2
3RXf6MPXdEup5OkBrofB/Dy25t1QXxz1RdSVem3c0JVjEZ8I69NhQCDLO9wWWe4Wj2nC30U0DsZO
ONbGwG0Q1SyLsAMkg5XmFQtVscPoolt8xC+OEa5lulFA18Gqgp0WFKiipCGpD/4qIH3bBwf0qtDf
hq5Qwnug5l4A+Nhq/mUVOgfIEsggNw6JnVdQaiFGB9B9UJqhXvjq39KbmXyaTzoaArbZumxy7k+b
SHlfzti99i7GtGajHdx0mGcYIcZNovmWcX+TxAReUIWGGQun1Qv5mE7qE0DEHYD0hqr0IAXqaEeX
XJL4Cpq3J39Wi6fkYLocqdfONXj5fpOtaJsgDRcmEkceuS7kFNVvUOngirVOZOkkbcDTlmDgpcK5
aJOVfPwADOkJ7/Ifp6bx/QRXzBMbMGmloHl3uWqVqcsNfYhPy8pkAsWZRuz7RkZISzQFt1uaj0hv
mykSM3YMRbkjC4ioYiKrexlAaf/NUzNlWb1D/IBO7oppUntP1RV9KZsvXYAbvuTTl/dq1aRJ6OBF
Q5MQcweW/wGPz9Kl2ra8V4Dbba6C4sxC1Yos16Pu4mbmNBFCW08krOfqzCDNNj/B+ejx8SyUJrVJ
72W0OwPPsLlkAZcpUOzsaop2PBMmOqJd7i0vj/jX06raZkWl6/b+qLYfy3B+1feK8w6PwCuTSKXl
czR8AXMVdfzBmejI3Kh+Yu+wd+3Zt18tab/boU4jGJ0uXhOwQNbo3ggQtpgwh2E9jsJ0KoDXBzze
2ilzeS/PDPaO+R6gBoKzOmw2UMF7jKU2Qq5DtX8k0ea3zgk7L9W04eKCUn67rndc7Sc8a+68Buxv
XCW0KpS6yfrr+MFjL0NJu5gyPIEcHzyLNCrwqP3Bu9pclrpdcTxA4qTwnFL/LbIlel3bvbc78qKb
Q+1UkykyxEw6M1gClxxMeInHo9LkejdnsKLhtA53T6LSa6FjQYsdlf0PAUJ71OviTb425W3NEtZA
sEID/zQAoH/bGO0Kl3ilHWJEuANV4W/6PsgmoA4QtJ+gI5MPgPdfwnlKOwWbXiJsXkw6EnWqlDxR
yXXN705YbsQr7Jqcmdz7KJOU8Hc+oHvqKy04buqygjopjm7wYLyX9Ost8jMY0DRcUfEocBtpiPZC
ChIIGpdpC5zBvmGqJnnvnk+9eIoWjAuLO2GCr9C8XIHOztcUM36TAFaO2lGYG0naaqz4c5Hx4nvQ
HIgkismJ7CkOvoOqX8RMK9UG/PE7+GZ2587Sr9PLtpTY81L3pEFTUZNlsvtl39gpmP/Rd4XhPYZy
Z8kdNOjR8bLeki8/jgpdpnE9muv4ei4IRUKtTONpLcKSH8h83kEtiXSOIDClX2ciLBGReZHhoS7K
JvgJssXOF/x4ZRqXQ1Q6BzX5/Ce4ARA+Wb8SsapXnUCm8ayD4vWHCBenSt3vrkEUag5VM6O9Jt3+
qpz+DQzsoJozD7FYp3sUrIeezOE8qHhOidxul6ZZu9Q9JkIkE9Ub1RXcntTF/rIiVZFgUCmcxJEn
cgg35eYCV35QB97BAm2cYZ3u2Zp32CuWjFq6O6O1K8ZDVw9BgmprmW/xaiZaDkNUCXiG5ihD0jwo
Z1lu6YRqs5TNu9ez5RnVlpri6lAYuYB4MhTvesQLUs6dN2y3QG+QiNBKU2v4HZYNrUtEGK7RQhRe
Lxym33IcGCGaOYb8lmrdhjjU4/MsyjWUiO9p4Kz450RviCCQQH/571ag09lcBoq6W0S/2I+xBGLU
vTLjTIOgonPelnzJ/tQE7UDA1hJbp13am0gPFUJZIvtgvNundidxmHyNxiixWIiUmFwqKkR5ET2i
SqLN7izDClhtXDgiO9BUFi6DltqsT3LYF+v+kF5gGwNZslvi8jqZ9Ew2svANcfmXQ5jwO55GfWJe
7Z61SQz8AFpEQyxYnlaRJ5iDklcuZLyfLzdbzWFqjxj1NWb5QCgtWo2l5Ad8usiehfr8rjQBp/uG
ZSlEf6ewOYJeUWTxkdQUkTOve12GCJBr4NOiqh+KrJjWJX0y6+1eDT9pVoJwRNFcPcxivf9G2p85
l/6oXgxNiOtZns1XA5GdhPgaYOymKR5CAWagYBget0amZN2lwhy9Rk0ryuWO4A2K2+5beTgLNpPT
OMuxdRHNT+CXT+mDsZILr/ZS4l+iAX4zmxCl2N12StA6rAEA++lCCYMeP4DIKVchLV/9P1oG8Sav
NKU0LuN36yz+okzegfs949ZF40Y4iSr8xuaTPR6NdKDaNJcBdDXbbX2eVouGf7E5Kc+SUt0RyYTQ
WNYtF/eXbFHtuq2cvVfbrX0/a0ZAROyFUixrnSvZZUcWSWlhIYSI/4DvfhpE0NiHdV003x872N5Z
C63aCN+fXFheri/64t7v2y5SSgpGG6bAm3FiMdTevIScs7sDiQ5X1/KQSZKazT4SAFIoXmr4utRQ
kuQWXkqfAvhHTN6aQRN3Bvt0TGCUelzdFnmCAgpMmr9fTWa4J/3lIopUz6rIoswmcWCqXzb5PhsY
EyH+eOqT229nNEujwfcD4bgOA67LUjvEq6ywTrJliZhS0E8Wt5Ug0GK2q6xbB9/YVtRLYOTtJbFi
jhKxmrfjaNmicn/u1fcjfsvKB+Uat8n4Eh2xpcKU7dxcUGRropbRJ12xQnQ6rN1rsTc8sX818ScM
khzpfijudePoJIU4MpTMVk3HCPpsg9kB1Mjrhum1osXDnDnAXDzYQ8nOGltRgy1ciaK7uGDVJTwx
aDWrM2eM2OxS4/HTyKLmFEXjyE/dTbWrozjfs3ax1pKlmzfb7apXgWGSrKrh9kwYh97f4SsnJEnm
klnY2k3zetZm5bWvgTfkwuoTMW3w/gurakDhaWg/bQAEjF0wIc1vkgXDx/ysbdxkMxHEDrpOwJ6+
YfwOPIjcG8vL2Y67uV6KLSeXlLPtKvtEedmF9qW+OjA2pe0PuQyBrfdZN+BOBfjoeUBMgeWsOnEH
tba4uNUFjhQXHXRcIOAmbIglf39qBSaa3EkR66Ucd6zEmnYkRvLYFZWkolbqKFK/VV8AzsvY5HUD
oruuXL2WwxIu6DJdv/88Euh3D5vqecT5r5dwTwlz7EPEN0HIEuiNAdhciJNGblTIgM+VowXL9/zH
cpVO+Fo/OHshGimGU7YgVopwTFrYyiINuckvrR++HKSFN7bGpsVD1lmijIqunNrJGbxawxH/sJXJ
r2eS9gSXqMqvuozekUuqkEo0Y2fVkxxL3q8XiQU6ZpIp3sI/5V6Wv2BOy0Y4EQp+31hYoub7CiSL
9/WjX8S278nbpdREyO6dh5FaXmDqFX8HAhpRDnpwYl8JFO1hl/jZSgxKdtmYR6oyaNmicWk2omqY
h7ZjvKKoLXNx8jr50EHM1mPU3pof3n5xBVGUj8nHCJAbcRY+IKyvigWhbdNeS/FQKwOQsGlGZa9I
6WQYYaIeQE9hdzevDKeQ02g5HtTLzhjuQMWDyAVz/TpVeeBfsUPtp1cIFKNyHX0Z7LGAcgXn2AT4
7df2+uhp54v5fcHS18lDV6NQrobWBWGzpfVhz6HJ0OWpakG56bGV44foE54TLe22Cm+mr/u2yn4v
jhDM8xW2XT+ZZ59Fq0k2yXfPw8YrJb/E0yhuewsVFP6N3YCzUUSGaH1jKxoTRX6jL3T1Z4wTC0YD
vS0ZW79dqd0sIRPzz0PD38pZ7QrqIUaLpGAH2pcbXvFrX6BwUa3OFMxTlU485cf6IrFTjp9FWxTD
YN0DnvzwH6068Z0V+dxJ9hrs4/Pn/gGl6oJ+Yo1/jfQnXkxmeMj5OwDROpRt1t8YeisuCy4uCwVE
YZv+DH+2bXixSEnF3dUadA6yFyODiN/dq7TQ01G+rqxOJ6PF0XPOWs0P5URY9XJU5+MRBZHtThWG
kUsdy+9YTxJ0e9fKqZL1amcAhslVoX+CDlR0FM3XiY/9Vss5i4wTAoKa6gBBTsIDoqtf9+0eS4Nw
6oGbUNYPt3vtNStciNuxYy7QMDZNXscVgiq9O0wjMvtR3hUJisRAQoPw/8ALIOnLebyujmOiX55M
esC28KNwgllCTa4VGq8gx7sF9paUEaWA2ygDFAfpElC12Ri0t9Yrye1AWHCUxNyEkuxdZ19j6AWp
j10YOLFZ/TD8+uprxRvAtMHDFgxJpTuHQJCe7KatDbLLAnCAeRLYfUpn5Gt8ySr32rIUXboXhDIY
Q6yM7qlWiH4mGM6lifnoPu6kEsb2Dki/j2yqMVScJMZSJyLJQFc0d7WPAvVHne+NJ4DQmnQrOovk
kbJk+ueIgVVk6EL/oMi0PBVHD3hDkFJy1pOWfWtnvNQa03+pH0pD49Z5Ne63H8XvOou8fvPCEMdL
trb6y/qcIboSsTZ+r/iepam37p6Es7Fz+c4wjlwnd1dNZQVBUj6E+eKDmY1le6INSqfpoWsERpiJ
w9yW/+3+hIPFKiuvIcD0GJp/eN5+FU0A1bMrV6f35aGqwIzNlL/xFtQFgvD+J4nOWHSrtZ6R5ObR
pXmpivAUPgl/+KismX7f+0fhGvTegt5WoQVMcRV5gl34nCcOq9k31nY98UhWOsUXfFvIz5NCkfaD
dkYfT+cUCbMxggy1x8Thja+xYHW91UpxrQkOAqc7trfyy+Yx5VQQK6glglbAA/e3QJ6NpXfSckEK
2gkn8/GtrredLCQXpPhHl7E5Ek/TmSDARpQnr88IuRezlf5MGs/vc3JIWRP1p28vuodckuNTyrac
b95fI+8PV8LKTySSmfpFVQGe9PKeqTvkzp69yN9crdC+i6w4xOxkIMhspRvRJbHD0/MIXj9TEBJt
9wuzOgEp/ndtF3YXm9q1VD67P08qRxSWulu3okHuGapZn9XJDEf8sg22ZYkfxEbrmLVTGRMkMn0E
AkziUX50X+KmAAPvNqHgiZ1h7rtYWYwrTok6lm/YQPBB6vhOVIpZPTptdaO8yjxr2MnGWhz4QWGF
RICwnUWrKr7h26ORQPZT3t5/60NGJQi632nLvMDJZ7mv1W1cOuNVsDfZXEGFFcmeJPpVhpP/CALp
e6i8vY7eUwR4ylw+6GBrh9nSm9l3a82+8SKZLoF/hjxiU8Cqg5LgwDJaUEaYLEdqy2E3xd1rqZXR
Leiy3Jc0pa53Bc9Ypa5irC5ZQl8i6g6zMT2//MQ67NksjQ8Lc92WVxo3D6K5m+o+7/VcM4FDCk0I
FV8G1mEfPZHpLMzvnJj2W+r8xCZeLyNjjWFBXpzTQ9jy2uK4KWA6za+9DtGvngdAgz8u+Ml1So0r
9wCMaN2+suR4TbCJ8DVTX4r6PofupzZkDDiMbYX4pkBQ403leg+TVUOdNY1UrBowu3iM7fsqQJG1
pAxvG9jdg4P+G2eGsDWrNw/49pSkck36t06kT6Y3FNbIAFId5HzlIws24c72wvT3KiRX393hhQAe
70Mcdb+nqYzhoGMJYVZJOe7I3Ynsj+GUd271LjXjL+kVgIGqXXAQxKmux1QoJkw5NydMhOFXGkEA
0RYWR1GcM9xLW0uG3Zz120yfKpVRgGC6hz36Gh0+5bPzvc0todwgKO0cJ9zyXC1SoGALkA3RSJZB
+y+bNipNKitbPjpQpgFEx5gT4iiQUUiqgPFxHQ1EcKu2fW/C/MXVThtM7TDwlSC67utF/S31j17c
XqbcN2bmnIajNWZymRZXZlT5FwoZzPr1rdxTZrG2aopa6rEfGC5L8w1vyf1C4Q38DLHo6CTcYSry
eQsbnZgaUmTGeUtEkeIeNTsxq4i9lr/WaKPm7ab0xjn6oFwNv4M96ofCMxJfp4au+cdTVBLP/P5K
aGmpyzpgfwy3o+CN3cQY7AuO5qs5lbGQbxS2v6PeCRLcEyqjUF3Z9NjFJZ1iDYTZKNUGvyc3S4qt
3JVe+6kYGZO5rJgsVoddXFqwKgawTbKvtv3RRk9tKygrk8czg6PlJg2F6YoGdBlvuEMRW/eFtB2m
7hhBsN2mfJhATqnyzLPNzVvVelr91bEkEtsk1CW0kOHRDzm+BjVhdYGuO4NvdR9B8ar4PLezV5cl
sFjRgMOuhRQkBGMj1TQ6NFZq8MzhjI83EpA7WIP5ZxXpQ0NTWLs63PP6PWjsYrH9CKb7gOVXVcXy
vv0f9HR9H+womHjl2omDpccRdZdDPfdc/wsRlWLM71R4ws5N6MLn+ahzNIctgpuwtwONTyeYEJHm
+sIyt+Uo+GrABHOd5Ehx3RbvSn72fgD1GZwLJ23IWYhUb5DGWtAWN7lXp5joKLY8Ey7Dd2y49NB/
Jox9glo+UKx+MPRaygNRrBdZKGI9uHsWUjVGvbD0IfSmvy+Vtl5xU4ap3CPPHlGpPeIbb9O9K8CY
JVvL8sNkOFg4hblpM0fGFscMAP4YRAu+pGVeZBVNuH5SX5OWbEpo8NwIktoayY1IxuvaCTdYM3my
0l3omr248/3sJxyR1/G4i1rmqHuLgihzyO6rKg72l1sXGjRX2yKBXUIz7jlLsHgwB1pWP8Oguq0e
jNVgEuzDQ1+/V5s0PGnt36DgzM/dsFUJg8MspyaMAq/q/Q/vtaj2IAaDszOjMaeVwRkhN9BSJFWP
zLJ6InnhR/CgeCmFafMi5XLlWfrGl8QYp2JW4+v4DEN0Jf2420yk2KYIAAfNHqXo2GNvA7COZPUW
kJ0PYHyTcQTjryqJeDeyNfEm2kR7PzandqYWgREbZe+BbkuWFNwYPZ3y9de25o7YQdBJoeFIJEXP
BrROo7tVs9sG77JiDnLS+RuyKKvqieHCgcSSiStQaUkzF0bPBUeNBrOzz/PuqMEfIlQzXriGkg7R
WSam7xq05pXOMyny80jYllZolTS4CCyTmjPtJDMfBeh8w0VJi6McNXapxUpe/+m/2VGfVxmoH9fm
ET5i1Pa73bcaE6lDYeprD+1gb9P+/NCiM4mzFMm6YLQ+ZhK3LJ06Vw9DQvbJb/R1Gl0304C/V+qF
lEtvREZJcdEsyb1Fs9KtvgzJ/7ZNaCY7nPSKBnGTrgs7k7Wp+vZWsYTq/F1isM1w/x/SF1E7Cmz6
0LT+C+OE6F6XHPLhOt3fNyfC7hHLO26ui38BblErXeEP48Mm/qD9LUKPs0TKPD9CX/vJzeOr7sED
yU3wZ42c4b1c82/LSxv6kUkIlcbmJa/ImH6Zk2rW5bKPnwi50n2cI2DLdQXso6J3IYAaSuZKF92F
kVaX35hYcuCezZPn74E5pBj2oCWPKtHzjz5omHslOeWjTGGY/cdybwYlRT5r920AoL0fLR0DjyDp
FXPRhtjRFXCIniKq9J2/OTdi1ZieJPjv21ofuXq5t8C5b8aT00JAko5UWLtBaPviBArgTjJMULKL
sIBctdVt3dxu9yD7Gcd3K7n0oT3YuCkdZ4TOy8vy/Y4rw0ihRfdjhO66YMO/qiB1VW/QJxfb9wFV
ibi1X1kfAIr0ejez4fJEpuUuzZ99S6i8M0JJAlAwUr8llBJGayO6t8YaD8QvfQJyNkV08Z62aHYk
nlMI2daereo8RXdoelxajho4k4Z88rDTFSGVc3y1ugqSX6H78rKjp+KhowBtFc8ed3AXNqHBn9JZ
LCwXFISiWsb+HImVsQ3Hslpg4XPqsOkGD9B3WD8cp/fXSkI9hzKt/IjX7sbjlN8KSg0mzaSruk1Q
SIcypgIbVvqXU2OHL4KyPGzob1GSTkqzheJeL91S9YDIxEHmecF+/xaUr/nhjLvJOHTHYo/qnqWk
D+gDGlLVJzAa/l97/E/sfZsvoB0kMmeO4D351JhcI4QZFj1yI4mdBUEfQYQTXkc9nKP2TuK23KGc
pKDDGsZ9lN24pwlFa1lOl+fTKMLe5eOrRPsGm2ytopa/C2uRJ34KBef6DFzwUepXywN4302loeR6
PlMdtH4UpNK2QnGT941UW5d1wNtj44DyXzmKMzohFpeC02IELYsuTlq6uVHjZ1LfO4YEg7iA3FRC
ceRKXaU7lxB3ZEGRjI0mmAj7YBteoYLROpUpunziA7DFqSJtVngEq6psVyGJ3cUrgysdt8nXmYGw
v5Gr73GNnTUS2RsOOsGDNs446Wnhi98ADa8Ee8LVsA5sDWYGCf38KFBOIUyhXyLwZMh9lqdPRUtA
MvFMnxNwR0gW0csguGmMip3b5RPKXwRhOKG5+YxBA8YenP2zaM7O98j6JirF3gkvRTGevm+lYxR0
OGhv7p3YIssLv0Clj0sfHmHmLEeltwwAaMa/v1W0tweV4dI7AMTSJiypIgq7IscI4bKLVjlU2Dde
JknIojTrABX6HY5trA/UcO+idPt2mLI+0JOgfddSXFgJIJO38nQURlgfcv/sCTJZyP8jAh0uVOfG
ZvYMQUfS+O6s0Xj7hPR2B7MAOwZHEqoH+ckBxXFp36mXYKwuV+7UmA3PPQHlCwcAiO7HKb/Jj+BD
6WhHng347vRXDtBNAcZx5uH7yOazEi7uPnHeDIW5EXcPmPoiXHRMz5fCtJiwtjiU+QJR3VmspLav
D/WOqNJx2Uavo7ljkmHqUkll95zYW1A07/AW+eAUwVOZWnotuojVEB8jCFk+Z+i7rQqhhrKjXILT
tz5WPcbPt8YImDcSyMuMJng4o6yp9F8HOwcNrkhbl4y0H4/X6BjsbCMCpvE9GDjWC/dS70t1jr6C
k9sOwh3mwHCWASa7+L//T7DWRhimSdjCRqYSutCX+aDuwHmRkCbb7qzOXBMAG87iY79KGdStJpkz
r3DCVxJwsSQHuh5jdLsgc7q8PQmmLBRq3lqEaoq0DU2fU1HcZeIQIvhECdyXKwd9+ic8QiPP52th
l1DTgv6FLu2nnDRaIKTQJIKHL03OTx2yrfZbGhtg7AIG0Oo5cDJyOtHqlwUVUO8FHxuGXT8LBP98
xZMNWTAkh5wMTfrp1/RxAsyu9/rfXM4Du3y2wSzdMFD/k2nHU9QRncJ3AtR92pDtPS0ZFrGM317T
0DlCBGSpH5vhkFWMFvHWsS6OtmiLcXz4XU1kbCJOUh3PQebJfB81lCsvXhCv6SuHTuJflhS3w0TP
qNXqHEeuNOtjWO/0H7vwGEaZFza0a0V0tvpzHwOqW8Qhh1Cyk0WlT/0VSPV+A8lE4C42YiQ0hu5/
cGgp+0suokX9uT99wry6s2avacUfov4FEze54DOw9CuuEfrvUeQLWg45qJP6gavMYeAFiBqwoP1J
MDrLKdm9ZHLg+grVc7p18Zw0a7csYsVuT9a45Y7xTSpxh6pGHzEK/iu0rxqUxrrvY3PDcv97pE7i
6qoSw0IWWcYKIlHfdLhjrmbZTTUwxhSqHNbhBH/p6W7GscXqkZLUOMOW4RgyYfvx1PSr7AFfKhZu
q/BDaLgvdrxql5HvkYQ2yQjKHw97TI4ddQRfLSxVgnjQ8JXB8yldERW3EF8LN2/HqKclWMT4z8+/
kG/eXq0PLWlwa+WRCWI2oZMxD92Nc6WHO4Bp0JCsHy36qJ0Uy7YIpdQG1PSwg0kKK46bN/1DaO2Y
bIei4SUxrJ9SVqSMr6HPzriG/lhaxPlRguBleyX7Bj/PQd8rfkGmM6PEaQB1bwtFLOzXxsXmNAhW
zjIxt0sYcIBzfq0APhrapRVDyQLtNGz8xOx0Ra5TXnM/BVq25K+Qyn/EWJSwVUBhOT/A2HgNVMPI
czmuUrO1geucbwH6KROcHmAbsso617TZI+YVZaoglgPecNDJg2ZfbWeuqYDodEHsGNktUUxgX4bg
cKl7nZxfO2pH4CFhkj66TvF8HSCWNWAIJd4jLqSR89dp3141iK36AB1uFACebWnoEiSHGgOjn8La
Ykr55iiEXrABCOZ6O8vsMBCwcXVYr1ihctBENNgD4dWZTGYS7vf5UNj/0+aL6PrWcyK+CIkAZDBZ
0QNyk8Ug2ex99HzFX0xz2L/45GKsoAaVh33BrteD0e5tv67G7WjxdLqer1aDWhvhj23YEBYj+lil
3ur7fMU5yGMXWApNjaAqZO6K3+/MJRHYxYTOfhcBmR28cBSN5jBU6cI+AEHMyd5lf19RNkYChvxR
NVjjsrCdVM7I+3oXHo3d4pOw7afofaRrMHUCBCXk8KAVhn44qwJZ4cPaR0MSLN1PRApMefW8gOsc
G1ZzxB58lUlZJviEWno0bX/hSwkFCtZEEH3l6geD8leuI4pODG+uwsrxZ9QWxNSUA823xODKpuTZ
wnqLzN/9KbsE/s6gWirLFHfhQpWG5/rreE6wBRBNTm/XN7Xgm+s6BE9JnhXUxhM8vFp0BI/PzKHL
sxvD7v1pdIQTFvmSrDrhFl0ety19e3z8+L/CL5d2VwUu2YXiPHcpRBNRN0V+7KeRPgeTml4TTjiD
3TOsqnQbfdL60WOFEWokXKtN7Xw9WG+TY1Rlleaavzh/A+Co79lLkz+CVulS+G9pFG7S0y5THSt2
8qUevYrBLJGULw1YN6JJcm2XjUydUMr32yXjmVT1zn1YPc5Ll2v/U/YfhBHFjyatkke+a1ABCHTP
/zSZrOGI29iRIwJxwubYHB6m5G8UIoseN7Z/eXrXhNHnw2ZUTgjnViITs6otnMicLYd65Dme0eCh
r7vm+puysLBPiWDiG0FFDNmswlGHTyDcGsfbG2syiJGTl/QTg9h7ZVZFA8YYOFjXOah75p4DWwN7
G/F7+Gxxdy3X/zlvHDsyut0OKa+mrefKsJ0tvkKvOdMNwglHclMcpBoYE8HT8LUyJMZhgqjSxK08
Ne0uYSbrY0ed7bTKfDNlzghmd/7yWUA0Q8MNJGYaHO7FWBd6zSpisB32Fcyxc5Dlso0Pg2XzXSnF
4kzJnM26UsugAhsOHiFSCQZN5Dk1TEsFkhGc18XQhUwQG69Gsf/aSdHtDBxfrwG5Hkify/k8iVrL
CKcW3EM1d1hEm4ie2+7bWBhLpk9YhFKgGnu/wBE0pasMnbygehhV/3CIUyCaA0oJ1D1+gRlN1vUI
qTPhHE00OebWBbf7/KHcR2VlXiKbL4FHpxDL4USjr06h529tRyybaiRIwbAtIKa8laxck+hcSFaV
ZxMuZjw4IIknG4CsSCxGSL7RDLgTwzI4wtDkSa7ZtcL0thdg6Edsjz7s/Oz0hG1e+KRIgQ4+m86S
HAalshoZjtNGVZA57ZSa07chJJxOmWsIur9y2Nu4ow50m7CtkhBC8g5DDpbOsT4e93mj78StB0mM
XjHnA3Qjmh1T+oAD5h/DDxZ2H/2Uon/i1jgcEnTMYMJrXsIeFWJ5ldN0UPbzSbBgRMPqa8vL1JmW
ifCyhuJ7noED1SoFou5ZXOpCTZ8gebtEe6+ubOZ3ReETu60oVg6xptqTR6/EERSZf5L79S3t8vE2
k1veiLoWz4wG3Bb35klKqsmndz8+ML3jQWNfJ6ZdqvaRJ7OH6ZHSTb0bmaOpd6XL/LnyYVE8yCV0
jGcvgIzIbK0CJaJyQvLBfT+cmXolliiBNbvrnaYSw15hQ1ahGyx1STqJii0hr2w+RTHx10RdEF3B
Vmk/IbqeINwAhsiU3MBDw+zJUY17VbwBZsJRJkT2HbkZ3fDjxCsTGMrEzYdPx5XQyyhZKZjKafhK
WytQ0YyWLWMOEUzOrX1O2q+piT7OdJJViRzUiBg/wHpl+C5LygZyVLowjKzGsogC922wSSTtRFvC
BdOm9ywOtQaG8rzsomtQ1G7TKUvDdH+CmQvQfCHLr8g9zlty1ybfSyxYaJZEP7LhgpTKgqQU595X
J0eZEhv/i+jg+FmUw21EZepzpswjdj4ugo7wM9tATPDGqd/dVD1Aie8H/JLWczteZXPvz1QBID0r
4beJpVfN7KgSHJL/8zZvVTmv7wEs0kbodIRKE6ziKI3kDraWMT+gQGsoJNHecW8RsR05PEWrqU+2
fec4if5hTgKGqXJeztwydkn3D49edcXE2kYdKIblsoSR1Ycup8xx1RAlLBGrfK8XvKj6jj1MfMaG
EzChJtl7wGGSdTabyT3iuLvMyDfTUJO5iQajZIBFehO/ooz4fmGNwUlv5bKvBNZcghcRgihlDdJK
EeGF77vsiZG6u5Cq2oFgKRgezFCqp0iF7UOMtKKBK+LKywCiklPMkPjcDcYOl0shvqyGVze78L+E
SUY2gVAhtsE5jHYHDd7ZM6pznm5C4qsgA+m7vejHdCNSHAnsXo/7Jxclovy9n31QMbLX77UXd5Qi
rCHY4RBxV0ouKnH71eAe6oqE0oHgklDD22vfmZIT7MC4Ze5tyr8ODItRq1NI9MhZLYSc379El9Y9
sEMMcdAhpXVliaU94IdsqahWLqW2plbJUg2bZmnxSwUHypfCyIMG2ZLkqAOWymcchLwovlqIYgA7
YPMhmSQq+FfUTvutGYVopACypsfwiPShsUf6mVM2S/UI7J2D+vaHnElItwN6hNYe35fGcMliuzx6
sa7yduq9nw48oBCLoAKGuxm1gBzI/E8gIbLYk1eXwdWDlPXLNYET10KMtZDrNtKHpqqHA5I83s++
DvInTKTVCX5mmWLX37GV3wf7GfKX+6tWTWuGUE+8doFngC6kuFnFz3VNQT8GLnd3pmwAHH9JZlpF
6BytO03/8Pbj1+p+R1U4+Ey6c1MIbvAS2u/hfccDQqJ/XBdXRotAUKhAm3tN7xlKxX9zFbvyh9dN
PiJ9VPAw0cKcafyO0y1casJnxi8dEs5oml7vFHs1pw7buCCHgqh+sOHRxE67KJ6ysak4UANYaM5G
CvhTWS3k6kMFmJfmr2U1BjVLEwmIjhd32b3rHcVKXInKplVizDlX3plSDSaDO8D/dy4VkKogpyyB
HyItAd4BZGEykDZzWGDVYUeK1N3oYi6tou8oMzt9aMeS3yIs9aeH5ZmKewJNu4vkxN/R1yoMo1ts
SP80py7IvExlEd/X5Gd1pLpElMiKMM80z5WNvcIKRzKyJ5uAJvTFBDo0MtEVGdL+JDpGJlj3z+VJ
KEvKn8q8Cz+tTcenJWH21XRDEvM02fQiESUgcIxucdh5rDEpVyDZJRuHBK8J3JFs2ed9I8lsBCZd
tvOmYFBR1AMNM0MLsqCUzee6p5WSJ88YDdwVpTPHvhFAtiAIhTdm9Kg07pT64MASk18FtCLdPX+3
gXNSnFx0vCB99ncr6OlC5Vatq0kyU6xedlLVNfR1vh/BIjNckhpXY6j3gkASmPsXd/OPEFF1b+JK
V9561CXKklFMa7w3Oxu7snZ7rz0wmZvNiU6ueay0/VSXA/sJ4fsAlT0lp8rkhcOtdbAreB4mOkK0
BYxP2BZbR0g0QMpfUrhif6UG1uerUJ+D9ICMuAGUYYJRZm5ICUNEyKh8Hz/HM1HnFd16+U73RTle
IO0KVjWmF7BjuMrQYaZBF50/z3BYv1GpJJGsS0MXtTX5LeymeKse8Pxy6NFDVm/JdZCoYm88SvME
CEjS6UWsAzR9ELsxRLmXrX1sSIY5ObIyzFDjxHXQo8bWvilRUnvPrIuDmiL1aau++4/A9qZTxqsF
BVCAJttCkdWMt3efzOk2FNMw6YkNu3opgFCESkjMtOvj6PZ9uVRHd2j3KvaI2gB5JLheTSdGpOwN
iJx72SIPEIcfEpl+LvUOu31D2NkNHPBCDxPjtE1XCSpm3kXK4My011+pCiltzvq9FDn/Jf4FLJiR
hCxdWTx978Fxz1DiXUiWTBOl/M6rPhV6Hs4ERNJlk8xW13i7hoO8mBcrVz78FggGf+OWYey+fP7w
Wa3YXIRvXA4S4z/VAxlLTNL47iV5+FpeCRmHLGN2vHG8rb77iBYBGFXU9TPDQqcYz4cpa6oK3VoY
8Xe3Rx4v5YRI+zbNoMJGLZKdm5Wlxe2MiLDkSbhqEsg3sNmMUauOBuCZju+5Jbt6W/BiBsQL7k1v
sUBLbZHvxfoqPgvXrmtKenGUDMEhVk3za8MNW6q7aMbTjJp2XeOsP0dYWijMoKvwTQQKNgyCmQT7
1Ok7o8ACHnoCUHxjQsvJSSRS/q6GI/jVg+IFoRRUod23BOE4fVBe7oWzOyZbvx5JY+ceVqkHWdV/
sOpsTtzDX0L7ctzLzsuA16r0S012rOXDrvuD0ztiF8xngo3PQKSJPnn2vN4OFvLU56AE/xk1UE4X
cLq98WWUmvSq/S6y8dg11HOb9yjTZ+Or5IKHYtjcrbNjt7ON5Et2uefXrKEBpk8KXK6tqwsEhV7O
heKsMb5FXjTY3iBCRoLCq3N6In6V6iAwGFXc75oNUM1ZCfIAASTu/09c7UG+WwlabyVETtxuYwGV
awtxkpSiHuqpxA9pUtqKoTXqk95yIldCr/rByGq+0wBKazV+hL0teiee0+pFX5yDm+iVyFmzKhnm
z4j1a7pqflY/mNRnHrYzEwPvD1ik7LuUlAjctgKdA5smWxZ7+yhYVsUqKqxKmARXkiOgKIL75dGc
9C6MdfryPSkj67Y/qUeuSbPoqyt6K28VLqnoZdkcHaWWgS5BFlqaITqGypDaTifY7Ve8OEfB8zrx
17yIVqN2x72klV1q2XwD3n6/a/z/xdTQ/UBDxSaBITF6cpJwUgTyu0mUblKeEGbIB8CJ4X7bK7bz
WVUbWOwVauL1yEdVtXiyGNWZWgOE7aOnTGZvZfcpXq05fJ5ioCPt4MtT21XRyDabEllmFVOcfUbD
qd2WvjjUDkxJ/ogf7k2UM1EfqBzEmhlZJsm/ulwlWRnwX0GIgRkx1Y8D1HQTMo2J5fO+uIjO664H
dCguzVv8YbLA0uFAeomP0W1MivjOuSdCDQxO8awizQE4MjplWUs3+plTIm7AfNQiwcX9vhvtS3T4
TIPYiMI9O2C6/r3MzCUt/fZfyFvDX24BR+aayqQi/Fyc8ti8N2XUA+WOmc7AI7fgyR8ke+GBXkL3
Wl3+r+PVJqEwDtB3Qbg8j4QnawQ2S7sqQTLsW5hkkyhd2ggexTva3jLckFJ1gkJkKzltGTK6eDXB
IGXfYcZ0JaibLKEFlS/SjlHOZhPm25v5IotJR/LCxsA6TxcqR7e44U1vbwvJ92Y5anhwQ0GBily5
GbqsUkPwq9eKUxT95whISSsE3SerMJivRfG7nncSDEoXUicshYyocOyip627JWvu1jzNQSJMV3iE
mzUHq7i82FDtF+PNY59LpL8qeo3NO3KUR2VLaRo+aZFQEBKKjc0pa4hCz5rwEi/PF1eEsItC1e2J
Eb5rlX/JeXNOLqdV+ekHCFTrPrJE3W9R52JZ7sXr5jD5TXSliSooUK0lmFC71n6aSv6klJz5a3S2
/k4sNMlPKRRvJMkGre9DFbtU6cH04MSy6klF1lkEJMR9jX358cDkhBVXP8Nj7kDrhqpm+sUkiA26
vpFW7gWsuADP2muji8N0Uua8qFYsO5XRFhVbJq3A1OiBmtoIG+deNPqEEap0QxC1gGa6Xx/6mTI8
nuhxUybVVCVlK25ZL007PTR83J/buOjyaGcUDb3fr9rI0pUum5zVl7ZKS6YxB2cQTLKsiHfJJ0DZ
i1KQ04yFqqnFo0ZjrhlyYBOJv+HrdGA8aa6M/hrVaLpHG5GRAirjAkRNxCyP5QtKv6o37NlQ1qST
vpyYkp8Li9jCR4C2l0EvS1JTkSPI9IXnbcftC2kOxhfUr3KqSkL3WaU11zhQg9UyKBh5QUJHzb7K
I7T+QUrqG7+WxGSf35+HPc4TnQQaXpSlc3E0pYmzQ6etaI2JIEK+sx3NmeRNrXRmXk2YAe/D5sk2
ZCTZMJ8mQO0kPksADPj4c6rp8Nn4TFblLREye8Iy5ObRpVWPiMyUp82zxFJLqW7wjS4yw+L13MYf
FZ0ElWQkFzOje6b8nqktHI5+na4uY9eqmShsfl2Bbifw2zhrRYd+RNJ3+vskf02diOGVdgl14KKi
PvJITP7zVgJ7tK7WWoKJg0112LzpBK/GA7T6cS0c30lc32rbbfRsTcfAr6vYf/636yV73s5LNpbg
Nx6Pcd+h2rwCZ4WBBhxr6aKkLVjqRlk9u+8+s9EuAq3Bpsgo5wbeNSw9Pg7u0p1pS8eVNdyeNP0S
AIMOjwzLlz3ryzeOUoQYUvdRdViQjIH4VCV9QkeBb5sAUFRj1q8IIqxL93+z29tj1RsMT5zCeOJO
sMl3hyjWi+nXUtGo6Q2g6JzpZZSxViLODARcg4UKKJaWRpJNo8G1sWm9DuVuBoeCiZFHIiwwalhv
4IA41msIIKLfO/v1SRNcqm8QJy7s8SmuQc2zSxjrVSuSl6YtnLw9RxTMiv3ge9OsXR0kkFBxC7dE
wStSGnVFNu8B+1MeC2aS+yv+kJD665b59ojNrpY6JNnR5QmWwGIzSFybvyYUFWph4FCAHxh/FhkA
WbijoMSskzy2StOOLgKFhsy7V8wYkrWIwJvHbDL1aeBItFhE5AkCd77JjMXfu0qaFIfALlp5UNQ7
/cmFfDv9Xw7lV591C/KC5SLSh9QLSdcyIIrg2MLKyDOCKOGcHec77ccSFbiXqtYue5QUHP/ChVD0
FSB8aVKKWDS5depEZkE26GqpevHps+jUInd2V8Uiz/IOcbiBM2vS7C0Tv/eQ7yJcB9G2P/bnn3tq
/nFbATQtN9FXXI9fE0r1DnOv5GWDSGffN/3du9YB1xcqGF+S4i97JHv1nf0QmWb0yQ8YsUVZKu51
KvC3fqBhEYsYH5i5u4hnSknPAeVd4zNf8dRno+sV/zJkzcqEy/B0vOSW0OC9/gilWXobeligZe2K
/9YfVWDIPOwDYtsLzJSU3M/5KWyDrb1GFub6aQqTdorxRHtCCGbde0zu5tfbQOOFxAScUctbyppT
5ctfRQCTQuwGdJeHb72Da7+ifgKueZfkXTGdjfzH0zWq8BG4xbllgGPRork7qwb/elbKJZ7zmc3y
KK2aT3Hrb9fnZHc3PwpKyfJ+EtX7tGGiZXHdxF8NmZwCp1h89YjiNtdOSowK1Wn9tRvclTwISfsG
CHLKcVe5isVseUbtwlkpIV7D9RMhTGfDnz8lhj2TcQECySPXaRvDQMpMBKffFwpJUlTzojv0iyEB
PFhR6RBYMcn2no/dwBlme3KgdKFy82PszcJpNLndiATGEU9IDCLJdiwo+gcIs8sIIc4kU9ANoC0z
UDMZ2eVYm0ByM6eZ28gSR9l3IUiNbUTMPGrUuSpBLGbZGmh9G6ljHHeRLLi9yfQ1LfHbycjDlL0C
GqX+CggVhWUHrWcZMPYhDQLO9Ot9M16+pc/vuHm74teagAFjuhL9xnp4KaXmt5f1X0C3ByZqMD6K
RWSnROpzgKI5Pf3nx/9tvHiHo6aGiMcTrPSn9igmH7zBe5XnNIySUrYpyzYuPTqFcGNYfeVvyQf/
NG5xomO9FWfFnqC19OWY2M05LXJd7wNLPeumSFU3axpqhppoCH5+byPebuKMOd9y023oo4NFXeya
TVfJIj2AOZpE4oE7GjITPr/JQkgi9L5ozh2uAWDzStI9te3D1WWsO7OZK2HR78po+7Kl69z1m4jy
wqPTkRXfNf8VCOnwK0P0BdiHPoZSQQyaSOg5klfeAsAEWihL41d3ufawxYSkhYLCaUfA7SzHTcx3
fNn33tks1tUD3wiqS9C/ypzNYQdQ9O/m3IplzaqYA24OJCeycSeTde7/KkWo6I7ipisb/W8H8Gv7
PkdbwOvOFxQO9z/SCeUsXH8RB0wiioWtDFjeTjPrvL0XOPMHiP1dfTBZR5pqeJ350nSXsVhy6ZBt
SMD7yQuqPfmd0lkfmVihrTKAxgOuBoIoBzUtKK5aYuWugl1jFidXh7P0PJPqXRhL47G1n+2anrh0
jjT/Sk9A29adqNFHO7qsuplilP/JyWS72z5ldmY0yQmEjzY0cHn2PnTU8w73YblL0Zvf54B9xRgY
lt7iSldy/wdl4iPV/8iPVKYJX2RGFldnPPK6XF7T3qxephRYfMxPQxlL4hud0CXsffIe17yGZE3N
plqVlwskTjNDWIMfhMK+lHphJ0drR/4RyHMBpBww65ZqOaXutPwSvQmK0ByN+LT2TVb2Qt6t+znx
Y+t/m1cBF6j5RndNUbhWP64eFIVkSuVsSPJkAVXt3oa6Wxyqr+CQiQUtWo2ckSVOIvbIHfiFQRBs
wBibsV50z877AvlrmMr2huoAH17glHa3xJ8aUDUK/RmuSdHzYJh+oxK8vuvNb3z3ttTgL0OyMsiT
2TFU2bfSHS7KW+LDfyv6hPJHpdtDs5Z6y9mEIyYlOM0+wbYopODqQc0MUmNUBY6q/IUYKDq2WUsQ
n7ojrUMxciteY0Q88TJ3ELYi27kzqAKrFAmYuUWyHmnCYHCl5F6EpkhSNY1TGdvCN6fQfnE3ftEt
bNWW6O4GWxQTp9jPFvJIvWnRUGDaeUcW1flQigbEYUWWv1bJcvlTGNcSoLhERhBgdYLE/RzKasBe
gupbN9v+pTOBPJspwztrw1WpzHzrTppm2XVgtSrpUL733qNRwRou5AvXcNixur4IH7UsLBuzFhpB
EQJ35tn8pbZj6R5Aw1JAKWM1QcI0uWuFJ75eSU4MPQPNyLqaJc2WPTgkFrb+qcF29SsPp3qAj1OX
5Fa7QYmTxTL6E3wloWe845YfImouiO87b8JXRBZhMZFKHeIl8MMl9nIxgERwk2EwxscQOMNw9B2S
kLucCJiqgfEb8cWba+dlrq6DKRTZbq/MEkKQeWel7Momhw6c3keG2nItpvVP1n457k83v/0lbfr1
i9dE2c6cEoVVQkSsx/4m19vQQ2dhNNJEe6DY2sWKyrmFXPI/taVyKgsugzXGjWY6X4oddlBjpGk1
15MlynZTsczs4MUJfOp5U6hNa4sYc+mt+VaAoeKRU93k6YlR/pq2nsl936vEV44z3igO7Q9Dquny
HJ33UhxY5FiGXTZFHUdNkzBHBvv1JvgSmSCnK3tluhVXvATyX91ln4FAgQkm+2792PdY9ahlsKQU
nd+FK617TPxumxp+yIAgMMv02XruxwF9r/3ALA/URXhtpmL1rrbH0jD4tB9clSxL3wYEAM3AoGd6
dRq5gaGa3aNIZpg65Z73MCODQP/Q9avrZIaJS9VfPwzcKSWRrE86DyVHHwXrkt7ZrvqC2FDslXE5
VQJqNDePuXuCc2GqDUgC9jk1mSgJHgACu38kPHy9NtCgOsHdZD69aU2tqTn/c+QOc+5W+crFhuiR
XiccfHnc72PCBZc2uSBGfdbBSBPVp/8wgcyyRwdmAg6ZqCshXWMp5DGenxsEH/6kVWYwONRysg+4
7uMGqETBK55V0uUgdj3GZGbEqfhb/BCw4LJKwAin5O8B4Awgu8xYAlM005RWobiqJKH5gCaOyiGM
6LBhKA1uNtXnpHvYWvNngut+49HJAasah8KZQ5/ZdlPmI8Uz9aK/yjg6dWQ9OTpy8Z07vlP0nU4L
xafSRynjgeLKsQ2fCgwNGSSxEpwKOwxSi9pADUgRvDCuUbY7FEeVHDeH2DgRWQIdqgzfjXJZNPtx
IDPWGQgVJOZbCJilfXwFE+iwXkmbEaYOMpgeovZLhguxDWU/9OepBH7bM0Mww2rxxOvsF5LbaZf4
AU3ewYXpo7+2lmaiOw/C7/kde8+dZbj6Y3f3vRTkIXA2goHuDA9+EuywAds5DtYbbeeIQoUp3gJE
ACOcRYzLGPV197yU5pVeg/gFvzsg8DQr5M95XW5jX/wFLunQSIuAR0VxwnXC24mbC6/0B7E+PYxv
hOThlVEf6AWjSppLsKByXOqPUjxztp5LZTnAk/6J+jOKIfpl7I408vgG5/NvUOJXBqxE5SL07Eqi
LF961tJnxE/pTnFSM8JGeNofPKm6Xz/bYAN5Gsu3YsVRPM276s8+ARfHxq5fos172nSAyhO6wmno
0KN02VLRr4GwFt6afNTQRhSuMLwiqwtXrwF6FK4nOKOt8T/y1c4BDPJxuIsRaJOe4ku65I2bDgN0
r9wESJT7vpr3VYSGEOWG4MM52Oljc9NjETnmmSqbiM00NnVGOItLje31YVvNg4zMX6H/PivqjRUo
Bx0Pq6PsOkSk3zunbaax0Zh0LgxhLOUq+iS+l5WalGkFzIsunJ6Gh5MsztQQ5zYfmfRq0uuyyvVQ
X8IqUcpb0rN+4rKw5fa7xaILu91DVlf0/3aRkt1RKYEaD9vkrkX2lCvcoXt+rlOwk2HIfU/rCNCp
GQTQbqODKq+gf8u40hJohyILLHgoBCXxpo5DH91cBpRmj3x1iV2EcwSaxYoThXe9pO8/r3CS41hK
SpzXuxF/Jn6g/ddUQVHhv3H5mXFMyTqxxHE7P8FWBbjB+u+ijejrtmr++kLeko2VsVrHkoFUO0Fd
wCT4Mcg2TwOXS4Awsh5J81aCnEDzLv0olltVsQx5ucJ0GmK+KOqQbcrEnSTz7Heycz7/K7m6q7Q2
lA6Q++doFA+9oY7Bj/oHZ78LCaTkPwOnIMKo+K/Ltj/U0OsXc3FtwQgVCs81Vro+OL9mzgxKfvE7
lfPQtgoiFSLTd+W4WuC/q3NlLSDqVLv5IWHPJ7XyfZTeAH+/Vyr0M/NGdb6Md2+5Lw+rf4s58cnA
d9WYq8VpjEjKyqwT/CYMk+V+gqwe2bbuS5U2UyU8GknOMYEqf+YckzSQd0RnohMo5D5k6+kjUyWD
+px9fOccEkcc34W5daOmkLO1ife9NEqXA8/0Dcc8ItlB5dC0RTQy5iWlRPwhnSANBap7Aa8vMw1E
PsGPa0cgkxskhuwo5mYJeWehLXVN3vQN3L1sYGuG9hJvkKsvhap9z7W8WjxlZPISxP9HsoAbWjTQ
ZBvIRDUert8xTIEkDTY6thVtSAImQIW54/x33JxJICg+na79+EOTBYbgcqRPUHy2fk2QsbOt52D4
C16DRFr4pomYrXorDROUQAZR1KekKFNMwht77fzrzH81XflrDOhGBvMfzpKoI2MH2olTcQI7b6W4
kDY9M9QwRETBm3jdF5r6ne5EcsmVOgR5jCjVzslXJuGtSBy+3Wg/7ppNzGG0/BvjiNEFTEf6uK9n
BXt9C0/lFdqBEZ/qHUee3Djwe5tS2AvnRahCpv1TT2+eaY8kQO6qDmnWtCZSjoRD/c5SaDuZvfaQ
8hOz+LsVGK+N5kBUPkNn6AEACB3stqlj/t6L3NrNftV3u2hxzUDZc795oWTWO2f04CN6STQ5IQ5r
Zusrx8kc63hMDRwmZbuaPkAnupfd23gg7HjiFdF/4koqfyeKG8k/xE+ZMRB34FKrcAmS0o6C07bK
3D+pu32tfBXmveoeUS5A9R6pqeumlozXJsvBR5xf0W9nVI7zEQX3T87GgVM206IHJ4nbTWjQ5O7N
GtzmoDxRZaF6K+kyZyy4gVx1gW9HtzFixbmFu4LcVfpWz9NINI4Z2QI9QBcLjxKH/nEabBgF8sXy
229flV7uvVJLo8WgEsdBFBDnsHo4e5lNX8/SIjyb5sCP30cOzdL8d4//uBLq5whCLbKNuFoPYq8x
OQikREs4cPp2A1gHPOxJGA6rusq3bConScecz4XyfojnOFVTyBqlr8v1SW7CS8cqyJHgtFfuCN0j
R0jsoOQ8uDyeEELl9XROaBVohI9R6FzpHQB7gU/rl/vdxWe8/N+ZSfipJ6BRsIZvGcqjpMrTc1jV
WrLToNJjrIssndfGJZa32IrdErNGHfLNV86gbLxA0sRSDv1QnccJTg861NRxxqSfaO2k3bYO7j7O
+C/Q2ujra7mu2emenVatWeC1INd8aAnFaoJaQVlmVU9mPlxBWdAcMWknRIUJjgXsRfIQiDv4qY1f
uKDS0lMi052HSREv9BjzCa/vCJTCEsZZ2Z5ljpFt6wG8k4Mt4eZEL0VI1OKigtwp7d/EPe3R/BsQ
/BQrRQ0Dm3s1bbbyRuJeZHd6ItYYrE0MuhMx1wnYQvQweI5T5Iv0E5ffyDF1bGssra+vjriXYfXy
8H1KPBzDvkvmQIzPm7WIfUM26vBAVLopBBdAkqOecS5PDokJmwu6E3qblM0M73UKRd4JthQRKIUo
MrOXaQqJnZWOAhCXqZ7cuEiX2zSWGSatbCR+UdI1xI35I9qkwvF2iaDDJHF6b6Mz9qqAB4/iCCdc
iKIWhP09++GdiDHR0hX3Z+3mEdicj0iHqBF+Ly4ORlWXaoc40UKzGx1A00tS9cWui6oTehOKKexN
uE1qFEpu2joD/8hk0UGiVIvWuiUNsuGOYGTB2jjKeuuu9oxTL+oRsALJCrU/MZ8gxprheqYv05Os
ZT0ZnvyvP/mWg4CFB/Pha5TGbS9HjZfS4Ys4vcSwIWkgfto2gqmba8C+x1VBjKR1UNk39r8V857h
h5fCd4kToyKEhc77yWGi/YM6jeuSrTdW/1cpcWcKTiBq/yLJSooqpRn6PdfcnBVJR9Sa/UEWBHZA
SZbFvdRYUzmdPV4IijIIn0MjJSfghlq1ffEnxV4TIEvbd56ucPpBHaciljbNzDIMD7z0O6feQuqO
YUtLdl6BnA9vBOeAdmUzfRzwOciEAg6g5KHx6hfeRtVgqLYd9wkUVjj5wOfviqBhhNyWDZUUfE8W
hIvdqDpn+yY9trqu4Aa4iI+G3uAEyiwMaYwtuWex8DEtLvhK5X19o8pMKkkhBFs3/lLWhDGhi/hf
3h9tKHXt+E7MhQBSZ/sGucUJoMAglqPjtCQahlWC7lCwgc0rjoTtg6Cce7SmYiqEM7nnhytnw6N5
DaadtWdQmkI87HqFNfQSzJCG8FAKN7qy0+ZXJvgdDA7CPEtiYihV6gCCecpRvl/VB26prujfB5NU
+7VPVH+lEQGwv6GuThZWPem1T0fufimdm7WCYvg0wmX6jDO7VJ4OJKQ1JecoB5NC7mhGgw0SuyRI
KWsU68xO8zAyqMYgUU5rIdP+nygozn4U2i+XZ3IVVo//fY6M/79je/QjjrCWeKN3s+z/EmF3b5/z
R8r1WCxH7sFmMF1GWXS+taQ6TmhflNxVaFKldLEbTtwq8Mkd7FzjOTxm6uVtvGrU/XoTmVwGsKGw
lf0wJvevtHjWPjm2+maMNAfl6ZjTyxHF2YOwGAp9PvmgaBz9I19ngGHh+75hQwxad/zUYHgIoA00
k/kx54fjVzoTIWQDXsotfkX+DUoKFpyVSJ/wIq74f97+bJOBjdekGZpcCvgJ5a6vTNH8pf0bdLi6
2w4aeFm0sjLCBkdvrhaTeY9TZI7dAaj7s1rMwPRqo5GcO1+lhC/S97kvzUNZ+q+uemNJ/2BnNd7H
8t+2Eia3uccSZhEcQSdCSzzLiComP9GhUWzDXSGl4T54Nw3NX+T1bJumucrANI0yhXZDHEc1Ck0H
W/c0Eio6GEX/1RPhJLn1u6TIiUiprOrnFV4bk7LR3KRGN6JCsGx3lMFUvZeqP25gEUO2WbEvfID3
r5cQ9Ilr8WtjIDO21SJPpwPrTqJGA3hHYCkHN8m8F9uuAOezvyjHZlGQn6SrUPPPyknD3l13ETsp
Y+6QYQ7ns2nLc8y6G/ATBIKXoZJaUntL3UtfoSALyQy7PZfw1TOcCDrXTxXdoijvo2s5WWZsur8I
ZdF4g1N0eiyiPuwA4VJcan0IBXmmFYNb2npGQ5YfFTgew/NKrocPNBkTzOHgqr2Rmk1lYhWFvdMa
vj/5CABprv4MIHs0OenwYATUe5B0Od2PBFawApNfr5835rV2Pl5VMayx/eu531loWEFU4IJxhgfv
L0t3Znp0QOsYxj1t1KteCgBWAScuqcelvXEWm6EITBJz66VJhxVNqMD9anw7HetlT+s+C4oYUzBY
v2X1mI1lVUKdvS1wf8Mzz4v2Zz2i4jYcQqEQVDNAPnJvHv2AMSjIY5EWfH0vpPxi5bmof/qPPITT
gPiTBheIQlFi9p6XG9BxKWOPE7aHRw1IeuKIMhif80K2KxDDmo/SrLQMdNucVoZVCoFJYKlY7Cqb
7tIuNTiLKpMrfu3u0DLgn6vFY6fKxtkhbB07hol5HSwTjPOtwtM4oKdp97/VdealMIwXmFq0ZwXz
z23ZqfyP7tqhvXQO1y8g1++LSw4AV+gBoXDlKRJShWKEgfdMxzRzKrxccxdEkvyJWj763pG0HprL
8+EXlALnAAE11NB1mzjMnDkqzHuk9/1hciFw0UyT1KcGiqjDOjdj3w9CDlmrLsEd4U/U/sjjj6i/
vxlqqTOz3VaQpfRjahwX7dNOomSF7YtNqvxSFsXC2aFF6nrLYtYldr12TrhfLfqZ88UZLkw6F2Y4
ou0S6YGI8hpedMheJ5xqsI2s689sSiv0eem5HNAvnfmi86dL7/nmWyoaYJdBQlGzaGg0F3D6eXNj
947Vy5mhj1S8sGIDA3rlZqniQRJY7hdSwbL2/7JKq7Y5bnDMiEksV1TwL55tCNq8W0OzE89/Et1s
Ik+pp3BzGcFwiIhWvUxxxXfmxxzW+jDvHakOl9aRfegCV5ohfjeQZ4/fk7kqTSed2ReLRUTJa5eh
kKC1wCaNgluBuaauCAtxX+JTQ8yWpMuuU/fYCg3BF1wPfHr/LT6JT72//gvG5dh7pF9y6uw2wYxK
U3OUwHiN8Cr8QfvSnJw/VnJVduDsLDNKqRL+yTZAFanU7DmwjoNlj8vKL1x5THocDQBDuX9UmIgQ
t4wY3cQW6u7I7Graf9fcMHpBxPdh+OWA+LAihTaDyheQx7VdzOCrYv95aR+6tg5MgRoG3TTGPT+B
+X2ZcU9hkYz2OUpsQICVV5pwqqB9FohYqIfwTDZggvPEF+LZQ0THMVz8tQN7swiNR87RQNG/fQA7
1O3nMzoB5RUVHdiQnj6X4QXAD2P4kp+EWMVp4ceEUPSxKJfMAgnmu2qKq2SZrwo6c7EiAHutsnkO
3CQhWccu+9fhIZ+YHlBB6CG5ImNLViL3sNzepJ4gsi4JYMd76aVwWb5TWDmuAMbaY4AbDkcfhMMw
L0oSdlIs0edapgZMHZUfs/Vi2ImNV2PGFhyxC2MpdZtt9TmoN0bRuhxatp/VV12vLrGcoaj+UO+v
8a3XqTJCRzl9dc1z8xpSB8cIyotVHyG1OAFKI7wvsuyalglGi3jnerDy04mJ/h77m25mYZc3NIWH
EKFlGlVmGaAxKNL9+qVOe3Vxge0zQG9IX2sHK8WF5gqGIPYsCT2wNzEkbtUaMiRtXS45GcnyOIq6
FftUkRP+vn4O5SHtGfphUrJPNoKQmInu+hXI2k2zN+YZSoF6xqHykkKre0+MWvvElbh3NaHZ9ozH
xvhrTHaa9J7njjl8Y7BUmTSE6KkgoD+k5qCRBGzMYcRe3Z4izX1GSLnL96WhCTf68gtSfE7143o+
pVbA/fkYSbdUVfc2K446r2A134WAqOfb6gPY4JxAwBXctv4kPNWrX5+cQARIA4GE9gyrNfEbHkkX
PeG1zlBZm9CPcx4D6RW/nwzFf93uszId/JgChA6sDnd5/0N0osObujsdVAFJsEfCexSRPD+JRm+B
PvtwCfTehfegcHtujSUAl2U3eko4sm4Qv9RHPMzll3sBCom91uCJCTpU1l0oKJDIuhEJHtmI5rvq
wrX026foiVgxoX0QVARGzyGXLVuh+B+QT8pQGJi6oBbQiByeE1IedfwUEW+dSI4jGdIkT7v24lLI
UZgbyTsSf4LZzXtea5ENz0Cb4K5kDD6l3sZJqk6EgQTTbHtSjZE2XzpUDCIet5a/1Nw1Y5ZWUhdO
KbFOheKnM1qjgsI9yXowO1XjqaFioa1lXEzKhD2BagGCSXE3ccqFKC8UZs4znKP9oWpRlF7OLYXC
0YPtnmLBY9DF3/8mYXDvawUt7l4bApFBLzFEoZm5dXr5Swd85ZdNWpO964cRdH+3D5cS8k4iXKUx
XuRli22UCv86Pz9KaDYbMFDaGBzJshEcPG3tcNgHin6o+RUovvPMl8TvSRCk7rX7RSgyDdO81orC
ey4+3db25FARW/2l7AWkfGepntyO7Eyv+6pdQxKOBaeYQNQNArunIMPyuXMVXTpFBTtGWfV3kfBH
T516e78vFVhYB4iF9fkAE8QLJlcbIaOMBa5KXD0hwALUVLP5iPyYrwcfUtVZbuV5+4p7I3pTji2f
SSGC/LeWJuGjiQ7MC9l2oLx+Kje7lyftD9KbhkRWijKic/iSQckG0JxAUUUCd+OTW2rbXR6N7VIN
z3NUyQ0F5C9eXF7KLauM+CT3HoXpweMGI8wh58Ky/FaELyb1h2zjzWPIFykdZ3MogE4qC8qv0Eek
l7nKb/AORT/ndU7gXOaGW216AeassmV8nPXScwAl9vMIJgQG3JCl0L/AXUZY3cWLfhGgVDChdw0Y
PhsYzC+QTr+1+PmToXqeDVyrzquJYp3lR437PgZ+ppKEAt7tlvk/Z8z2oohZvUyIL75R7EVFwJq+
n6hAnhbRPZ9ff1poBAr3paSNz1oijBSyuM2Ps+snG6UGBSliMebz/jt2q7vReIyx24uEe79DGAoR
A74KqC7xUGfTsGFR+vE9ik3hM6S64HkyftKw8fvujZfxz6kE6/b+25RtrzNw+/5KsimdnjH3FSBe
SNRLgGrgUPw6fvcOBstCyxDUS4KKgB4gpEssrHtJCYLsVaFp9wm/pfUTdrOyb2lrax5pqS7pm/oK
xQ8RK32AGGKyWBKjd0Gk8qBEU356puUh0fGYFL6oc0wunuKWQ1/S89GuktOnUrhC6mTk4Ar1hEyW
6G1TWphFwTluuoGSeQNVAOljxXfRJ03ZrZ3Ym1ww61CUcwhBHewePf24O1lckfAvz9IyrFkYpCNb
hgVfMARWs6LF6qbxv6Kjs8PA/Ew2QYCE8kF1AdjJkT5nLP91a5ErM1kuM7KD/5W+l7nWHSRgNhJ+
fUQN392u6o6dpPStbvRxkJ678r7twprgaFcXM5b1ezrC1asfVjkIaPMpqryjJyi9GLGz7a67UynF
MYtbZXAvIBeRtxuZFpwfJ4lWHzY0Fz1vYv4GrPv4l8KX1tRIt8VS9bnfwiWqWMiRtHcG7Ogh0Kvg
xWNKcVhQGdwq0SuIIx51OVjRDJfH1YjAoV9DCnWKADP+EyutW76fdQeBMgB2zVJUzUTXFpb2UvWU
e1Ne5e1//5Wl3+8utMth+vnQM1u6ZzQG56R9Ac1ZXIRLq1id4/oTfH+F2bCkbBPc42MQXycQa3fh
8IzexS9bZbVH8B+/faky8Icef66+25sPoR1iOSugTZrD93lVCk1WozINHaoTnJdXMFqm7TuMiBPn
fq/7Tpx/96QsarjelIDdgUW94u+cmcZ9j754mKVJgQst2vP95ELr+h2Tqb/GBMPhfs6XOqf4LTKS
FxEMg0usTAYgLHJoMPW+nSc0iEuFsYE/Bkfwlf6xIqUVM7TTOCteGIHz9rGg7eHwNyu+tkKmgfAH
rFjRxFRTEQ3JlFdop1uolThAQbLUT6d2Jqhq9vJeeu3qWMzllQRLSUmpgwPcl45gRb8UL9mKXERd
9sY47qk8kuFIoVvEN/SrlfBlGwkipn+xRTAV48FshMxLknKS7igNt7XwXsgjE+SAjN7k5NYT7S6R
wHTaXl12sWJIKVgaofgbQerFT4PDniJs8/EpE05fidoPz0A7FdSFe5jOZngOcJiMb6SHQIhLx9SW
8fK4DxsclE4MkGaHYYZPuZcDlKmvgz84YqWIsUlgPGQ9ABZNKJQQlq4svJGwaXI78i1/EaRt+sKU
54UKKzt5xT/MrgXgPzwXePlH0pG2BQrIpX1PqVOXUB19SJVAkUph3e9VH6YQtFb3A+bxPIDEumcA
Xn+qtaJLiOsPpkLULa07IfOmQ7rgVtE4Q1QLF+iPar1EvIcRcrRZ3D1hIfRUAshD35J8LyKY6yZ2
pj/MnmEaPyKwsX2eaC5Gdvcg20Zx/Ws9UKXKyikv075JknrPXgHse5XNtRAo3WV+f95ZD9ExMDjN
xi8aT8BJhMuYppylFsSPcyfqMOtEhWbjOU3XV/LUvy0Phl2ThKWyKNuYe0D3rlBwfvnAIiHxC9J0
Iqb7yNBhghP3PFCMaGDgEuMNGXQE8NeIo7dqSUPh4YsIDY2HBJc5OrL+ADYTRBhbbNTNuavXFfCm
Nq9dJB+zgEr5bB4viKGHHhZIUDH9jFZG/lBZGmPo6O+0IBX4WNkAK/bPB3pugu3HwC5ziJGbPLWF
RHBMdJyjAJwgBogxubF/dlyDX7WOyx9tknWnbUfxXDf1SV34ksS/pJQL1+XllUCkqHs4WAG9AVXf
qQlMt/m2d8J9aiKMz4fk0Bf8LQr+xLYiUjxUKMDPAqnbY3pkcHqXlZcB/38ncAjwEw7LuS7hggyv
Qc7EiexOALdqvulkyoxJ9B+sDDI7YLVsjk4RhEtmuU1ucbCFrAvW4poV08RZfSwn3P691sU90iDl
sTpPxEToBrfXtqhYflLUIyvzhyx5G4KTOMVSLeFE6L1wYhFD8vnFIn9bYmKeatrtsccfvACmbr+X
Tcg+dS306rFFLiMkGgMdJLNeNuQ6ji32bt5zkqq4Yd9fEuXVZv1uZJRZIGVKFxRO5KwEiKlzUYww
+SjeEjy48rI/pGV/YXvohGPkv9G1tEmDDTbrE2FUg87JrqpXJdVWfDBfoavhif3Ehic1E0fvyM3T
mXFknqzSV6rPVLuUBFTpLsBw0hc54lIwyzrv3flEcaQpXtLZ0QHCJVge/sUDAEjQiZifPuogCaRl
0J0Kq7E32e1DPdtFKDzdQMVWwOWIt8KAJ8eNH1eaemwoirFcEgq+xrNJvDCZ7ZszkCtX6U3DV4e2
o1rVM/FAy7Ej86jknKnPh83pMPGgd9sn+V9B/l3Vij2bsWY0Tdt/PY1mlvCYeVfMVD24Ev/X1gFo
dFihIjymaG27XuG4wR3nBI6FK1PYm1hQP1vg4JvOJY8gIqHzvMdAg5FUo+yOyBBpvkhvmh6+hS/N
e9jLUnyyKGn97nOhDt/0CI+HiKH2XrI28wLL09ZBEq0PgYDeP8FESA6NF8Oq4Bg8n+FILR6DBOEC
rWJf+sXrfMvE/7P7QeLLOXoIwUivw3bsc0jEvFDTytW42/T4yM9hPd5rBDyRXl5c9ruEgXEWa8Mb
SzTlL6omyfXY7ajttpo0RBwRYvnKGh3caG4tNt0Ep1ibjuHSRMjELfwGPVo22cSh6tYmddTfqJ/T
KJdJ8B2qEzzGxFAtldNaUp26bDJtvthBIHZct/DMjQTFWG6JNuea/Q+B9JMyVe+ufiuouUimQjvV
i3zzyjd83U8BDP1p05Q8rEovOPyT8Cq1wXuXcR3XSyS2tHlev0BlUNvf9pIKLX+ikVRjx5uJALRx
/D5QGB3ADXtsLsxstg/Ua+KWKDQvwnrVa6V4dzUv37o8ljgpoXzB6AY6ZgS+nyp6Q9UDVyu8+dJr
6BVowYW0pLNlACssZYsC5S42Y3JRoehduQUuFmyuDT5mV7se/KTV69Nvj97ng37uDX9F0CG3yD37
n8yWws8rY0UCM8mgvWzLUlEZ82i54DDzr7xzOFvjicatXuGRbZWL1GvDIvYnp6jlmXR+t0+z5yTq
55Y40izzDrRgCbcEGlRqsZuurjDoz5VvUxJHeuK3fq+CImnoWGQ8UvR7ssU5tnnAZHHGw3UjP2XW
JoJzUx19KTvgnmAxpodlZiVIfOZJFJqcuATkkek+XPYHVMpgJrOCLUt74Ccn92keXvFN+tCtDSbq
+Pnl2s2DEBj7z/Oaw6HzThPT1pj6p85eF1mDIYlGYgPqAhnW0OKFTofVJGqMeg7CPkNNNWhLo0op
pHglGirBV4MgR8ahVF90loaCKYcmUlhbIy3ZLSOw6Lc2paPWGlFoQ4tgIisCMQfIpa/H/rmixwCx
czSFDmusjVVNTYE+UksGLMMJaT9z4nDmjlHmOxhxUHw0JSTXw0nkmFHVEWgapVYNIwg2jnC1HgzL
iOJMXTLg8LEHfuO9P9ObD1NQ68avclfVWyENPpDKVjuVoGs1u1H9clnEE9RP2jdVOTjh2Gkbre0J
cXDBpDuoZI6wS/heHEYb2nbxyAIQO4tJFP9TIunIuxphxIBBBu/rsUxkzDkrFmzDd/HjYagTM5T6
+cj+792j7dkhTSwtAMDYSW1QnxzGRkyLBZG2a7O61rIWUZV9e23TQYqqrLe/TI6E0lMEs39cEmxl
64A3LbHVRP8M0KjMj93jtqgRS5H0MPkrzXEgq76syapkJDdSbr6clAiiBWclkJxY9ZSV5cdWzOF5
QTZ+Pm4MMDEtpjH6P+v+A6t/J5TL+QgvEzCm1n5Rf4YWTEffcOis+nec7JQyrm4sQ6Al55BsWyuz
af/2f675hlW2f5LGKnah82YXSOWuT3T0Bk37KdYt5CRAkW1cLuNo+xO5p8RUWgCjp8avVpO1S2wG
n41wIDLFui972W8BIsne8Frgr6tjQrs/C+gErOFIXSizkJROWdCLFtNJyYQhybma8DeMgXBqmr6R
Ass+vvotoCcFjGAY42ecJ1bAEYxUjpb9ISJY31jCfzLr6lmR9qNZTVHqCXKLmajtl04NWr3mAuoC
kTJfPjFDueTcQqPFUiQHbjV9jfRdNhuTD7Wk7ixp/6TLkL0eszCFNSIYLfUpkRZun3+IRpuZbZFK
BCQW2THxcRDrB4F/ArSzNtMAmxgscTbagsddTf5o1c8pZI3OEIjzuTI9sHqT2XjjHA1OwxB7y56k
1kkM+1MhMhR+g5LX9hOYDE06gUvXPGjLJznmOJFOlwhYiRvV6yOOMYFQI3RVpjVnbUQx+bqaN07P
+ZdC6nW7VqNIp8C47FBl1R4QpYgGrQwb7AJYNxxt/r2QG6ps1gRs/6z8b+xcvxJkPOPnD5DnU0Qy
GLb96XXzbqFiHjVu5VeCJKrxZsrKMHHhjPPU4vq34ywYeRVDefMn1K1us9paR5GqYZiD0+Wp/3zn
lf2lqaY9BdX2PNzk+iCYdYehMHfT+BN4JZJ3J5WyWK3e9haBQ8fjio9cDjRXWO/BBtzSDrqFAUT1
Yone0tXmHS27+TrV1lKP0L56cJTp5JdjJdC9ZXd1xguOjiolC7JWxTEm6r/PAgl7yZijUc2gchjK
WwMEqdBMMAhaZsnb1bbO0vz0Xxfqmo2xADH7JoTIerRaTfGvxRDeshVqLpFqA3cEAgTT1neg0ZUf
KF+Js1bfV2o0QP9/RCnsS7wLYVccu5uQVm0GN8aVvQ2lwYxpjQjJ0uppHdYGhPvra8KohsNFvsKt
zhpJs4IkvDDcngulwSm52xHZGcmVaSqyVO7Demsi2536k1NDTZ9bW9R1SnGpOCmqsUWH+lrDeeMb
mMlC63X4q5zt41JLr3sNuGcPuqc3dC7zHnkR2AZQ1xNs2ti2NAsZD7V3qd8lNsFISNC7vtSXGaGP
O9TrkG0gw2y1fA3f+Gr8SPlzCFNrttpKjgYMDtI6DZkvPsCDUXUZR7peh8+BzjnJ4VZzvk19ls/F
ucCerOje6HJPgt6owxmyL+yB9vyA/sMbWbQGfa1gcNYUX6PBBWDLupj1a2nKVSSqGVIYdMgnBIIZ
un349E8k8Fl64RcvJq6l+kUerAPF6wgYhvNasAQ8dolpAwwYJ1bhVvaVF2Zm0RGOjQT2dPhiOGz8
7x+iaaNx3P5vZjRSthscTR/Hdqda3u8v452BY/Y7ehyA/1cWyKH/wWqF/RvVatnG+pOcKS9N9RT1
OVRFCh/0fy+0ctKGa9WzfIYIN3hZJvpJjM2ugOgPXGCyqdoBXcLVRjFIsnJetbCEaK61vyYoWFKv
V/KVmwJ7rrhr4NwSr0b+GcoZr+G4WcUemRdkO/ALLiqBBq72U3Ea2R6AP2MahIZ4Ls+1lCYwR1rM
32RYg74VP2rTeWRZFIWjfyLcX+Zubj+OINXA5+CsqN7hL2kFoZ3m2EwpaOmcCTo8AqIVC733RpYG
oeMz6/qUHSWQbTEP5rW6drReOjsSehYYctyzlwY0LAm9xSPRepdTgOxIphxqDPfmusxEXMLQdfqZ
jZHSlWw3u04j9azKv0yAXnW1xGzhTUu2R5VsWHIzeZ1THzE1jVbGEzkR2QIrra+oJ9jiVSA/s/TJ
uhr3oRkhaCPWr9Pf9D3JRWX9s4IFek1MbvInXmDURC7sVty2lxpzvyyFkU80T4p+wEuir+E/O7f4
R0j/ksd0Gw8kYzDmv3sLwl7ssx9Wsdp8OE1Q84CDnXW6df6tU24pHTSJvEWSE3GJPnkwbotOM5W7
WLAncYnztP5NyRXyRREFX40DZ9M1FIMUoCN53QXNRhNfguR7SCf0e+6Q1fwC3o3uFvw38fGXKzZW
TDIivFx227gB/geqX3EIRTTtIVO9bs55CLsR+Cd8UW3Ekd9wu84K7c//Lba/JtMj7aQiCPNKgLDd
MP6+sxhr65yQ6O33ZCX7rM7J40/BfNYKeLZjpxw/Tgf2np/F6I7X9dp0I77yevskA5fBS64qUsli
G5/mcRrqndcBZQ/NBxG2F7m2iwtJySz229S9FvNmqdzQwE080fDO1wQFawb6utrJG2b94dODaYiv
+cC7CKBNmF2ka73iYipi1o/ZArPu1NkabAxlQq0zIfxHMWk9dacKs6skAlkZjRVfC4dYnb04GmHB
kejm3V3VNd2N9ZH9xkCddI9lJxFkFxdkW6x6qMml4jYR0RFDOkWUMTT7mdYT838gUovH86t5t0fT
d7tk35PM7+a9nkCm8pfIQ81cJ8ajjLpNalKNTADFt4FqxP/jqFwnSYXU0Smkkz/pJjp9mTHnQmOT
YsySWxHfub1OKwMTTvZ6qRI+QDpTAIOz06BT89ggB9goetL63lEVWDLEbD15ask/MbRn7HKrbe5o
sHaepA9ZgR+ZS+sB6nelw+93RidYYFUvWAEsLiitmq8CgvnDduyfxBe8r9CuWPDI5HBf/HeJjeXJ
QgDtW+SQ63uYZ1i9n0eJKldLyjIKDM8xJkxkLdA2kgFnaqCsDZBMNTjI4fdHElBzLmNdQ+QL2jJg
jkyXzeX9BZxS4Uc1d1uzXQfQyE2MnZsazgq2WGvwWyIklm1626GhCgdEmues1MHoP+qV2AWFGa5Y
ZYCrimNxIC0kfmslAxNHSbwceibV9qBGyoRkKIwyb2huHlP2j46gWXLXFEjmZgbd4PiPe4yEoQrZ
9b/GEPmBAmP7cTPJig4cKN6cwDi+mSCFdcnkSKAZ/feRhyBB3iene634sCW1WayCTL4Oc/ObwyEV
jfodov18IATzYT10B8UN2FyJ2i6AU7Lfw0EsqXRx/WDHpCGMjqFiasKcNNMDHKE2eq7nWkGWchVW
DSh0swt53t3Mbxo4qPEzo9sloaAwX1OgeKVOUMW6nEjSGYNYxJkpRQbM5OdYMqB784v0GAI2jdbu
WtmV8xHa3yVLKr01MyaoyGapc7aUi3B5VngrCPkKyLJy+XqSjdB3TrfWPejWol7YKk7Y04ciEoYc
R0BE0GEvyP+fFZxzs9e3eqUeEYvzROhYvVi6gVAKJ8qrSZP+DFjCBhkyaHlmudYMbPqrjerir6aB
qc+Lg8hBL37/6Npsq9nlUHLncMoL6bLCxV+/zwXVW6822cXXay75e72CT5/ayENqxAdeMs5NFTIe
XSeToHruCvJFpI9tCw2vwXSWxsWyyRadgIUkammMMeEOjdB6QwRVCtkwkXrb59fclWWL9DhDYAM4
s6gG37KTNGWqq1FxhJDy1jNcJ9l2IWhA8m8ABqkpBAyZNw49nG1dWlfOsnV8wFGn/2MltUIY7f3J
mmdTAYytqqUN/13ODElUHB8/HpkYSoWsKbJHIfdJb4rhj/lPz4RgeYe4nPQ2quMY+4vaOKHrk61h
5I38EwIu1MzB96QT9dgTksSLs3mgBIq3Go0qT6YJVPJw63v523kOq2j6r267O+0zw40GrKpsFRkW
PXFt0gnwD3oKFceF+bjeaWK1LqGcDaPGE+LIRSfkn/4Umx1WsQqPnKYb7tGeWWxrgQH8hgfahC02
slw3g356uRC6g2Uvs1YCXjcrET1fviSbvEulHyutyBMSHXhFYSfh9zs6Uezdb+AjruKE+UKSaEIw
qdX76Nov3zBvCYtDNkx9+N1CcU3ZFUKBs6eWLZBlvBLKrAFrDPHMegLdo/lA0yIDivmyjhh5gQ8l
X6yrZ/zb1oZ3AVFU5bxo+0frrKmRI6euvPtSWf9YxcY8vGK3j6dKOQUwtJw9ihwF4noIg1hleLgk
W9Io2OCr2BFuMYqcACNWlOfujvm359pzeMF+wPP5Gse1tsV1OIa+BTjf5xlzVK1qQoVwh8M/o+Ag
8nJnJ1cD8qppc4h+2xoxVxKgh/XziPm0eICKm1lO6B3wIgXto40VBn7DLV89DjhZQ+4TEgFmg47X
xvJP/NgWkjddxnE6WSXC4E17emcZqMPTLy6S9do1iGJwKTax5ML7Lm5pJ0RBCxnoXUJDayXnKj/o
kuUUt8t9XzKHJGwPmkP1vrPBBRVJkCdFBtPjgXD8Wa3BZSVBC5NLfhmaAAaN6X9kytngkwyWPktK
tM0/JFcqg2On7ZG+qgd/PTM8yi50fxi/G9cBHCZCfApNp1s8BPndKTSvACkiZ+rhlyj8T7n3NUfW
sx5K+Ob03+/isINUkCk77SqQG0p3Dju48qTmMh1AeEN13ofdk/UyeD6deLVs1GICQsqMinEYC4sK
W/QcePuj33acfWn3ibi+olQ8z4RKuV7asUHjlpfp3DMLd3FMltpQIk1xqhR3lRgBffw9LgQnHOmF
eX8EU8ppNLvPTwtCBFfGRs/8+6fV5hNzzEYAnhHfib7dt9uuHdiv572QkrfChyq2cNRkTWJPRtAP
3AnlwwZdln3Y1EcXjVqgA+X0Hvcr6gj0hWP4bsXRfCGjyaV95BHW3IfL+Jc004V05DwH13Am8+jl
CI4FQCc0NYLQcsIBi4vLHdDxmk4i427kPYer2c24WT64rTXR52Cil+myHDv+DJLztWTxl4jje5tq
l3jY0LWu2LuSJNdvpIrMTSU/H9oTDyd85XyUyr2qhmK1T09qTWjHle3dlM8yBlDToRyeN/Wknf3S
aVIs2o7DqVroMkZ/b6vEesoYpEkBFXjYOAYOI3+TSGLPoGGqRwbsw7tGP5f31HE5O8sd1bibOcsj
OhbyohCV31hf7ukXJ6upbdzVcYDyrsEJn37xOTO7dk4M/XI+M/1COviszrM2AR6oRX6kbTmkO9Hd
7U4LD9sC9gIsdDw6lx4x8FfPjPrw8KZahe120+xbmKP6RsBgLVFkY7FDk8LKOVSqh7BBtqrooQ/g
3jwHNbvlN53hkskxfL2Bi0XtRJw0qkDVSw0qewepR+x4zQHUAvypHxnnWUSyjRNdJEtDo9q4KzRe
xEWXObZvk4Dm9MavaA3nu65Qiwe8h6e7WcKk9gQgq9JAAcECfQOYwL7WQqUFXlqgixnQS9GwfBcT
3bYQj8+dVeC8MZO5TEz5oIiD/KbfQ4VC4sF0en8UyheAW8OxTGuZrHk06XtuegN8VMko/ZX7m2lf
Rfa3CqPpqCGp4wEzrqRVoHAe8XE7z/AthcQjNOWBp7LySo7Qabv/BHNYfWeP9RHCS9wSlJOJxYrz
xGqm62zdfdk1bFMubBd+Q87LyqVw3MYw5GHl3RQBFzYovggKZLye8Fs8G7+3QV+MBC+0TG4yXA5g
HWAFj24WgsdBP37IQ6X9oR8CIjZIsoVNhSXnCy+UTK4cpC4AwnWaNUQO3LG+2/5shjM5b6ucI9Lx
q5cNN20g0KuO01IPDh434ingh9J8hwqipXQW0QSgVJHva0YdrME5mMtyoQFPJHe/h8/xligjqihs
XGHSks6Wl/alGiIq4gVvLUF0PjYh662LcArZ3Twzrl4qdyucFPQlAo4fFOGqICDH79ErtSRraNhM
gvFR8KiMFCwI2QNX2r8wFQMQrbYfphqtjUJTTyk11jBCXQekWReJogy66ehDIOW1QIyrEh958rgd
9LBciOlqC7JKS9Vzg7irnNL52YQb0RgD+expYBMtnRCq+h0lpbBXeyGNOFFbVUXeWdYAmJ5kK728
9FexkP5RYSOoMRO1TCy0gX+RcHs4QIGrfkdV4iS3jcYKjAdm8cjucbVZire/2cgyaneDiSjhqGBh
m+wo0h7ZzaOWYuCeHXQZ57yB09Ob03wR8nO7vymqq6kP+HhwUiyk66QAao/3HBQeKVfKrBG+HZ8A
FsjiroYLvY4KgOYPKlD3o5dwVQQMZzDByr/uyoYCyuznRRqv/kRgQyKIh358EGDbmeKtrl92lEUM
lsqjoAefFuJKpr7ipwRzcK7zvYcfDuNjXmcuessWLH7NTeQ8HWdYhuovM6cJzHmDn7dHJtMTdR0H
SdBbhlxjw0sagYvDY1uuoYih8F0y8CiBZolrbcirNcJ8bvVsJ1rx1sQebwxKfqseV/MNA0SD62Ne
CGLUIDaDTIKnmR9QUlncKy8MZQ/cr7grMglNYPAEil0K0gU1kdqqT9HGDLNMMo88iJx0pBYg0rek
R8FqYeKUUiqniBVlvsJJ1xhTss6otLJOtYE8TfcpF0yLhnCc2hlDQd9KFwiIjk0GfU2Rq7Q8AOKP
XRjRmbBHCwOJvQ7CkY+fsBRzr1DFjpnJ05qN6d7I4K+NveFJ0UlM4ENnIFsG8u63j1RvFbheIkt1
cF38gihJ1ZmrWjT19MbE1vT0PVlWmbjenP9zoPyolpCTTOmZHAUiUa3n75PMc/Fb6RRHScBsA19r
PkJegJUK9X3pwsBtt/V08OueByDVWPsTDU+NMQMbqExpbZNFYYbYgCvcZAtxN0K07vegE5R93mMr
MREmvMEHQlwDxTw3mMAtYDeDOasis/3r581y/3e994tbUnvQ//ZWA2AYDZ8VvWH9XQzZxMiL9fjB
1Knp3P0HA9S3qQVr1tVTspjHERhbnndxA3fhemCi1e6MUo/K3QGhIwsUiA/CHgIPER7SrjQOjDdb
93FvELDmX0ie7i9xM5TItPkyPIdnm8UugLFUxawSuRb3SNu/motj6kUQb3U/lamn+/nqG1qpaYeZ
+3pWiCUtCGqZfMbcEsoWbgVeWzsseeYa/qS4C3jt1V4CQIe5vGWFuGG4EBFdnu8pA7YxL/y5cxd6
0kv+uLjmOGb/6zMD8BQXFKoWQgK3D025QvPGZ3ebWGEUuJ042c831WTo23mCl63bVR2RRvVKAJMo
dIY0H56Bdeq0Fra1cFH4k6lwKAFywBTVOBv1JePqISmzmOz895AKSq4Dr0QmPwnpZl5pGEIkV2RW
nvB+Bl83VavDWeejoHPZl20hMrdJIwqLEBcqfLAgM1/c0O0bvHRYqxIlDEX+9T3KQ/1owKQzRMG6
gayQVagyV4pR31Gb2h15E8HlZRQsKpTu5eZfGOMhE5fVCdG8Zt1zgZ1yuA4OQLd2apdGWbNVPvJ5
oW0ltPQn7RpdJrRpGZPht8rgZY1KjiRcgHl1It0fD/US+bblDtDHTUd/uZLDSiJN+inWMcAGQ9O6
VE1RhqLB3Pj3GaI05cvJSrRkMS4yX2WkmwOf6Xw1+YVZ9UrBoMi6o2TYh7Dpi7cnE6/CV1rLmETp
+dUNvqrIv8fMHRu1Zv4qloXw+JH1nHZA9bREpy2XtqbAHOcwJeFQYj+D6Ive8x49Dm1jC40tVU/U
jEdicURoatW/U8WoB/AsQSxvoXaB7oqsxemPMFFpJngjHQ8fomPCehUWGGyXF4wdFBTUfgh4wPb0
5kn7GaYzi1Q72V0e4qJJzh+H/XgCbjJtZDGw/3xcPQfhmOofnnNzofqxFLxU510gqB82QOUXVn65
ibP7gEBm9AGq8Ap0OyqLsMNSkkCh9kDkCvlcVA4iyloH3MW2eIreFGzSgBx7kycjMRbrR+7Ud6Lh
y501NyGIistY+AWAPcqsIqhVlllLyjbD+hayJVSSsqooQ6KRWKwX8ooIh6IEww1HZU+HDvewoaSl
tgxHGSppOHMa9MYm0HIOZcDLtQFcEICcf3bRmBpqZ3j09ny8moSptSVYqdNZ+r6U4UW7uHB0iI/w
w2qe92cNJGx89X41mKs3vFA6D11SPiDI1OAblf+ZyTTr1q9Qo5E/gDVbzouWnMa5a1aVBwm1ka7W
fI68oOXWCi6pj7CV2YR6zGNga43+9hdd0sOechFKCRwpRGhKnEbeYwkDCRZ21tJFCxHjcpjicvtu
/QhaLD3y5nthNpEEfLjPmiVMP3s7Z6zgHpN4vPRBa7NDEV/v/aLwx28NA4qumX966hCv8jaFlJDA
czFzR3hq+XGGjp768Cc4mzZT0SygbPEDn9rBMc36xRnIjlVSLDiHrx9q8bXPBscRljJL35Sj4G1t
rlDyelyCNLhCMGqa56geQuqJo5AlYh4vefI86CdgyeaQPxP6mEZT57HXx7PLHPte/qwWebfLE2Ky
LRDp+WAJ67bl6KeMhXLziFPDQbL4VjO1/ojzCyY2T+g1VmnN5U/OH5NPXiJg/HBsmJ/utBu/vpqU
jIdrkLHWY1mifcftiZcfUDvlKu4ggR4wvIDeasYmbvxKPpUL6ffFVu8PMRIvVxN+iR3+za5GxWQE
cl7UeWYnMAu72nsEy2vJSPBJODmsARV79iHpHKsAf7bfDN/agIS6gtOAUZYvns4eJ02oRzfZO6D9
d4NckHK3QKLw3QHazs6FuEOTbIEuUKNZ38IqItSRZ9wyXpLJZmK11dqfWd/UNe3UEKBY8zQ2JDX9
fcY8qgR9yX5DtCZEo4Fp79MT/v5KQWjgUgAEl+nHrHU9v0j9pk46jgKQZMs6q3wuNpM6QtHijeDw
Ibcwm9+astUyrE7deNxnlNCpbDpnbKxRRS0tIVQJqYyY/gze3gHRLR7niEeWXTLYGjdGxUPxVQNO
niuk8SlV2mXGBOJfTAfGdtpxJFM03UHdk6Z41A2Ha4088MUdx1qRu5IFnG8jVv6EynluE8Eh6UnE
obltPBwxEghCjbp1bpT915JxvdtHawpoDIYFNgpHWKkiulG+TEOq2OPzIgy0IPJIuiiHhHKq8baD
7zSoyIJRxAFv7d+hFcvmgEoxB70FMaT3rnWWqgC1iGZFqyFsVW/qAGMnK8NQjwHB39g/XDVVdiyM
RjvtSrH2w9+nYr5gH8gUC3+6Gs1xS5+MibkbYvtFYeCrPfGW3fxpiCyw4uitdpz8oDQc9dkjF/IS
blqwvekkfA9YO0aH92RYDEEHwQiy3BKOdyqtuOAMvU8wl7nlVX2gllgBILhzkZzlCu1BW65bsCEq
iqz/AAf1CUQE9EtTA8xZJxfM7PTl7bCD91qlJILu+ADFfR4Uyo/0onVAqmoVFGheDKNcUeDe39R/
haGhE9ZDOG5Qz1fYZyLWb3lMypqJkCAYEu6X7ZSpe/QQdzh8wBhylDeVGkXBa8sZJoe7k6zyYSYK
gGTN6aOOLNlN6ezaCp47Te4vmJEyb6GwupghKuMexM6GV04rOxkpTE6zZrOnhoRWH+h6Q7LawjOJ
Gw2ifkgmwMX59Bsi3fdYd+GSspvxf0/traNaweDTysVJ1+0yhy9oLkEM6QIWKEhmGXZbGoBum1pK
B5pTSRtPAZ1HOtcwG1HZ5zikjy5Iq2dtMsvrV1dshrFj7Kd5ECNCvj4O7FbdLoQbcjRl9YfDLbYs
VfeN0k8rr2GgUsyCKWgSFrmPW6kHGditLXeQhbCwzn5bCB2+7NTKnXCIdk3sgjvOK1z8HmGOD4EV
Y4Ag3J+JVxT/lZuO906QNt0pqZNGwZc0dT82dnpeOsqwnQnhVwaV7LoflXMso2jIqV67osGfeSrH
FOFyc7YKr93+9gL/bsveIVT721RBCgdbG6PxFBn2lDm3s+fEwibBkk819dFkC4FxyQLrliqUo6DQ
mIZEJKMkZiOhwNEF0vuhiDNIdtZH6jSh9hP/ImP59KgI0AmSrVlLD6tL9lwspX7IA8FDfjKUylhF
AfOSZBGpu/cfc0HH+xGLNRmYcPu9riHUg70Aa7QVuUehrOh6MX8/NilLO/Shj6Qyr6+o1dQ1jB+k
mb77ZUj+BlRzY3mOFeW7mjv1Azjm+WPzEP0+1hZaUOKK6ljmz9fcmbaOshH7UOFYJd1yQFCAoXYv
ZDJzPKrY5S2R/4tLwwr8iSJKy1PrRH9hY098/TCPcTblSyV0dg2QdsltW73nZbJwN7s4SMLiPSg6
yYIBkL+v1MahbM49J/WB+Y4hFbXiRwsXxzgorcx9aMIIPwvDVBIMF/VF7/ihq28rF9EvasfHTelV
kGeMgXs4aRlcn7indP24/HNX8EfhGBwDBKaigORVDN9hCstem4sbCjBuATEhLwm1F+TYqwU08UX0
9RgMRE+ZnZNoH7FrVX7X8JQ2hXpKQcMb3hWd9MR6hFjTby1Nex/YvOuC4Svh64d7GTi0J6AL29rA
rHKyVqWuj3P11YqCDHp2nflTLFzZt0cjd4mdvx/EnIFezxsZtD5sD9zBOA2BTbpc+E/jU7ILdZD7
NOAk6sBgkm3wYiJn+uuKhcLBNHj59T4aqv9AIhPJB6at+odpswDQNUGWJ8GjxVKe1OY18b8aaRrb
7wMxdjpnnTpsJdd8/HUgNPnWIWd/RYKovBFz6YrlJGSBdt35HkgsINsnJ8VFptIcE1j6jPcsqTF8
qgM/wc6HFqDn7HxjwPIh3oWtePrVP7RIQ1+mMYKgMB0PwI8jKJk/xNHgQ35PiWWcSnR6eZ6Ls64q
bIy8W5UEssBBew8pAB78KxTOH+GvIgJzNgwvvMAr0AtinJleTDo5YyxTv3z3CMgvjdthiBxJ1FBV
rt+ryPK6cOZY1w95ZZ55Wjon+TCSAFR/CJwMy4wRpxXnk43XVrXjUIXXivHMkwBS1H3OpIShyZQv
bnlLz7TgnUEIjOkra49GVChrHbjkkLudeniuZDkGLsY2PyqpcRmpWoU6K/iloNKPAeOZneI6MxT6
FYvj1vsaEDzucIieRQM7G9HBJqZtIh975Q6cffe6PifYUbO2wsk9og6DTy6XrTIE0bbSRjsExlQS
3j/w+mWBf1II4oWwHRjFpHcq38bId01rF0IakZWquPhmFNVE4+FrhSp0NYNXf7mn12H6gsJYwVha
qMxOuoF/66wHqvh3/32+3YlTPR2iC/ZT15ObZgijEhwDyKYc/avSvk8p2TgbPlQaWyGEY6yrHO+J
w/HFilpEi3B1rS81TMqiGEDYjd6/NgFGA7kT1hxmx6QpvrfH98eEUU/YYXe7CElNnxgqEylTgAQa
4v7RxN16sL4WyHHIzYbfKUi9i/AJEpbscFXxpXhBJOKOIIFA2xrtWJxa/jqqv95VdxO0EnBUeNpJ
QJhiOLF4pIpE7A2xrQ2VuM5SUTUs2ZTXEkYEfUvZ8WplYfOJ1BIQLSOzuz4UvokemZqUCY6gVwbH
/7khtDz3CgpBAX3BYcIzlzsIaKMvKZDmZEFSu8WM3UtMC2xQL/+BRJo604cncFtxIWxQxBmEV8xI
fiE4zAZuwD9dVwz2otIigtiVWPJACd6zVrhxw4Wc2e71f2knQnj2jVY+CIMqvmIvNvmH0B8KqZKV
hnOBlsPBjkn4YxEOv0h315FS6wK+uWGrKhYlvTd9xCm+qoJoCsZXO1tNrumnN4h9kV5hgXXUd1cm
FBPLawye9Ih8L/WT4HOhNEx2u6qAPmI3yVoYsvrLUHT3IZSTx6I8uql1cW3HtMdVo38YLUQLh7n6
n/FxblY1QgfOEDN98Jpsoza2yvJr/cN00FMKbrSGnkCPUwXJTZ/xQNTy+RnUUmPCDe29a6Vfa3bB
21yT4HeLKvs+9P3VO8UaGTTn+wSiEJFunaw7gjs8Rtz5san5t9es6mIzNk2apnkjxLqzioKUl72E
BpQYZ9t0+b5AAqxRkTC6G0CRm9a+nEwxrYeyvYblnOOYn90WxKH+OqmGichrwvcCKXu3aozHIUSE
GQ4GcIL7HX5T96cH50VlbDvVQeB32FMBaQLZCeCnv1ZEWAGX8e6DeiDuGcB2DvHGP/giPzr6cDO/
K8eNHOyXKEaEwLuRyHwDUL2Y7LGPszzK3Hyby1wPZC+/zXlgLxqKpdJtSnNRSW/y0qoRZaDugl7b
SGos4hEt46/eEXf6qlUbu7V71CK/tod86EayI1o/KEztaV//CJaFcwB6wrLeMa9MPRYNE+UbQ9Qw
P6H6gZ3Cw5tAMRlZny2go9hfQsxstqZuV53N4VrVpkshPV26K6N+r6VvgLOptiDZMAbxtP4bw88X
OQsQR13QKPYX/wJfZglbVuEhfwPtm8tjWMxDsczRCuL2NEUqWfTZ8H6GKvOx70lvPP80JaM5ZIRY
nNIn7IzFOhaLELcwxovuoZmGmHSUaY40eBq/zHsuLZuK+lBuXTvgfjO2e04Y4zVWR4sTseIbSAPZ
4VfXQ1f49AAWbYzbSYtDroc3TBaTCA2ncWYwF7k3kspm1P+zM2Av+6ytDbn/7oalKfnlNBIzQAQ7
bPVA0saypyTPqC7HVzLZ7sQHgppqyf+t7/M69O1HeLr3YjmyllZLp/galb8rmRU0C419BsOQlYIZ
sx6aXXVW3zSkYcJET4o4421mfJ5jRMznsZAc1wdkdN6Kjya09/dsnxmMKrDK4u0eFVOJPUCqcMCD
PBfulv/+UrXnj7arygTB8zamqw0D6ZuKD6jqrDcWHqiHEfUWk0bHwPsp5kgzIhL8cvycZy6ezEu8
bD86WPpzsh71snTnlbBrFN3BKu3/Bj2rMM0Z+mmP2Zufs7lRuX/oewUjHZKfcGTWDdaSlTxwiTG0
vgBQFvXu7nrEY/5VSULr1ckmSlqxIBtcZTRLIsJU3qFfdYWb2dCW5U4ulM3eOEM1qTBVN8iZO+Zk
UgQE5ug/ARGn9VdPm5mYUypumUKBjaQgY+nas0RiKT4H1vw5KJkyePfrTuZftoSWgUWHWU90uz5p
kNMUFJlJQAhynB3prws/jpDhnziIsPSiKgtjaxL0vHFZXymoIxzJQNwDRtJ1EQkRJjLEwGbADfF1
CpceEFGnea1YXT0uXgwiirUEHOeOW8KWm6xi4ip1QU69M48EUgoqcfN12ufmzJs3QK3myTZ2kvT2
kXo6DCBXqDjqrwgzwZ0XJceGCLCpxdDnEf9c09D5tjOm6vekHD42REcp7z3y5ne80Fgy9xFSup1r
DwvzLODbQTc+CBaneoNeMuTZQBfbs2n+423owLXqRvai0J+s49YVWE1hkkEVihUb+FoOjn1eKSBX
4SNvGdoe6SH4ychJf1AWiKV6BXph0U51yGwIZNf9NMKL9wRiXDcjAYzbIOAof9JD7Q67EyzZT8s8
DuS2T9x09v/YeQudwcSwk79QGvLjMUDH+0HAXjaeXhdmJJEvjv8rm2Ar5glBw/lKPKEAMkD2HNXn
BtWwl08eBRGYLmkWLbjix6rh/ddyi7dE1y5UZyMtMAtjj37qWCr3TVa5LmfLwEmz/bv6XSyQJhSC
lbeECpLnce3Sjf1S+PyheyxjQ4Jpq3+W/5NYeCXeKFmpFIynrMtxA4ZT63N4W7yIllM0Dhh/s3yU
DmaEybRCAoHdFJXiUU8F3Q/M1detBs1BkfFgI8yVcobEIYrA53092oxpKK20sqPnoJ9EcRguvggb
7sF4imOlQk7CAPmisGuCZmLoJppjlOg4KSNKHHN0Hc4XB8P6rUCFLEcMktcR7VMWXaXKO52bd7Mm
7dbSDy6gbQgQ66TUFsHjLuPqX1t5yt5m6CFz+ADWaVuIFm6GjP0uvdvdanV45oY1uIiJnBZfoa4y
4nktnc58/3ZJLuhikaiuo99Uh9Rf4tDY6kiNS3lFW/ifxfEQQ8mDGs5tT3W6dLVh5xG1buexA9FH
B5NNiRymi0chZw/wJtqqNqAh3cs3Cw16rCzoswHAWqdRrfwT3t+F434ZjCztnEgDC3smrJQQ6Zz/
dVLmQxcTNRBPea6rupLQoTUifY78f1kwwDyqcrr+OqrM8c/GqoBSsn60TjRjWHtcdnY0qk5WwXXh
vdSsw7Bc43+ongob8xEauXYs8dd+6r/6tIekDTIpL4yw8YJTI7VLXS+xeRCSzpYxbAgF7JPUaZUQ
+LaY70k9bO0nnWDWvmVkGbSfwS4wcke3Niy+++5+QDNriTO2TD3EgPgID9Fpg3rpztTsAnJothoh
TsI/TEm1gd51O+/uXZowExdrilSzsw3H/lmQK6e/YQeM9T0KZ+nKIDMDWp+d8RXd5YzCgsaMN1lY
bBiOY6OwiB3AgTJlab3MSCQyccByoJLWhA6QbEUcLTy7LKqk9NBpFU+gnx2Bc7pvXxMg71nXEQDH
/NmV44cTAlo3/CK3sjzUY8HAj2WnPdHcqX09oWrIRyC13DX4nYqvci6hZor+tCalYFDtARFz/XgT
XTJHTvKLt4BE8tTy03FCCYj0ziev70pO8w0OJYVz/yjyT+sCNpyie62s0KKzKATD0UFbZ/XFfI28
HfCBp0AoRZyIaAtyBg9loCCaKPMf7R41UxKcu+nMM2HGfeHXOh+Qq+aRp8Btki7/bZR8sF51CuaJ
RCW/IgG8JbtXJTjz6iVyADp5G6c7CCq87TJYcubIqbJnbbxoNRAGwuo9xPY7QB4xxYVCLDNj6oov
LXHMk8LT5CAzBIWHuJQPK8Klmdf8uTU/mrk3yXOr2/PzTYmDQ2v8rXGCp/eeflJE16MKJTcFYOBi
3tv4yWVraVYxL4Kth4frI/1UMGLdYd0fi0TgNPdjRow7xTEFB4bt9bCIBhkZwobZrRtPrqw1dZr0
4g2CVXCtw2xJZCliyq0mFKD9IQEETHpLtc9qZTNN0LvdfcyoMsGpkheo1EcfVbjpIX6LuLt+Dxal
g1w0zn0L/uXzuwwUx5iC4mcgrGBQk/xgyWDH1HjQXVQxCN1oEDwcZFsZI1aKTK04Zd8Iuiq1PfWn
xur9lAvO1vI4ATx1n0z2WVBJcqCWLyeWQKFC01bIQOxutVOUSDNB/xq1WuLxif2IqncGO/N6bsel
poeaJOgsSAY8IdVGiE1cApNlBK7S3LoDwNYks/9KlF6Fo8YX0WxWITwzqiolAl2QuLOgdET+llv0
JZZuX0b8N8AhngliVy5WC1RLhmvi+xJlaDcxQh0XMkZ4nFoPUcchbqcc4avuUfd4xoxVbcdWLc8T
dH5IO9l0eY0wXIKkZct/x/hFRJv2Gm7w+PITtJy7teBBEjIRNf7gmZuD4xCD2CPLY3A/4QJpWKU3
suirvabuXjNt4ZnLl11mFHTfcs+nKa7P3Adp7ahJRxNYh+o2e+VrSRTfyqpd3+0tHFoFQWRf4E2t
WQ46k3RBdk3Qyx4WD3FNZ/5gOlju+K3Gr7eXjeXYE2ySW0+3PUdCbJrTtGGQSgyYVY/EhmM4BsW4
hgDuLsp8OFEaTngvk7fLegt74i2e2c1rxlqP05uaUVOoLAObaKpc3gDs5+q4YEQY52gevjuf+mD8
/Aw4LkzXfKrmW8BufFN9HCvEEIuGfsvHM24IXkGUNWE5Bk+OikEfQTXQ1Vl37YnVD7J/TKsTQaPn
ahiYxVbkuHUmZKAICACm7M8qy4tjqqLGFeFjr4vYmXvgROOY89S+PM9Tfc4IXqGtzlbsR9+yA2q9
8LkPSWkqCHDaCOkH47UoxW4tHD8wIDheqG/92AQSs5KX6y9hCV0htSM7e9mlzvP8/2GFF2DdFydP
i1dvPzx3LpIp3jWnHF+ZfQ73rj4uvGVTD8qjNfqmqul/9Sv75VwxKswPbYl9VQKYObpnCFP2iwxr
iFHNd3FoP9tg01eAeWYLga4o2UGzqVVgVpUEhYFbCIzEDmjB7UcIM7Ne8yr0Y872Bt2dUXNGW//S
jy0l2MEHT9GkrixAclHJl0faTiA6maqrbktoIRQTw2HOeM5rEMMxEBBfRoFRnPmQMjsGqs8ZHBPg
XJ2XuK+hUJtzDnwdY5tIkwbMaSciJJvBZARm+j+UTlF834KVsu397CxZvusjrkmEVjPKjaxjflv1
8qVOf9mq1q5rG/Dk3mEw4toEVurzO+H+Mi+DTbBISFPIMooMxJl8Qa2AInQ7gOEydt/Y1pJMAU5y
re/N0NPlO90mPuauNGe3LMhmyGJFBQj1x+wSvoIGlGj8ryTCxF5lrWZ9pdn0dXW5PTDSvofOZytB
WHaNr3AM/EE9GMwArM6dy8hvivbYe9t/3M/0ShwIFTtIGFMHsyUs8XpPmIdcstEQsMGCE5Zpmg27
WV2CDuFPBHGn5JiMPXvr4f7EZRQ2OMNxz1m7stlIJfOv4EdS6pUqVN5/gENBLifdmS8XLQOvATn3
PHcQ4DNC2tpqdZFvanARDp/cWLYWMqFFCukMaXPJLDyhgZ2xNVZzRYCaBj8ebHf6tVz3hLwZ6T/o
Ssh+b5UhSD3akeR2AM4JnqJ1pijo6PNCgNE4HYXcInQ/tk1gEN8KRTe5qyKMsrPnbDMVysStsI7w
BnK/KeLn2TfENZApy62VcNbwt6yK4xz4/Av7NkAwoMjd/Bk5vHJRRCPehLZiJSYWyQWjZiDQ4kkQ
efA3xnPVGGwsiIMeWy/Ugh+sgvPpe2ey9yHP6qglQ+w69cAza01MW1gHX/vZVfanzbvmWAvKhd7q
fgsAC+pz4/NT/Z93tmLf+6qkwjLXmJQ9vzvnW6X+iDLx0Ol9j3cKgbWnmXF7CByPt3h9nuCZi9wN
OhKd2wDxs5qeh5QEvYcBRjGeqyESpt0Xc9zJgd+DBdjaFLd9gSrI/36iG4YO0rnsByG4utY1LZAI
dlMf6dYn54xoX6Cu5xJVPeAmhMbHKiqFPx8VhskYM+3lzAvsEGL3aEzUn/G4ntcHmoERGY8n71YV
UklWTFsoF5TrMwPTnu8PDs2BGC02LXcanZdZjb2K6NZv5Hgu/kGHh11uIPqGJEShdf6RIs4/rykq
X5Wqo66bONvLd+xqrWP3llcfyVjOiKw8Z7Rw8VtZudAjsBpo2ECUh9fOgntnEp5rLvoPAcsZYjpe
iFHvJ3Pgk0RNBtOqrBI0rJLqxfnVbpCDgEv+Vdl4rBxiT4LBba6gb6/QxMYTUSt6AozXzgO5Xkc+
/yP9ODdbMlqeC1445/yP5vNuVD/P/er1ywIkSygObbUakjoNzaBviQQX9oop1/nYku/BWPKYcM+h
ieCfbI3uxgpgCBKfl+Zw3TUVu5YT2z28jcparOzLNP7gLwKjilo9qkLr1vr+ERdBinWvM280WeBZ
f42bix7Ugv2APhk9tusaP7mVRuR7G5vgFH96F06SJ4HoutDKOeu9h29sJbycRJ9YWlQ4/shHAmLZ
E+/PGXBqEZdwAC2eU9KFWeYoLC+a75MmTiqzV8EiDJiP+XSWZMu66uPEcZfLcM745rCZv3mdw7Uz
hmsbwCSe6zeeiiY1aWDYwsK8bAS9Jujcu0AideQYcto1j5xZW0RVSogyOy3mHofcqnaT17CKKMnA
fpUrhP/WgEgJPx1H0D6zr4aKJnHUih6QTvHA2/OjDlgyRPT0NaSyfoE6q4EAHZCxLrqW1XYslGVm
5O19SwMHExMWKxg0pg3NdRx/z/VjHEiH25Iu8DO6bQKH6FhLutNjf0cXmEnlcSqce2CoNfCKgS9o
tts46JiMXmMrP4cVyW9Yf2sWoLaWNehTqll/2iPzlf4L02BsRf4Sg0s2Fm4BAJMtWsk412+DKfru
63pDNN+uR/GFeTHVTGBUFdVdRsqnCZVwCv4aEGITKtEc+MKFakyTYQzEBJ7SvOJfQXRPpVW6Nw6A
38yhCfozkOtC353IYpsoTcHenWLMMz2sYtNEgxMIuJGaMVWo0/cksFsKCfsSGB8evrDBP20j50bA
vO/VPxcy1FCK3eX6mH1L/iIbDMDUmoZQ5MjRC+Oza+A9gzscCgPcaxpb2GBVYH9B+I8cJh63PIS3
6lNN1QyyjR0WYmCIkhAS40ED1Qg5n/6Rf9d4bWhAAXYzX+NnRMlrlYq1rJr3YO7cUT6kcGmrPg3m
iP7D3QXLCj4bmBwQKWVu7XUQVXNsfD5sd9ezEF5cRGWsEopAtr4ex7oVuePuzZtJV3PMSdw1ulUd
15pLd7B4pflWmpdcTlS2ctAf5Q4XpaHPe2cK7RfQO4VfAUFa0RN0Vbc6wq19s+Xbu8bCOAgZR1vW
c8wSpVQ3GzFkSYkWcHdx7FI/wwLFPf8msy/gmtWK0EHtZ2+uShgZVQYNAcuKXQwqP/CYTLqHxt2W
Lxi7cuvkb0o2v46lA4HAhLRnmjpTZtBnyFXO/KLxPSjSvb0JrpNa8MKy+LtahE7pOBoI3IBodpOj
xUlZ0bFguHnjqgEhpRb3v0j4OQrFTSIVDuzOH7P7xz71w9HEUW+9PBimCZGh5gD0SYIOb+q2irhH
9IK4yw88svyACuG4IsDVYOWG1PVitKvRA+muEIq8DEQTg83YZS+obIcuLAJ/PpuAlA+6/TuXha2j
dspnqsraA/o2eXbKGdOsohUVxpvB5vr0QQ2tUOjduS3rGnXGb1e59U2fV0a/Icb2C1tEIS/qGHQJ
Jaf9LGLj6W2Z3MRkMBS0XKXhab+fkGXiI9Qc6TXbUXDny34tvsVXXP4LvCEQ4B2z4MKC6tIZfsbL
76KrUG+tBokJmzFew6aOJ++H8+nfvLCBIcHmBh20w2BWGjdiuQnoyGOLI7457lJrr8WMbkZ74D6s
++YfetQ5bm/4pRAQujHVsAkLdI2S9QLti5wsvLKaOKHaFUaJNgJKft6U+DIkoNYWwLNl/SpGNAu+
zen14FrNMUG1ZXuPoHtUQhx9jmEjILwHPKQnCXjHHhViaUmVbiQTh+IYf0gWaAdpw+dcjBDjwIJY
b/b/cw4pV/Sz06/y19YXrBOEUve9XEe0EXoUQTH0Rc2p+699E92EiN87y1957BXp6dKtHv4VrJ7r
jQHNl4O95SWcOXkfSDK7ceO9AtmMwADDlOzck2zFWeeI49+XNkb4CCyI6GIErw1nz04VooSC5tcl
TDrGjf5jYd+Lqc71OjAeqTARXWSHZMDPDNmYzcG3sQIdMxD1BNK+wO5sBDz2DjS4MHO3C8fS1+pw
tPB99LQNs4NLPYIV/SUWlqiN5cFIZGBh8S57wldsgzZPj95W2MpN+KrTLuC0aNKjfbnTcmALAOaE
w127PxYiEqEkm1kCojZRTokrNdwLj3Aw7mE2zNbPVzk74+OenA5pIP636xF8ZKMtDL5ZaqQh1I7p
Ph/uuBZf7RmXG74KqOaKAbiCv5FoRFaDeOJW7Ozll6/ZXz1DCCn7szeymq5FalRgn6czZDy8xDhS
5jy993odFt/ov6eDcd13YBYNF6bh2MvTMlSvQ7c6apygFcz97oGnDqZEXjToH2mplRatC0Vl2PkH
66wgHbbqGgTy/QXJbyFIK2Iq/QHPaF1UWmYtcajFTV22kUjIFIxyrne0yIB7V+GKjpPoBeLHZKqL
b2pI0rWAj9ztBzPuiUJ3eC0ODbzrLbJuxoE75i3WyCsl4VF+2BEo8SJh6VrHL7/kcQyBcMs13NXt
9+At62xWijs36xzZ5FKE67h8jqSDNKXcz8Ncyl6DqCDCcakh91Yeys0IgVcYyvb2jRE/eeeR2UgE
KSeUc7aY4BgTkmgZao6cv7DltaErPSj0iI7T+wMwUELQSxAUM6lmwzZw6/TnLACO/DEu82pCOK5a
2kayjs8P6hV5aG3EgAQJP2oX8ItJfaqKOo35tBDoXjRAwY958+WuzYoDY/lfN6dRM6nIYUnHiVoc
v6ExNPi7wQB8ivyUI8BHbZ9mEh7Oe4xLtVfUfZLm9n7s7nu9Q5fnmy22QItT5VnqqsOvPqZ2x7N3
obPtIAdWfuOqqwdRZwlk08jKAMpqgHngp8djJXN5VPyYzTcdtjyaMsAY5GMcE54K2ZWmLa/E1q2R
pU7aOitzVnPemsb8A/aUBR4odRZFitQTIs2To0/fRNctFTO98JEaeidkBCjScZp93JRJmjE8fom5
NE67MtqteiVlkUUr3EDzwxQ/XYlCkIZ7mQidO+2zfyHVs7XcRlvEtpLyBfsh+fW+bdXuexEsE/FH
xGVEIT65oUAnfzemWyB3hyHfR7FfobUV5/nPU6hqnksL1Pp6amRNVTt+Hn96srMEBtlG9yx5Cl3j
iSHTYdLPxLygnvG/fOOHvqZdva3Nd6+xdJMF7jf8d+U6HJHR5AB2L5LjzVy4JkHNhGfuciEmw/VD
UABRif6/wIekIF+DrnvqHvrqnnctiAz7kLaHk2roDAt2NDf8iz3xF6B7aVEZN7+cGxGJfeOVblXL
HbHb3ufjF7w1Mw3QtPELvJgfYXrLQSOBdlT46TR/0hkIKMoliQcAMKG9fUH82BCsIq2BkJBhuXk7
XgoIaB1oW4nPFnNPwIm0yRtmEh7+egzqc6tA2gV/uuMdHMJmvYJJx6Z3YVsSHgbRHwnVTkzJBVJ9
ceafoGb5gq187+Na4HWkmbwZJCCk/xIsCre+8OVHcFGZbFR8DyVPwXLoC1V9z6utgh/QQ2luCai5
S6uTdOKSi865ClIT46QB4w7vtec3WJKOFoWppDUZC2jme4i1Djk2OPG4HtFPNNISpHUNht9kKedi
ZBT7vefKsWCMF87P92c2zpN7Zm3A6fRLV8yQmZ84I7RId6yrooq2E+rt+3n3GxAK0wlBe0+C1Xpa
gQK4NUAvFnk3CuzePxEaFeyrS42iShznx2ngkkVe3ggLd1qTJehiHFMbSmBTfifgIoX9eDey7b4D
HdywqGNxmCkm2d7CC76CY6P3c9logDdrurpqk5p9TuW/QWdmeoajS2ZoLx+mu9vcFlla5WqLNXNi
mTjrq/kcFaSt4yDSEvfhTAgxGznMq9j0Isn3XeRvTJQXkSICC2fWZ6OvQobsCI7hlXoQ19wm7sod
qTh20bqgxqbrIH9KDpmt6Vmjbd/28dH5hvPkJViDTAOASRW2R9Q6TkQBLUnKKi4OiGgfXwSX1Y4I
93BmEBDI6KOBEeR2gv/2W+9E0wbST9gbe68VAsWo+yCys7smKWOu0cnYoeqp/NIAIOOwuO9WO59E
ekZglfPZdK0b6df2HC0+2I6G1msY8pN99QXU0LGmbkH3+vZuq8cflBmEze532Kepvl4rWJ/TJbot
1qZl1NNYDwT2Csih46vnX/lhx5R6JVtMYiH48RJquHIXU1SyMhAvs3QVcAbNdmNA6wrJmYqscfjd
7lLyf2qkDhzUFWkSX8p7+Ly3bHrOEXFSsnJn8fjruX/M8iASWVgxn/QxZrwdHwMpdIp/6b5dXP8H
fI9HEZ4CWCaJbXtGE7XGr3q56zzqtvog+RA//LrCoz2/5oqoQqLOkKqoI+bVepRDcDLLwfd5i1jd
EddErWJxGEvX5YkMwsMXdkFau2ul2MwW2nUbZ0L+Oopya+SYZh2GoOppAg3X6UaXWezOi+H147wA
3ikprs/jMnMhlFQKsH0BpwYl/1cU95EtriGc7IiUbie12Ir7tVvt9ZsgOt52q3HijD6E7AAOqUur
rHjoaz3fzT8O7zv2iwsIg6MhU2K9jgP+fUoaqmS1cs7+XzXtOWetzolsrZW6/cfX8jZV/oQyoRa+
gxwBLhEiSJmR6l44lK8JufEpWsM63zrYoAhBBV1P+CuWTGZY1ZfIt34FEGCLGmeKj+pbazLuRWKp
SEF6+u5cipd4WhRT+2CcW2nQdltzY+pxVWPdBadEb+muoMybYxA/++Q7a7AeoSjcnZy4VvJb2bhE
wGzLuLKrok6e0lHZcRn+MnU6AcaWKNi5DEhyEJVrefee/VT4f+9SrVCmRyDDGJ6rOsPfLPvpAPlu
9vxeWl1HjdLexVFmMLUzkPjBbMAhWv1ptOHWqRAes+CWL0uOdCyHzpUYJdSzYMqh5PzownHgkynF
JbIzSZKeSHv256Ylx2jYvlilRdUpJAHZHjh9J2tv0v7GGguqLLxp9n8fT0yMSnsbQKSZiJfFkDEw
Vh3tTg964I5Ej24xXA5SUSeREzTssiAfk4m6/esYPrX/VZvHXaCs4nXoXHlruyKc15+TAg/+BMJC
jYatFct9lN9Gx1dEzWvUOvyewoh7DKOaA/cjkGTrcyRL3C9hW/fdBHUIREqgn/e3uiTH0ytoIf5Y
AlehHyn+heyoB7vg+kBp+015p+0iO8eA3jDrYQB+7C8X/6YDr0H6DMJaNVGpXncJAN2eVfzgAfiz
84zVhnbzWlWQNasz/o14R2S/v/FbO/4whTKrUDtiJAKuv9yzhq13Hcbp/zCq8jG7xUuUmJiFARWV
8rtKAGzUFqo0aN+oXB8x0Vh2EP7zwiP0EU9Gdcu0dztsMQdP/VnTopdPVrPRs0aM7MJuyiHqEeFf
m5JEDa4JQAGdm5pw+OPxm7eMOOw/Kb7EhqUn8p9g41RQnTK5UeGERgV5cKbxjFOEUhgELi/my69U
kX6omQBcb6/vPhjPCig9jsUNb5JtOQEEBcCINKJYrUvOrP/Y6xYAAdhDGp5OSCQvUnY/Q79Lwqtg
02D8UlEvX++AaS46K86pEWPZEQRKlIok9ryFuk91FaxCZh7nrN+5aplwyPA/Qtoij0yJE6csFKZS
h2QuptN3QC64JPwk/AuyTcTZf5ygaZi6MqUncmlSrNqFjEtOyii2ljav38g7fl1AKAtIgQXiR1dX
SXZRBbPqWdwRlhy6YCCxSvzx+ucTbrc2jlmhzk0pfABto7aOul9K7fhoegrSV6DH2ijJ5t81uxfu
77yO5GBMu4WHblamBKNqFCuhAgDzab5IyOmLFMr0NjMcMtt7cpSJuhLSlZm+sR11177cXUlvltg+
eIwsRG9yXYEZCUEtR7eCdtrXy4PY/X1IUKkYh626z5kYv0xrHH5LpYHpt43FMVxI1FzP63E2S/Wk
FxnDjxwKv7N7Hovi4UzzJ//6LXvLd+7T1KYzn7tzMNi40lZ0A9sRW+M+3Zeb+BKQunvzmgL40a3T
NaLPq0rmBzwhdbU5/Ab5C7RTRz4T1jxKw3TqRAf/ceaPtlz9kHMb14OSYJyBBmWYwz3aWkKXuqWg
bF24S1Dat4MUO7lWhXOCre7YgUvaS0sD1sx4M/YsK8f5O5RxeT07lF0MZiK27mZJqV158wISD7Lq
Pjakp+vHPeXOuMzhaag/BFFaoPIFElFFPyhhitGznZHuQxd0URDbgkAXvCFHbOoAwvHV3SpsSYQf
eMwXrYzysv0C0MOrnNH/W0/Ai0teOLef8mimKPGjw6/H74WHZB8f10PlWPYu/Zn7wp7fAAxOgshd
c0x5Ou/h4Mr9/vvLdYj/4u0MLmjJIZsVstAFFtmL9dwwDzwu8hJha0yJEIEzlFQPD7hhAeAzT3g5
Q4CeNXG9VCfyereJ2qPOL4DTnwbfgGOP2OGe8V8q4S/87fcGBaX1TgDiI1sGtsICAGiOLdGZPxGZ
kXplfNNdwLPhkFpEBjYz2VG4q4frR8aedZj+V9Z+PkHKQLmHlL4QjKUYuijCgftGmAZYVQnt/QGk
2KsgrUoiJKTSTZS4zgnqYJKr7hTX/SpvLRi1+Ppito7ilDRdAl2La9SihYG1Gxj5L8aNzjBcrohD
1uhg5tAi2rFlGZhDG4bi7u5S+usGmVrGDw4ph2j7SXqTNXHUkINnhYVB08coUkwLBdQlmc3CXVUs
/hnsnLlhk2PaJMKbr/wZORSpamxQJ8KDW73IyIaA5zCHgA4SGi0aw2yB2pdSkZY5lI7BOe2rDKlU
VyGavifjDswjWtj9Itbe7a40pInHvdGO9mo628J7wKdACCSSvJupCHz4oKyApfJCfhnjEOe5uLbS
kfPOsc9NTAjMi5ktv6oyULh2pCdNzQkBvBBCxqTw4UQnlMFEaOipRuut44lZd96QDso71aZD2kVV
XEzgdUFuo3RBss6lXq4YSGaV+xZrVzTeekkjJgM0cL8fkvdEQc+M0KEnbH9KMJ5tSAargsvAM9P9
UuL4a29hLe3cKnE2hvXWNI3LSGgXFoHVqUTuqOchj89Aml1Ca8gq2/yAdeHJLbDbWFXB0ac7J3vf
oStANuXFnzTYZEAF/IqjePfWA7YRf6Nf8MLy8AvmOV1WT9C4OBTjNVMSnDdE5EsxYBQRbWpSWj3F
wD75GA2aR7a0YLWY8ZfhaNhHvDN3m12cVkOqLk/6szoiQrl9UFFQKlI3bwCoL9bE4QckYfKkMINq
iJ8Bp9wLkVAFdQFsCL6fYfQahkIllM6W+pxCJeePFqz+hZDTaOeyQvn4xISOcQJPYa0ZKcgN6VDJ
i4iZiwsfAreDbzPx0REsMtzZD3qW+cpvyOSXBBcUhzrBonQaWbkhPahQ2aBl9Iyy8QBJLTLD4aS5
/VcDk1uq9cpaWl6MzEkTxSznL1XJ4CJe2Ht52AKowDEzu88KkxpxeE912PZFgVeaQW0KEvxO8fum
CsgUOnk2N130Y9Y9ig0x+A2CrIWgKl9Y3g+Xa9YvOxVeYE/E4/c64TfV9Xb+L7I8H4D39xwG8uIu
ytzvR3QjgkDeebBGEwX55gSIHL1qIvZXDfsAmxDr+H0Flh9v3oMZd72263K0geuUujUmjX6MaHN6
16VEcRMxGXOUjtRXO1I8I8dnCxoYe5X6osYKMImH8i8S2E8coGDTffTkvtOhn9JrFcmaLd7Nru/4
nc2bEMe4t8nYB2/WXrtlhuNn7SZXA9Fq6h9qtHHMAPtBEGYgoiNgy/Ahd/PGyqzx3Yt+mzJtFaTz
sGfs8cJI5mhmLbl8/MT3qjqcqe9HYZFEz0SPMhMC/L/rqrzPDnQQuYwLOTtm9o9yBMpnVck5T0mC
vPfncXBAHKOArSq4vK2RQ0Ds8Vsl18vKwFMfkPazuC/IYSE0QPRJeM5NkJj1UoaV8zAu2vwsjnkG
/a2OCJ9rulr2JmLyxbIZb25161ravcLd7sEqAuAxM0+eBX3BzR/U3C82aXcidZMiOrEJQkhCIALa
Os78YIvt8qILOpT9gaSEBFEXFWkM2QR/oRllvUD4TbDwFpSR4OP7NtamNoKLXgH/+LS00/9/nI0r
GoftgzxewJcQn0ARHEZ44BrfPmNYt7xRfgcJxwccjPrk1uzwNbCcJ8wlk4MmOoEECNps/FSnrgFH
iKAm0LXPyGPtSxQVznrOBwGWE1lealqrgnNbZpJnsFCsLTumt0hKbNzVf4wXuVUO9IGHwEWtaRLj
JgTV2XJe0Qa6ceaY2f7MEeuR0ZwO1VoWAZ0YWRCOQQyaGSpSiERYBREViJ0X5Z5SKWPNvt/6C2iM
ZrxSXf9YesAd9FPcIQFIbVjuCxozIHUuATfdHRK8W+H02BTeZFucZHh35mUrowsewiPJXiMBesHd
sPqayIGaR0G4192e9WweDCLlw/JfrdoRIRZkXCHcNTOeFUwaOa9Wixyqvz3JZR+uqPqsHITPPOGL
kJjGBBLyA4WNymhRNJiAra37UZTa96vio9LFmEWU0mByO47GiMkffkHyAit1EJYgAoXFz7aHY0hF
WlRnAgB/QfZ8dTE+2odVhPWeVq4dDhTp9yN6acBYo8GF6mluZNN9Q2wcDZQYoPp6184XTQpkjQyW
s50dVYwnYlGfEDGWPBBksUbWYYO22ZCa1+Hky5qww6aOOp8fyW4ZfR0RqRKy0d/SOLfAckv/coOP
+aBAhjQufNZ5iWz+GMXgzGM2gVVkOKqRr2Aode93i/+7I1vBEvpyXRlO1FDU4L8QxVOxG4uAHxy2
vChJnnpbuOtFmZvgalKZPNFlFBwgZew9DZVrm4yGulqvQpWimtmEBpmExc4fW+qtPHRET3h2/DJn
zT0rj/xxvcmChjX4brQrsRPcIZZgR5V9hMNaStfN46AP99q9hfqCJUljdsjSR0JpUui+La813Ztd
7TwmyucoEsEPFVf72DCXbRTrLltQBycwpg1brHmM7OGfZ5ej6bE6zmtwMnksIhxkURz76TcliXPs
81EXmiWOLeFh49B2B9rjkqSWc+aGCRdA3ExQRdq5WS2McPyL5I0Wq8Ut4xTJDUa1CSGruOW8PEM/
2QN5A3/IgkuzkXncjhhe9OkxceH79p67iEu5NPvkSGIAsBSXXgqvvK1v4cYM63gVWGtBB85n5bKU
plASwT3Ws4pS6yvsHAan4tzbvVP+WeyTVHGEtWjc9JoQR7Ib/QO90R0bUMPwVyuUMItrJtJP5OTo
UXW5H6s9XBVo04JO55sZGSTOxXD51jeD/NRb4NeU67ktEfohnAI0C0JQft9iW719LCq0MgOL0diK
XrnahVK/AI5wV3DZ4s8ol2iD5ccFU7tXE88NZcinHPwKkDy5u7MqL50ZKMkK4FuusynaDgjXDvoc
WuB1bnjppd8yx/lqtL2Aocjgkc/MDutYQlwLS3K7t/mu5OmuTwZYHEMKmK8/Dt4rQLkXOCvFrAZA
vxGZ7E3+pTtznXhURKht2oGkWSWsv8+mheE7MP5RvLHrNJhZBWV0jb/uPzwlyL6/WAuJf4B8DCZl
/eUQh4Du1uXVl1ZulG6i0b6ZT47MpJwD8iW6csJQt+2IyAHfucUBCAfbnCvCxGk9qFskgHD9Rke6
RtFeK/VlHCT8J1nHWVKZ246MtftS2EXexajsMv0xtQ+SUINqSWwBEac06SEIfHbGYg/x+ASDXTMe
Wjip8RKgFujSI+xcBbW9a+I663kWJvrMyzvHzs7k91F4pwZ9OO0QVBmbgq47Bz5v4Wz/ZyVUo1+L
RmAKvUaTUaHb0o5oVI1zAUhuC0hIFLwoxdUyQZ/SVA3SWvte9T55/l0ElowkFS0hSkjEG+uGerpa
CW5YRNSV7IHleGMVlPL0017vqfxUtIv41UUhmIYAh7h/64wMYilP/QILkBW7tp96V45HqPfIFSAQ
mgTAwcQ6S40BeQiWYggZVN/L+u2OUdqJd4zjxZzj57m6vQAFmQW5mj0+PbyUTx1/RPr8DjDF2JhU
4DZA5gN+wBDzUSf8DRtQnpOokkAn5x+ry9l0yaHHySLg6rRPkL96POCTckPK9l2ia3ggWo6O4YRu
tMGMfpMp/YKKebWTzUxB+HkuTyPGDtlJe4R6OOOCjO9YooTwdDwYlhR/LmDKl1EwKGbwP09jtK7b
ZU6F/MvDgbnHz9lBJgJEm+qxuSctC2tBrguhVKhOLROflA+Rx64J+q87lluJIwDdblQsDLz/5Jvu
JM5dngtTW3adhbQZ5n5ukn3OrKYomO/vWsPW4Ky3FJ4iXJbTWvb5e+qYcK0LOscWbGdFAaJoJGA1
86kNEE9YQoxfWoFipsviRVEBNElmbcMhHUILOVskF62+2KwKRKCXWc8Qm5p5wh51j9XOfQqrfpU/
7LkFqcguKWn5P3VOQlbQ1Vt9ZJgBLwAzbCHYw40QKFAFs1rbn6Dm+fE0Y3MUbEapG9ki2BgHNQrU
oDQpMjJVHROQ6TEioopWgPE/cQkjwXrmaZhxQ7RBUzSUQzNIp4BudvKzCSEAVT+MHXVyv614oaJo
6zKeHHuYhMoPwekJdj3VpOHEFAAweTIMS3aqEBObDEGTg75lb7SvPVe/fnd7+tk5zvbq1Li1f+NH
RIA4+mT63dyxqggYIuh4n7uhlAHwH0T8+GpiYYB7ZPy/zIHIYu1VUCGxw93r/lgQCCMmTLJocJyB
Mf1U0whRK0+WDaLJ9IODpN29vqhkszvpVjyIXPbdCgS2eIrDP+6G5uMId/mnX2egTzzZ9y7wIdX7
7hSaPjtwTIqTWnfBBYeWK+QHUs25nKYRNyl9oj24Q6RnMYQf36AxDrDfGxA0HYJqDfL7HsQK8q9/
owqYaGAkF9KtdFVSRHYPRZN3rgh8AL1a+4kuYUkik2ybvzlTlm6/kqdG+tctpl464UMNrVfNcDj1
bvCUHp0WdQ+fkTuxlRMcsZTCZCc7xJeT8Kdsu1SsDTHaOaIxUfUAZV3lXUvCNIDX5uY0tgyPcGZn
U0429CFiNUYwGOSzpikj4A2sKHpmG1+hyvuWqeyLgMb6GBR0V62UVyLaB3hX45KVZTTccHSEZUxx
oCt4J3P+ZKG6pGea0QCIEoD5Aoa7EU3kqRFTrEY/a1LktQzCB320mPJBjTGLLDnBbbMbvtXirgZb
itzCzUuzXdzgm/zRg33pEsDvvJ68XMwGmtZjiO2lZEK8FG/ogPaTHFhZBTbHiJi6wouk0v0+F4SL
qhY5BD/JVWxxCt5hTSGTBRDqQwG9eOkq3dQded9nTJ7quNWPlvvWkwwSaWLvAoRr6cgjojCrGKop
V9YpqOOyFXZZcOEV0bgrDOEmzadO0C8a8znLdshbuZY8gGHpDy5oWtgFCOSfmmLO9ytTXuEfmHEY
Q8+NowWEt6GnbD/O5qZ2/WHYmrA1A+uCWRX/Cb9b+UnUAPOdKxHNb/k/6b4v+XV/oDrbB+DModHO
zDOvRYtQzrfbXsZt4SzKqWZ/+/s/ezvHG0e51saWtA9WyyDBFYFhy7gM9cgp5lWx3L9LWbtgW3jg
ruVUpCrx2CmM+ZoQcECfwxpZRjX4yMpxJ9rpcKhoIrEbj0xhwXjMsJbZexNt5WEpA5wW44VwWljc
gHvPhd3y2b95yKDwGQZQ1AvOfXfuK5e659JMAcg+6wcF9H9L2B/1iN4gahxTytKpZULJyxvjnd+H
QmRegZPShh6x+rACAF+dbltwCGh6mWJlrComEhCKZK6zO0RNzhF9SCOlyh4REpkHQTA5KIfnJYm6
kItM+Qa/8Y22qHLq8yS9ukApTPlGlA6saCruiKncZa61wTEyeho/NBUoa9ykDjsA8QD/I2az3gjZ
q73rf8gEoMgAW5DIO3zJuel5d7OTV9cLJVhYY8f0T5JCKcOTamXX9eT7J9eTN9OICeTj2YKJfsvO
N9GIkszobJUYW5dxeR46YBvd0ZzcCqAe0oZMsOhQgY2T5qNpBK/5nHmh6XzStDSQeip4W1ui6yPp
V10XjWZNd5VVdpsQ45IBiuaK1pQ/TVoFFwPTGbr6sR1+MtDgk+zoVp1ROjCsDIKdLIecNNdsHgws
8rw2pqOxMMVffKPgcpvVT3nnTcv45DCXIQsLaWWf0Pa85yOIXFgtvECnsEolX/XLQOd7ZbJdV/jM
puNeMNL+ld3sCKkEhDxM6j8sv3OYaYsQcjnb2LRs/tNgzg6kYi5Tibj54hROKWSapvNEKxZ+z+Lg
3W1Vxb/3PmhvhCDlazUIfqH7+Bbi5pxJJrJaoS+sqDSD07ieoXUzg0SDwP6mmYmcRon75XEjB1lA
DoJoAocTJPnwRwR3NPxmh0GE72L3yMTwN/ACJMfnR/Gyw6FJ2j5OwPYjpc4Do93SZFpIKbHAeLRA
EDvrAQRD9reePAp3o6K1q0XPrhgvWX8bUkKujGngVwCyg4VgzpQB8r05VZsGWg0MQK7J/csTkRYX
U+/T2ncrtRx7M3qbv8aNrF4hbgB4AL+vqOMzlG+wwQA7UwUe/OiUvB3egs2tHxZa/lAq52IV/Y70
k9wypiKgPqYYxVJwcIWPk0jwxXnGd+B4jFcWZ0t+ioZzF2iceM39ZtjfUDXC0JsB4jF3vwD/QcVm
Ggm5AJXGK9F/WkqW9j+rfn9xnWR2ep2lIfCfOHU2xqSVyZ6Fis5r7GaQXkQMR6GrBsUbSCPGUx21
QI4Ykg2mGcVVkKzvC3kFiO8iKg2fNQzM+dms04gaGsZc/y+DVVmwQgmQ7lkINuZh15OVVWxTsBDp
UmwxTdyRQpHB7dU8/sDWsFQajQA0SsxZlrJwom7Qbc9M9aiwfiRjXCAf0dOYhKrTsy8vlg1PJj/H
TBSn9tLCaP/J6ewBCN8I8f86QvzEl6MmXwq9SS53/3zIcuy4S3c3lCtle3dQWnNUfDQvkJ/T1AbY
Pbfrk51RCVHKl2MzN7Ik4rxYc4UF7aEv0grBZbLF6wgb1tO6XcjltUvKr3dT8nelibkCt/DOaubD
akfHW2aBz0VADLWlWkZii2WCTPAjXV4H3IXFYXOAPb4yk2QaLq1MDxdOvcydP60YRBPJ1L9xVzTo
vfy3CJS6tLw8EI/ZaoOBKm3JZpcM4RHAaBD/9OXfK4+Q9bzzHeB1Sv9xP0enAanfNzfT3lmi3HZ6
os95pS7ASlfGUcoHFT5DW6s4cRxKFxvkROsY9p6xW9ONCzcGyFeT3CB3pMvecXtMS7VU2ZnJYJqu
XLHm3ieE+OpfpwPXDUx04QS/Z7OHnXtQxmm7pkbwTtuJGKY+RollaKYF+ppHnGku/IFTaXVzC6jr
QeRroxcoqwBrU5Y39PCsg16vsQtIFaEqhb55fFlRslOt8jdswmIFVNhp3ZcfAyDyirFtXqt+6OOB
4aY1oOq6sYPnV2ERA7ajBlz0OlDgTcM491FkKCvosXsSz1vIRLhshXWnxl0L9SUDnZ4l54i0KV8f
UFce9/ILPbfaAt41p3ZxbRcYjp0EYngWxmPrcLf7B9g/H+xUrJ0TbAufUSpILQ5XVLBIrFOsPvw6
tvILap+FPJLpRnOvXyU/wqS3Tia9/CQysVDMgXWOEH8EotVgNqlWLz+9s43CEIT54aXWxwe3Qzqn
XbxvY4E9KMrioQvSsy6bV2tHsSv0LIF8ACBmWfMuD60/eAnfI6Ng0C3Zh5CCEJ2RmDSkVwmrunI2
zPbuJyC0avpp/lUU7Bwu7Ad5jFTAnnhjc1lHl4bADpoDwCvaDLBIO84jsuUSDsuXbKkZkKHESRpp
aGRIwshm8fvtaZNtQtxB4fxwjnGaa1VPXMivKDdkmMyS/4fxR3R1g4NdqIxFkfZsFCl7R9K3waSU
U/jvug/HA5kTXQCWzdjQKWYrskvbZ7v/suAQLoeo2ca0WFMxqGqGSiZjw+9Rt6GF6pRGVt/0KE3F
NXSsdLUNYy+tCKHqw5sdej9rkCNPdjEd6Mg1nw2IYvTFlXXs1sO1vXHBB82FxcW9rSxMli7PZYNC
ljnFKzTD7llPZf+ulCdOytEVY4k1OUhmD3qitV+NQK936grAbLWoorPgqYOTm+pVyyz8wkAabAAD
DyLvi/NxYK2jYgY4tdwBrSknbCl3ldTXNnZJ9risMnUI6EWFibVvxAWVeq+1p5BLKzWDULwPBUcQ
0VaFUgiV/UBk/MFqFZFbHxgj3gzAVvMqbd/WKygWE9BUHe3Pq1GbofpGQfqTILWYmohced5T3hmz
BXP+Rb3LO30PDpGx112i4fcRt1jiNyZcnomisXySSzVaO71gBoza4/+QqUwKCvHeaBsAGGSigt6u
c1P1mpBFOt2mT9kLtEBFJ37kMh2A0FDpPgV3iSt11dNoGEl9k6p05lYY/zS5VcdQnmCAA8YWIemc
fAQalwWCbnjj2+uRg/CWeVCgBfWoKFD8JaYGAjvOp6PVBl5CStw7E05xo/FHLl16UnP471yIYRAH
g0ITT3vm587zD/yxO0HcwEjQZBJDxSI4+IHfBP1oomGg0u5W485uznGbIcseXSApBbtFsQG3XzAp
ZpZEjxsRpQn8Fuw89gKlK4zZkxHYnLxlBcM8U1C+aVFmWZOMgQuGdMFGstpJ6LYYE47s4iCstguT
6v01fYQ40ay3wid7ei1bae9bv65yxCH09uqE3GLH17JAOaYFPiks1PCj+VXi3W6a3HYtWE9Nehdl
/wDmXkit1ynZCg5yE3agvP6CZmz8kNyfdroSfC+cyzZnt9YYzvxhTbipoZrC7I5o0EljIvsmz6VI
KZIzyH0DYCHTjS+/kITVI2ecCLJxR+lMGrRxd87liEE4Hd22yqW2wTJOJgiam/9ZmzWHpnBi+Enz
xOGAhj7+VbKtomq9E345M4II6tgg4gnahG1y69/eKpc3McDIeLxEK/4oYDUe1oGIVZj6/YTU+5v0
lCyRSYReSlr5Y7VBHspSVBtbL/rZhvyPta6A/EajuCjva6F86owezLpdmc4Z+sSDxi5ameDRU1jK
tXB7bf13e3OC5FULZjUFnnifeeypVNIN5gXZsgTDPAUEfs4GmrSuA5Pb3ihsUkLM5YsrDUCZ4x7e
BeIf3IQXYjCnI09dY5pMvPx3CmZDxrY7//6IfcgzclFV013NCTn2pOVqjSqoBJ4OCCmry4eMCrmx
sZXOfDdftzL+JLPRY4z9GScw1FgbEXhviq8RyJbNcSlGtaQcddQBXmG36ODdcAwlVBAXuvdE/Jkx
7z7d0lKlNEhJi2B4oTV795MVwncmQki2ro9ggwHZ2idIrfDg4YuqaYo/TUOx83BvCycu83Vsc21S
J8pbHOtmX/3UyMx+4F3FQ3EkRIIOG/WHnjIwVN3rZiPOs4+x+IhO4/stwITzH4ecevUWAlrP9cSB
S+35UIxfeeq9gF3C9IC+N2ukY0pqQZ40+KhxGWtQtrMlAccMqn/OUjvtzrGHBQGDKKTp7gD6L1qU
rSFL5HjhxOXOW+B4DeEaFr3BgmQl/7MxWbn4K3YvLplTVBS6mmGD4mpszvYMRoJfB569GiGANyA1
p1bD/OlJXcCfDGICCt7m2DtA4o+5/ZgTJxMUIDlERp1hMKmb21YjA1jC5Ej+9llDp9PQ7Gb9EkUb
j45KVt9m27mkGaJa3OYn4gEIcD6I7gn6s4z5xB+L8c56EgSYuMP0SqadhBOm60zcKFT9LvyPdWAm
M99qeOy3omFhO8PjTwbKqgwdNJ+KIcrVNkoL3MOxZED8HD8fgBDS5QPuD8ia3lF3h5Nlp4aIlB1Z
GY0iF8vNKEmfqqJGY970DxLmU7+dO8QYo70/eTp5b8/Mo1gJWTR4W+DjCZnuMhJAolqKbeLUhPUz
tchRQZWyfRhGJFiQdp4qAyjZeQMyWydrMMMDnuvhgYmd8wwPWXViS/aFQ6sHbN8Kxu1G/CLkvoPo
tHnqNts6LWLgM24Mw8cWbqzeBXXmnclXll0QWxkBrxRV5zWb32sWUrDKv0bkJS6B7CSkFVXUBUek
gS2U37OYFfRHuOfcnfxEyab+6Z3bP5/U70DdjRLQN7iApi6+h6jtcIkjSOshKXOYgpT82VVU5i+3
EWk1tKjmbrkyaNPk6FicJOUCnlEBmB4/f9urF6ODnG6IK9Wqi6GxyJAJ8fRMQgRZK4laGcZNndkN
rXj0prHYh0buIS2rpUGqcBczneSHFPL7M3GBq/IsAEPglflL+TjgM2TtvNZoZdjmqzbxgGmpZqop
HFUaPwTUzQj09DuLagv2iBr36oE8boNT+egCfjRsL6lu5OeyH4nNUszyc3DSkDM/wNU8YjVUhrqQ
LVH/dsS4tMcfRZMFyePExTDwhWZj0l9xBbQlIisOHu0c1mTKlvrCOsRcsD6p9bn54vB/uNxvvtjz
dg0/MO7drdz/LHpY4dc9WWm00AajcDitoCzUHZ4zsekN/JXtoXS+hBoIlmjGSB/VeTCa5H5ooJD5
72uuUhWz+GeCYI4c9XnCXLgVtDK+MTrsB1ix9fCAxVuqd71w4vA3NaeQUbQn7CjhWAI0B07thlB8
7AxUInMZ+sTHrwAE5UqIFwHMuSSMBpLryEnMVxemxaufCPTMUV85T1b+ZaFlQmvApeDUOPiAdwky
NrwirT0dyBuGlToy9ntDi+m/XF+r8Z/EE+Mj0spzt77fzDcCk5ztFa87d11cW9EKAUbKWTdh7f2G
Ch5P8y0llMiXx03H8sudrwNzx/yeqt0JdmE8XI0yDy01T34I07Vfb0760DP55/aEhLSptYyUOifc
wKEeOlPESkZ2fz5IFxdlv31lAczvBmz2v3ur1Guu8yCRkD3pDzsuxwWdVJaN7VdsaWixGjNE98yZ
AiGT0BLj1hqYu7bcAYKiT0ruMLE95LEqOuroJzRXM8K02uVVC8ON14xxHI2UhrWf9S5sjlOXCfsj
+p4eoVOzRmQiCb+Vjb7dlNuxi0p9n7gO9WaDJUUse6OltmRqnIlX5U/0QQG0YuIqF0xpTMGsv9xQ
iP8TRi44srywoyTT3Bt62gAjiOcLCe+4aTk0hKZxKbYb/VxB4DRG+L9vdZ3Geswoe52HU7bFEYwz
jgfUQMO3gSrX9O3uSfdrntOC5TTXVhUo7e1K/UPF9famsub9zXdmEuKtHWuZ16Ugf7YXgLe2GBFD
fAF7RSoGIlECuHStZS/br8nxZ8LPfWv7F7RSokjw/X6dHx7NifArPhaGpj1YbfTqRrt7K+VSAV6y
hli/+KuudRl2dOSwpd+aWo0prm7bv3kupJXYsrZO+yNcktRKNhlYKQPvxJixVKeaimctdzdletx4
xbLr3h5fxLabmQbV4YS3svtbTzOnnRrQKBl4QWUz21wY9OHU4Z0UUOtUjj98QsWUWikDR59u/kVq
NTb07eKKrSbxB0XOw07G16TYdhm9DIKgUWChn77VvOZSvrS/PmjHXUCNfpvQPIcztN6l8gOTOk5p
fEZxXwfTz9bi7sHkl7vXT9BYRsomgZHChfJ9JaJD8jWCzkMgX7wW+rf+bGqBc1KK3xNXRWLcAz1v
muw7pk4/YGQ2InWzludd2nue19B/9aLgYo3/4trG7XFyyWYWedn1Z9gbuYZEtJ6aIwVTufmodhkW
+fsZQCLpyZFms688ZTB/yBmbP+6Vz7Pd7hm20RJorQbOxwunn6dpPzTASznLrTOQfYvHBvUyKrX3
mrd8BmrrWGPRnm4GBtLRWUYqjWDRG23aay+Yu03HQ0AThn6uU1G/4vaS25BocxuNZRHqG60iIFol
9qZsON1EmlKDXucnctQwzzIwQL2yad7BdCiaECjhc7cUp7kucYJMzsLWr1FBlf9LGeCipgUItCAY
Ohe4U9xv1gEWF1vqvLqBxMj9Xe3VsIRq5dyuK1GO5WTbsJ8nr2GBH3vjkv34bXte1TIPfh+5HGme
oN0IMDl08ApWmx8HoczfKTFlTD0xddPcA6yxgizqUJ7QJpJIHCqB1ttlow43MADbF9iaS/nOJrS2
EtjrJ5YJWfyEINsetwSlueS8/fI2L8FGNf7NLTKONjLy/8rDm1A0qtxhn+4pHcmBYm/X+0NDHaI6
CmUcxMw9YlJSj1WJ+cI21Mrhdsx0R/dPqlh0maivGSFm/2uP0f64sgz7mL9129Muqrbe83Opia0E
0E6j0WFqhtV9OHC75+SoHN9+ubvq14oHE2DYa1y6oZWxyURYvSXDTeVAQueGzjPelajR+D4Js4yd
8T0wzGiGOd8/VGXbUF2etlkcGe+2q2dtQasoVzlGU32eGJKU2aiswusic+dAKx6vl0KM0uzqe0iz
CKLMiHqiA1IzUZO/QzBN+mBe3ndkIIs2iq2jl4HxEmBnqX3gfpNt+vZSJSxKyhj7s2a+mrRifXMj
ojNl7F7VBJ/NXtwiRb4UAKCb/8UbyF1GAFwMdL995T23QAOCM5JWyxgIgEdRPl1s1eWmDpoyatlp
ogFPIeNsMdpy1ou86NjVrFoIakTmpZINH7f04RwyTn004i0Fb8LllQ/l6UaGVNiAH57SnThUxpx0
aFtowDwVLMx6jHy4CmtU5oOK82e2iU1ti2YLuiX+Eg2AvaJO/xBXrFBn3mLl6S/8h7r1Cd4G7mW1
MCJEcSToCp5QdG1nUU9hGC0efdWUANm32nx7SEz2znvbNASk9YPXhtEV6KFz0FEJAdFPEorkC2Sz
2PcQZPJ7j5crzV+toycmhxjUq2DKpG4NyguICo96F5JXnG3Ua2clFXeoXb3yioLTQc2SBURvpW3M
SWB6p0i6ukJr6Xj0qiVBG8q9BBNQX8mRUENSiOtS8jWLIW8nmiUlnwU2mh6MPLE6cmegfe5H2spl
xKXx2gWnq2ZJBnjPCZjXOqKX3/JO229JfnaoUqc2rmGijQHQSks6m5ti1I32KcydH1nsMqI/XKr8
27svwnXSxA+4ldrBE0/9ObxPQB2FH4QMR8u9HYRrCZ9Cx746DcbTM4R+OFPY8mlu7rpmroczoF+S
gMfFpDfNbecICckgxbmV+2wQd5GnfBKquGC3GGLYydZGKwIKbMFXq2FbFxV3gS7aN8ZVGDJOVB3y
HC+YoMtwU+Y116x0RnZOk3fZiyGoKKF8/EDaYIX/Uk7/7hXdlqmqdR9DjvXtUAtTKFOjLLmevnmu
BJ/H/e9Q50yPExya9NBCDpFHzp+7I8u0/suEfFy7M5xrhnZ+CoT3AX4NizbKJnURZWSrr5+TzuVN
AQQW7LvxdeOKkqwr1ftL2eRDo6+4oeiBP7Fc/hR0eaAmgMiwc/nZqcf8vrtzMpczwrqavvmTJOlt
CVivoutQO1k8jnfwf+EOL9Y2tp3BUpjIT7rX02gxaYxuwYv8uj3QMVUnk5WHtiUebOnpS8b6YjNK
Tml3Mwrj6i1bJYr0uGMuDJ3BHdBMIDnNLsWn6J6TKdJ9iTqtLn0XWDqv32y/qZt59SZ6nCCJYXS9
K1ngfzsbuhEbNERHiY8KwrFcwQIQ0zJQ3vREOgDhnmqn/xvQebFPpyuDB9IUYJ+H0W8iCJ67EXvh
qE9BogIjEIEx0nQJUu6gTCccqzibkSc6NPRTPk0Es1IFwKuj6ZMq/NOaE4x1X608OiZiCMNT2yTf
hnL7Ypl8yBJOgK/QTgJRJlQg5eKDE8bMLWlLQEu1H+7iGV/MxGczi3nFbOJbOjkCo59dBWJyC3VC
Se4yD5G4Hn+dVVygukjktEGftLiSByK0V05MOs7FNRVAj0w5vOFqTVxCEA536i8IWBArlzlBLYky
eqN6m3OTBAk9UnCnAIY8o97sRIfxPS892sXkR/wJYKWDyvspGMv0Njsg8axF8d9MN72gU9Xlu4xf
IUBEQ2bvDZAXOVIoYIdT+4C24AuPLRv1udvzgBwzuTWc2WOrOWoUpmaB9avFVJNAZ1zc+UFnSlDJ
EgSBBqHWL02deoBhTUaM7MEYsFZQ7pnA1B0lLCk54C5kMOrBqPWhJ+XpUnXwM/K2da16/KELNz+A
LLawiopdAZNmb7tNKNNeqg2H+lZI+WfbnZ0rad+mZnr5TYJ/MY9n41lkwT+D7BXmds6e3e5Mx8R/
3ecZjkmvxlMvkLmHah5BI2gKzKxjFsf+Ct9EAqxWH7WUXU8RjUzJrsDwWuhCHL7ESn1v+HU+IqBj
KcmGcZwZTFI8WpsaHADFsLGRx3qnaH6sxWfc4DurT38+/7GwjdeTa8q0S/OORjpblSOIKI7NiT3S
eSGqh+seKG+5eLT2S4VrZP7G5tk8sLIAsx5oqnQOqSoFL7D/hQbzFrysaIzN/7IM0VdKDBwb7lo3
T7M3E6kxKCWjUlRtFDHEbTldhkU2ZB+Clwtjqkn5+03jhtJOVvv8sg2fRhpXfM44BzVa0usyXP60
38zFcBMuqZrmLXIt+C7LhD1LbZ7+L9n0iTQx1v5HcMvBhyhtPe2SkNIxJBVijBlRwrygRL0pfra7
xIZofR8M3DZ3j3EYqCRQbe4UznTS2+3YfMrJXINsDbcfuaeMj/O+vQ+IK90ToeDLisjQL4ciH0Qg
u0jh345aH63Mj4kyHfMeeLbRM5vGAmZisRFhsbQT47WqC+5BMdeNXOXiIk34GgKxxVSQus1O5S7G
S3yGqCl8FuuC1w2ErncRUgVkuW8zDISTKf8/sopTzsveiThB9aSV4sybS8EwosJ9n4Azgs/yxnrx
a4OMQrpwJEwkyleHEhLEIiph592NOyZTXTh05ExxwpC/vVWIRkjSqCc4uyyRa+zHxbT148EzZ2Oj
yAtI0G0XLRztPme06vaJRCQJn9Ojq/PQQPycYLHGIWJn6xdx32uNzeoypfl67Xf2FUSRlMv1sS9Q
QNxrfRmwuye9qFz1qGLwfm+mPOb/b1ftEQvPMtEyT3xCoMHpXd8/8uQwwYiPiysoHMwp3hW4Mh0S
hxYBLCySWqzOTSDvZAsi+XITnEchTGt61honISiDZWeoCEXxV6X1NN475JRO4pVV7B1sL/iSEBen
G5EgnTlDAXAwCevGHnIEgE9zeJXUq30b3VBn+rnuulj+pa9y89ceqiEyDfuD4+h2AwDptYvayn/A
JmRkaJonOKlnvox0rseEmHleC2jyRTDpK0OHR+CY57ofxGz7dT47QO80Z8SPEcQ/usKcpvHGzGNK
qoAT23nLBpeSEiLURTrvUb32/HWMMgR/7xvsOFeBAaMmV/shvV3cCMB5QIgSNMd/2nb54dldjlEa
U6WDc5NnE5pCa3dkfUd7B/mnii5EsrmXz4nxB23LJ71gNZfZmpGu8ihSPXytXtxaRJ0M/WrUzh8y
z0fnB2WVa/hYJglNKqSJ03iG5FNDw/qdI/+BjTni3IAcpXX2PTkoNXH02BFAXVqN1J128Tu87/Fc
GnHr5j0lZHUyxUAgbhu3tqIHj77ulW37eOk4VeyXemJni+jMOIDhCZZfC2ek7LMUAHq432hWvEOm
J52aWWciGkzDqSq/+x4K7yGEEVajW9L8nRgJTqfgnocHnMzNFMM0vSsxRE/9fkMfXuVZ20huRb6J
2nTsHi4E5Ipb7mkwbtj6WLJa7Pa1KmIrAg2+VhG1QiT5WvyM/eiaa9ouFZ2wnjP1L9EEtjtzMi2g
iQGybd1Hrwyqmvqr68v8vOSCeRMqxNfm8kzPA0rYdezkmJUph3P1MWueKfsomdtX2dRufBaRJcck
ysDJWp7WrdVWVNXk+ENKwWo5Av24hhTFPxcIv2h30a9SyYyAoTsD8VfnR3sCLegj0aLJhS/e7NyL
f0XDtMwwntZLpogOIAXXy/ydX3fhEtAx/jeoLEu7R7H/M827tQokQJSC9LnDvc9p8+dgD/ZuQkJU
MHy9Qsp3hOvlBPxo38vYTSMIMFGNj+rlL6MQHYu8xfecKrwTZuiYPe4JX0o5BT5o5/FtLMgKp2jm
rQIzxV7MskqpLybWfpi0nHai5ZcF4fNJJPTHLBUGLTQxlIx8XYYFj2IWjgH51BdNBUDVn++eLscv
EHiUWRn9K1iyGSc396RVaq+Yc0FspB1gD8p4IsWKIRSXep9SzltRJRobvB6Kd/yG9VZFHXK2DfhB
ZDDvemUQYXFP7AAa11NR/aiwh/htmKKp3mifkZmoHqb6p4UzAmiJIjtEs6QlU/dIKpGVZHZ3A1Ow
vg5AAYqnGht7igXu3JWFhKBPmXP7eKN8DYS9soGMhTGQpa+imY8UkDin8PN7h0y4LS5ghIewVSOh
6Bwxwr8eMPvBf3zH0FzPuIU4xlW3bpzczNAWVvv2L1V8QI2PtwWLU2SZi+lWzMND00S/DcOP7DpE
AyezN6OsWoI6Kgy/f13h7qBVj5kPx9k8znoF2sDXG5jXohmfFXvjYA8pC+gGTmUlDJWTw6lLnyYd
nPs0C9UIfy6bDBQooIh/Nout1uoC3+XzeA6lE9wnWH4uwUNwsiK+lpzdVZ/urpLuM61KsMPouPYu
AJmvEGt1ZPqJgt3VbGeMw/0VcDzaMvZWTmPK2lwRBGMfWgHfsfr/vhbNGmFzoYym7fh3coJ+ikNI
0OiLF+QIfU9vUWEvm/86vtNNiLEG8N0ohwFaw6E8z9Q5ICaRYf/w2b8BFIrzHwZ4b2++vW/ruoOh
2FuS+ESUEV3UNSzB+E7ZLVb4xnEPnj5Ap0CmnQooVz3J5WvdBVgwiO5RQbL7RdJuHfHpECKmm9Hu
eeK0c91PwMMV1amb2Hpft5/LywxmG/mS5MiEf8j47+NB7jNgRRJPs1AedJNGSaSqKwVQjPATWTmI
ggtL2qTQ5/9CHv+jfbqBMTzoAh24IJ4onZt7HgMHbSzoNRA06k8tmYvPpeQMExGjl7LPc9Ao8JZK
CEsdqD2HKO1xRovYA4hbA02OupkfDS1zyijBENKhnRJJF1BT3D8Yz0z+5jilWgG200s5WL4x40Yv
iwTsc1WMf+tw7HLsKqw2Gw6zwYIiCERP9Bh5/jfVAxBvYN7jMU1lyo4hbu4rseEiHwLgA6ABmzxB
G1wRIvoAHIW748uZhqlyEEriUB877bu4nfkIsFu45diz3dlpNoey/F/zAh3ND8CuwVMcoFWfEOw4
EfXfDvaDI4dcBAGpDWwcawunYjHzj+EivEF8i0eM7CS3Jh4AGX+o5AfNGylAUjvai+Z90vrMCmh+
Vu4KgBoNQIy64+FsFK9YJrm+YNlrpKxSyRdKA5271hr2khAoxporHmb/ZkogZFIgfkW+rnCGytja
BEWnKgDXOp/CsbbGVRi0SMpNYZocnVbawpYE8BG41oRFutxITkNwmOAojo6qormFLjos3ttl3KOe
PL38kDh1YCvzWFZk+wsWfUT0STr6mlye9Q+7ngBNWoI4LsN33J2senhFklNR2geNQYJn08PbQC5g
oFp3E0/bTV3D+F/MoQHcKUfa5mRNrETI9iNguHSw2Zom/QgZhsa36ScHL6ELkJ0KWdJN3Gx3TybV
3p9pnyxfvzju2/OSqM6R6VMHeoUajlcrMrRS72vBvUNYzaNGni4c6rWLoTzdedw63lK0QD4V+GgL
ebkIVHtX/1vB2qNpccvc3a0VBsRwRge8Cc0EqSTLrLlCHbS2BP5n9scI1a/kvMbQUM8ZtM39qxYN
vG7Z+S7DJaLgotWXUA6zPBW4EREF/09FLuFbef/JrDvj/d8vzEeldAXpoSLmsukc03qM78OWV7Iq
fJnfb3NDEGB8rxRIRGWb8tBpVzhPbtZ4puHRlG6m+e34a01cxJyC+BuPJ6XQo+/wKnwLVllq6CH/
wETzgGN4mV9YdeK7zuMr0YPP0Ly8niqZ197cLAlAQ7d/qE/G0uEV+A0pi4D6cO4Dl+IJipkbQbrU
VuDkU1BOJd/azxcNk6UG59NeDsl4mU4kK1E+aBMpB7iYBMFcXfYVDUJcQmWE06oJdKhkNbnjWmST
56Ci0YqtHhCeqyLj3CN4PbIx/CMJqm9D8je39hG03kl+83o8D3nAX1Cfle7d7GzGZo+PUBhVjOlP
zqScxt+S/QoQasjcHgtUnEgNQSI7glLr3hObCNO+MsqjfEvB8RuXwiXI18gb+eXLOWnZJVl3/0cH
6WkQLEjzkH0g6OGgByHxdmLD8StoRqbvw52wj4MbtSHFLg6IBRz5t3hafCUZ7sPX8IhxXzjBwddZ
5TK2j1u1+R478Ueo7fSr4eVMc76640yo+e1R8wCbzqyeHszJlcLtBwXBmiPZ4chGhBUuZ6d0ai7b
S0hklrgFG+TLTfFHg0wakj6Fbnm5DEV/TZxLuvs4gbaHBoISpPxkyQ/YgTvL4dx+xRiE4pQs+inx
v5CLGKvqV5z766ETjDFIrvZ0ujcyWiyu/V0pWPPt0JIK6HTvmRJT8W8xzdAAaZlULDUlh4yJln9p
9bxzOzAaH/VQ9uXhfVsa4WBOvLV22TYga5Vv3IwwyF0MaRYyb2DnCeiRBAvCijuv+8LafOipA4Z/
qGa45jMyrVhbLneQfCmtPUXavJ/XWs+8UNJyU05lBS4CpYsNYHmUIWTMOQLHzPxZkf6EAHh7Vbr8
txokJhVugtYkSmDKdoReipJvJjMY/wO+YkWxROFlAhL3gxLohGOvBSvuuycM9noJb0s0KumroPP3
TZq+bYPrFp1LzaReW0JamE5cr0Rhm+wokFufJZRyBsirSM34O7DvVFWKeVVpCa4zRRgYqR5r1z7i
q/wCw11cRf9WAm/xfafzxf4F5+/JeQuoLA4Fd+h9qdbCNGyg7OxEflzMifve5omV71dWt5LY0eGu
hFz9ZJwezzb9u37Qp3ijo/2b6mJjzLvMD1HCn0s4/N1BhxINq7+AqUvsRPg9P2+FaeA6wlpwmH7t
bEriuMjCOlF50KUSCAT+WRnEf05Oo1hAwZWeseXrrtSkHWzFu8Lxc9l7yLeA39DQD8fCuVQsRndX
iBEebMQwCgDOxTFCj7DG1KF83GtIqDu//IKtcUlooZ2yr45AiA2ve3jBtWeyaOuO6QSuSwr5PXez
gMLyrrSZWltT+4nE2Latp+runHGYe6d7Vq890l6eAZPrMjWnOB6apBXps2mVIfI4txi6NpIE+Vm8
Na4dmtcl9UG5QOm0WT1Mh7fRRAif/6OiXNY4MjbMuLkVQU1eTLQqJl8z+KLHursi4u83i4T7FNTS
xPW58NszQmbC/4/78QVFSahU9FGSpZPvgR43YWrtRaAh3jui7lvnGPJ7RUze52/N+J9UX8pD3H3S
TT5RlqhuzkZFgEhCGaiZYCCTb6kgHQqbp731iHUaidl+pYt1gTYXdzDIEc4GhqbM9lMjfTEzzS8Q
U4JQ/cXXGh/6EI+dyEcVvw/Ubgs37fT9e7h2hW2DZr8PTp8CGXB1+/jqtPD0KHMZ/6YgmSQHSYr5
eQtToIbhgJbF7KZNMkPG4h1fxA9kBi2jjdHC9p5AbccWvOQncraImyRvM5WMaLGTnS9Q9eM8B1EO
A89p7taXj0DbiwA13HhakN4FLrPmOWhsvu0UckKxkcQLSYburloTSKrThAvmdljFNkSqa0ULsIVs
qnc/0vjkgru3lunsJqJZeFW7xuCAI7oQg4TKbV5AYf2qzx1qyQqs+CBB+aJRYZSS07fhMxJRqE21
4AXwF1XhvDvvfzUKzFnThL5jmgJZS4kCjpoqKlNliYxZH+FbbhM9YOdLc+39ayZro2ZK6SEEYBqY
FYVV43I4HipTSyCB0vwMtxFhFsU487pKNK64m8rVRIBAWzQ0giQapHYe+nTB7RF3ilhSvCLyct7x
litMbGkETXTjshrD9lV/49p+sXNXRM/JJHM5HXyQ4FWWFz6ZW3md+5HG3xvfof/o3OFPPC+hlE6l
f58VKzYJBWGPy3vkLNEUYrOwHe4cbsBA2DCvwClVzCVioIHiy/Mbp0GaBUoGKvNQEVCHlcVGIDyo
NBvVpOa84RN4QAtqwv392be+hp7j0A31K0r3CwBKq8PXY3TCzW5bRrluipjQxjdCVNn1obZJlNd4
CRf9axLDGBuGwUFNSBCLdOFW3X2ptIqRpkHOwkvSH0uE0PT3D5dIo2NwD7ldhwHC8ieV6nEn5fKs
hQvPmXjyc1vX1DCCpsF3/Knq8mhYsY9eOF52r/yetX1hWV48UibZZxgdUMTQtaZ9Wuoy42fIGhru
zwYLt8pbo7aB5xJa/z545f3VyMM1mwe5hNFPNsFE6rYKfOR8kgsrmqtrs38I8YOHNRULIOydjIsM
lfombC22rknwIkeryT6GwjIjLnupU46irCy+53iAqJiOkbJMQe81a2Kowe+/BHKSr0z0KNwyAbnd
ZFVppjkoHR3vEnKyeTv5FrE0Uif865FZDiVMEUlzvcVkOGhRI8bzK2CyxHGAsDSpcdmuGNY72FMJ
/fYouTSNsmfUhRTFcHhUyhsYHi3e9Ikpmfxr7r8x4SweiLiVNyzhPqMtCvCgii3KS8loeNCvDleP
BsQS+hi/AKlW4plZBpg8e8p8INdSRFYGQOT16YM4ujrVK7oOZmEiN0ICZGzscHc5zsQVnEiojTIT
0d/6+41wXzHzV16ae/19hN8WejIWBtiJ5S5RQZoImPwZZfVqWUjfuc+Xl5voOg+TsmQWy10pV65A
yfb+Gdn6FjCA480VRPM4BbUeDp7vKuuYWuL+OzUdyBviKOUm+Zjs5kwi+ChTNkBwBPvoOavrZVAM
J0tHk+b6M+dX18X/59B3ddFuoFBQsetdThLn4un41v8F13omWEvWPfIDaLqqR61VYWSwe+OFToVw
/OGEYuU+GfZvHWIliMlI1myde54gmwkG8gZx3Q1oPZZwPo4sFcjsNJkCXqW+n1474BMBWw9bbwb8
kEu2jkoGCzf6oxfWXZhO5q9SMnTpE+/7I9w3WdkEAGJNp5W3Gw0dvxL4zKnI0d+WFXXj958zRcEt
PbWgL1Vc7WPJskKB3HLDlh/5LTXUzxquPifMhp12jU8sHWAKdjr1oxx5nPmafPUREIUeNL6msaca
sulqrZLWiGPQQYX9d4a92xtJQ9VR9r4yAtOuVXUiRYzPZfcYC658jW6dksWw8YvXzu6ZgjF0WW/S
w6IeSP3m1DvqPgvOXhLZEo59x8AJOL06fMb+gU8TJlk/czMWYEdrBNRfOhUzZ2QpbdY1UR6YqyLd
FKIsuLZofYjDdFN2De0qHZ3EdyUVnv9KFe6jxQpBBJBdkvyO+x4/T0M4k47ZSDO1P675DoY+LhtF
8iOkiWUR8zHVjxFiQTNgAWh/xJDn28Qacheo4/pKFMY1lm/UTbcxmBHWUJYqSIMaWG0X8qdl423s
7NDimBEwi5BMBGmMHEQTy56bBtegbzIGBfIT0NFr+5I3fIEYrZuTaicRbEpenKkgVaof1z2YZC0a
2dhm7GMgtCJGbpFra0L70HtMQq63oEM2J8kV/aSjwyUAnTVAMHvm5mth8Osek+IBPpaqgwERufgL
Xhk2lfSmXJOIa+HHZJip3Z8qJaXEr7+QfgB6/AGMf+F9i7sbRiuHgg0ru9GJh0+4PklN6oltZddC
T7LVlmRfHt/+70dlYMsZppvHYdm4pFPqERy2cx2t0aET9HFhkcDD5quhy8Y4puj7XblnmJukFrM3
B8hljq7zvMK/JzCkdfx2FBad3BbhXNBCvJux4EG4oF9lW6M/mpWBsB/vpEezCwJJbH5IJjaFv8dw
bgWGRA/a5bKfDvgSmMlMeOUtwkAlTcTrX10sU4pS5bQHMzYtWyyWKhhmxNLRPpaVzTljqc3cJ6GX
hcNElo7B9qRWziOYKLo2aEzLL78ZMM8EWVZmcYFDlaSZMYufafGXqW95OKhOcMrOn7dFCga65rMH
xqykOzbMVNgD9IX9+4s+6WrIZ6dI29Wgy4uAkajeSLVPaoDL6ji5GPi1PRLOevqUsr/2RpLkxDgF
7S02YyUerKvcnzXxKlZ2mZjNEXULvmfB5tCA47XygDSFO2LvTdBwTBtAF4mfmJgMhPBV6SljrdR4
rZvI0ZTSPoXrtE9f+q7tMNtF+nVPGW55kiZArYHJo71SH+lpLg+Rwj0nAuLGtPIOuMxQZBM7XdAY
+HFlFVeSOddEjdcAmdq3TbqOyKoAEa71xo3kNew7rz4wI+p6j0g/ID6emgjzhZEVQ0qT1/SP5mwW
cANq9HJ4iInNS86d5+8euhySvFP8oFlCThw1KkJIRyYZ+NP276UwJ96G7NNUTLZ+pFZrzaa7PC3d
FTO9pMJ5lctnTmYsSYl9pNBvbJKylYr7oJiiEp4+iZa5UwbVdlrj04i1XE87zMMsLeW4ugx0mikd
2umtGmS3FjP3Arjo8Zfhrl+kfWOGHPFUO4cnWCu5+EY1nrIZcoijRgtbJ+vw7MC2chysNfLK6mQi
4ANovC8RS4aqhp574NZwpU0HHFSYLZ+ZQcwA+S8RV1Jji9SQCFWY4gifSijL4TlnW7nYfHIAMI2/
dbQTMi058fBGcCckJXtHjOD1k+5+/O7/Ub3GwhKFl1CzsE4kWydO6NXasH2s3+2sG/XFTNCjlMtj
QaVdHCySlpTqJflwKZlsU/XC38DP/0PpAqXBYg7AIouN88hKDXCCYlovPRQEiHGdDsvF163/pCym
YuiM6zJ65JqrzZSij/X3mLIeBMo59k//5E4778sonmVRCBwsjUeS2/7T1AwHgCfNCR/YO58IPWod
5ifJbVkVgvx83BvGRZXZbWUFy21yYA8/XiU6twp7HTy14HUPVCYDJPCVML4QbGPIqeTLIDzlJQsZ
ZDdPExpbGHJnijjhgmodG1I4oih6PRvWuDJoIIGOFAwHqfiaTG2tjBWglkg3Bx4zsbOTzXoElUjS
7q14QsgpJZa/Jii9I0H9vreK2mKzdz3Pc5d91P2kdghClZT6Gc1ix2mUpx5jB6p/D5pbOD2Yu7BN
TMxCogFm+ueTkIrbQJX7gmYdP6ONwoumtFHdTMQXysvO2/waj6zsiAQdXESxETWmpTrlu18byf+s
7+9/tEIHXmh1e29sjGb1OIw1PZ5vz3vhd67VH7GE/ebCdNDP9tmikZMfMIdCm0o1x+/O+D4Qpw1r
AauO6xx2FdYg0vVusuDaF4tsehdqp75XW8vfUyxFB9KYFE6awWz3JpzmkJWKId9M7HceDy1w0YBb
7dWaj85x4u3d3r3mvYB5wn+qrSh3UamHu/zTqqC0ocqpnnkTaKsfWZu692hNIESaWyAr34ccgsoz
Q31uTEhe9ZISQ7yHp4IpS17EuM1FxEiwUCCDd6hGU0ZV3+qTvdKhR543MCeD4rKuZQK5tXAuIana
qPdvvysVz1ZLbTT8Fy6FirigTdWRyrc5cr9aQhbeCZqjJUHoIkSA5LSQ4w7MWZUMXW7DzwMPYqKR
zrbtG4mj0pF81h+lbg6hj50pfoF/DM2C0MiKFt1ZtJ/k8Gepm8wH/gmAFk7JNmYPu4IFiv9DEx+s
1aPKScffQ2kUgdrnfgYhpTknAdyS7kzNSArKWmMOaxtvrE6m9vqffGN9Rzrz1M/WhvLn7VS9Sk1h
V0Lq+X2Cs/ZAtaEr4zsByocmg4BXdye81HzmiE4NJzjRQef2hSNqb7mnq+d4ARw4wS4BORObKGHD
1LbBpFbxq1pn96hPueR0MLE6WVE7aRz6keh3p6MwYRoPuSPP6tGmxvX7ru/ZmG3TctfR1CM97wFP
LMeE/H/HxZLXTyE8U9CACaCHhhrdXcoKQCz852X6Wl2yLlvwYrKR5Sdoql0OqfODptNj2S+6jdqu
ALF39h7T/VLkyEBk0PMWqzOAIWfhopezCedqQwbS+EQzSlUgQrAQyNhj8VPPT+jeXEi0y+ZdS8gq
r3fbHvS1KSZmjCXtFgrZGR1kHKgSxA6uTN5nmnOnpfEEpPaUa/n/My0069WiGvWbcWTdvVuyq1ic
m5/OkA1B1ML2mX/vr7w2Sw+FCTGQmTy1+2OQcI3ozoRgmCEJy4rIeaCKk+AEK+x4oT9pPE3BY3sk
PEigbUCKgSlgCJFmgIZK42v1kz33mcGDsybFV6wsGgTYKAohZd/qdaBpDVTaCQbv6V5+ykSjZd/p
KK1YgwuKyTAl8Xv+AWCAOndNk6u1GapYNJe5gdBF4whm5UmH+hHw7+dsbcOLDicm/oKO/T9eUs59
QtoEWKJ7tJo3+8OPCGfyHB12TZ6LVsa9jnm5qo4XHydeMMbHZw1LG2MToEkgable7kgCPlm+gK8u
ecZLSSpxe4EIfppIFwVW/dOsjudl+Mupke1mETTGq84dSBcxWXDwx5U7ZiuKocF9cObiwOq/U0vN
0VXYqggGOFW6LN0ZgEeX7nR669xIBPzC6+1lqcwg6QSK4Zmiaf8IGJ/GFqiBhidC7+h6N6SQbgnO
lHNXuc48V3CbMFkZ1Y9jE3hPISKIiOsa+SA/CcC3lCCgkZkMCQPIm6dZPF2ysoXZHKMlBGy3O4Ev
GQF80JEAcIm4nvLG9289+z18C6IcMqBv9JYjAVbsOrGkMCc2lTwebSN7Gkuloads4MymS0c+b/+8
4GpNR/ncv994o6P+6lG+g7oYh3uS13EEegyKtiO18ZvvlQdOLui2DQBUi+2iZSZ/Tj6gb1mGUbR2
mECiuwNL/dZ8huVLe7AcG9aZeMHisz9MHr1BN2t3kvRbT7ouJDpdukNp+4WuzLSTa+LFjXl0fopz
HxRgbcCC66a3bELLxeRj6xaiMlmKADQkfMLxPcU0zHwzHfRG2/iJC+1jweAz6MIf0icL3AnZlXqW
u1Btd74i6o2OPnPei2AbbLGGCt0rq1SbkB3Hus0jKID1fY62Y9W+ny0ZyG5ZntXTis1gee2zHHGE
sk7QTxzAtRl7HChCu2euBsy+kfyg/XnWxto/hFtPg1/VzKJHLDWwJ7gSsYAIbrbUNIQcuRpEhhb0
OBnm8ccB8YUjqnOGS39HbLRud8aOtpPRv/j3kqHqR+Pj5isESI6FcQJPmMHGlpJHxD5l3VoVHbze
/BNfIng9J0KVogPd7QTdDomm7mf9CWX8YsPi12pfEir3UXFjUQ4NBtkaQTS7lHVFZV2mSVrGRYbP
/oEdBpiPu20NGCn+tGRq0BfZ3gUs63OJSXLjHBLNbhZFz2jqIx55EBGj53sMlS3GQV2Hcy13+X3j
GIh1zNyvoQLY+GdtDFPvWqlSqLGlqS92WQ9k21wOnyVsXDeQPoFSGbVMOsFiPU0QhjFx4Nd8+QLs
OnkDaZWXJCcfPmUtmWCzyDeT34dkPp3vvW+CYF3LzdPGtFc525pb5u7Zl1NymOcQ01j/Y19iEhGN
os3Tq1ZKdjO/2YdjEO13NN2UFkU/+EGm4dqAv3bM4AAGbudKh+fsGnGnlnHiOJnIntwmru2x4SJh
+WDPb5wDK0bk6zX3JtujPWACOHBcqpbFTSp0HCJNdXJMr628BDGN7dZdC8or/r74fT+LhP/iXmco
nzx6yV0Yexvo/O/6O2hQX87hIvi8buPwwNqqompFn9oIdEBWRIVZa3rqpOvkR4n79bu3mv3zttPX
xBw4QBHPBvOx/AWEU255KMEhQgbf9DoDicbfsCZUM7NK666gfywuQvpsCH3nXMgHUblbq6XEKYa9
PpRIBK/ieLeI2utlTr2Wqe5PluK4rDXnomXXoxWidGUtyfuOoMieLaCacAMeuA1H0PET4j5ohDeU
l738DxHqp6J7FMdabrIdSHqiZLnwB3yjSf0TRa0bMsIn5iJElHoPeVDI2fsn62be6VtWrynQkTx0
ktAC0Z1/LcHstZJGFtPEZfoi63A4zLMbVk+qCEPrlpbKYEguNl7BB9Gln+ZLluzyO3NFescDFfIZ
zp/WMTeKpoTO4LeQL3du7rl14vE4nJZQg6KsPvM0rjtxAiFVRfpt/ChcTXezzcTVhp401r5flqnJ
UZzDO7UAH2FSVu/P8LTC1FxyOUH0g/ZuqyKnwL9IkzLVqVHlNUWQHLS+Hdy98w5Cny7asiWA5sIc
zIu++0ipLQZzqD+ALSpyM49p/Uy95MyUmmT79UFJWirNQUYMTxcxy+0hojlKgk4UMFxwcxldyNy/
bLDgiuPPRfMUjIWBPFewUIq5JMwPWPq7JJI6jmEgkubgq/CEPWyoeBmDr1dN4kj19PU4Yv6ncYvO
S1G9/lJG2wz5YIIy81KvZf7Sv/2tzxZ9RZlFLapn3FAjZNw4s7XFNdie4MBU17cznS6xkbI+N7V+
zVsZIuf9EbUoiiHq6MRZGaQyRIZ870IBbpw1zdMKcuO4aRu3X62Y/LY5kYWzdkr8cDwPmle+9hzI
jxS5122M1qQh8LKniuGuV167DCJ+cZkyAZmdviskM2smOBGbOpRsSXWFfU9oK4pwHzAb5lAD2ZB9
X1hUwK+VwbO5RPZZT637cnUPa0LPMfOTP4QAAgceT0RLgN+ESos/9yyLrDXbWjbTp3jryTKc/xCo
qhYuHzTKMZzq2UvTAX8sqPTfv+obSq+Tjo30Wonqvv/dmI9IpDdGp1xwcboN0pq6iTJXEAEvEKpJ
PJ88S0L2J7s2ahaKSFbHACISRqeyWCfTdUiCGijKO2FU/BtJcGmN0nEMEWVs1tAWkL4x2T1YYflY
dxFtwRA8VdFDjAeA/9ta7M3KhM/o4gUz/6ZsAIYrvY0tSwqt9pssm3V1lMC4wHMkCV4LGLk0cydm
Pens8DHSBFlz301RjJ//vd7h0u8FuOQOUjCHfCtbuJXpuBthSGhbnKGs/RF+JG9hVX/4r9/fD4TJ
VLhEfJlKU/ZgdmkHkd8WDzGplFBU4zLa5UbaA0+ApV3c6fX5eqv3jiGwcAxmcX/EA1OR4FvJCaJI
sGlh2NKqtd6fCvmq17D3ec6lwhypkXNk7bGwxl6w0nERuWkvH8sVjCb7jYFeLOgrGhRqUc68jV/4
P6n/WBxoj1i0yjpm6OloO5S6JF20mHVvc9Zt1CMuBI60VM0Nk3ejfaMkjZTuRi3yzxGA6hPl6lI3
IPgla4rzj5/myUilOTRTl76UzdYLJrcGTQHRcP+jp+7uPfIqt3kbXRiky73u2PGEESfnpu/L23TP
XUbibWdTw18V6AwsWdezsyiChz+aMeWP9VxpGc8A+o5/tcdB9L9AdGddLTHKaxMhlrUwnOkHY+IM
tUt6VxSxCxO8mqMlxEOs36MNOWoIDoo99hPTjcVCKXQEspJQOIiF4xD0WWWvwda/WgiUEi1Xg9NQ
7jna9hkyv6ve/4laL08GarK/y10fOLalgGwWvs/1kaB6FQKebBdFEsvQzC7VvHAvgcxgYoAHfvhO
a0OeKvK2XKYf5Jjo91T6a4bNOgo5bR/K1jkVxKn0Q8aebx5T6OkOYElmGenL7MFSzBeVz+fp0Fm2
vQkwkRHfOdYevBs3yxDKe6Z2l67Qucc72d3PkHNEGGWrid8R/AxPY8mXkvkw+CvFdLXHXKGxRQW5
isz7cXPk/Wwj0aay3dyvz92KyzNF8NCseqD0zQBLvUOr8HmHJaUcajIBHel646aLr1Iq/2GtzxT9
4ViOgQt7QEy4ZHyLq7AAfsFfBIZUWLpruGsbkVeMp+92JFvj2CoRxT64ly1Ml9ayUd6J2PeT+M1O
WitwpVSu8bz2J/5oIluwq1PjGN/SiE3qfEWm4wuRIgQmh1WMBCrhGJf2rNi0wWeScFOm+joeJfzh
imsSf4qCMIPx6HrRQuGYa7kjA5b5p1ZNwbLfM5UvBtYqEEOAK/M1HGpIP8TU6Nee+U8n+uU0O0PV
F2yFhdFjxw1zC2R5jgClitypRu64bNzvkcURi1ziV4MfegXO9Qy7KHRrbEAAc/WTGOgB9MZbql1J
zdq/Mfhrj7WMe5v4hNg9IU9XtkwQJATmzfQXg522NBf/AprTTCo9Huy77TYlzIWw0hpwAQ6Z/cdY
2kC4ZLod2gurrbYMRZY6bSq5i4hrERGp/FL4/4tuAqGYxDr1aPSd/Pq2ZyuneM94USYLuLw6RcY0
ZXtc13qT4N7W9o6/brteK9eKHyyyB7p+/p6AvIu6J8x4JQLv2fPwu3xk9C9mF0+kWvSw0XDPriFm
sc70KkMYCXIpS3PWIv9OLMgeu72xVLL7VTR+P0sB7OJeFngpZIYjfIIrSksh4zNZYs8lsa8RhcV9
t+kjT04IugIdJ+4bwh6iSOCgLA2NOnioC2ISnX6bGPdk26Em7H7ksvLoLWOcvWdXWsxtEJUfw3jc
mHB7TqofWiSMYODegLvfct+2uCrneXtuFNhirbZY7XdE0PHYdHRzSYS5nD4GnPao9AUIqErf4Tuq
wkXyw91vc8FdlgACxtVXDRRdJHCl1TVBzZb9rQ+acQVCsJGthpA2KDookRxSTcRGElBA/UfZ6DTr
vOLvf3CQB3povb1a9UOOM+Dskvd6FulNlpUdZMVXayMDO8zIinvnKrtNL3gtiLRj+sOKN+FDR0Zy
onluAzOou0jPgNh1UphMLW1oK9vVxeIys2eYy+FDXKnMCHcDcxo0eCGaKnsiJvn0WmWuOWMfXxgk
cjtNm41aq5s4EBupwqVzKkRKzCfue+qrt/b/iM+/E2XtKJZli/dNHzYna9sCndXbQIJwPPIkPdfY
o7KP47Ykl5gyFslDeAtzIV/YHcoR7aaORmXpLxhWopaw4xL9PcsG1rhoj53tXp5ziKXug17N6yMf
BdljskUKLDbXHN8Wzb5RDlcZgaC/v6oHKmqMPeuKShHDAz7LKeVfdfv384PQx8zo6FNYdLGwZ7rj
LyynNZhln9RkPSCSh9YpXrNBX1XGB+xjE83TiIaXKSXwVI9hh7N8tX6gslk2xqrFFwHXg2IVUftX
d7ZgCWvSMeeNy+JY3gyTJRt6UVegT3DM8vBsHjFp9PpVtiaAeGRuLyfBN3EEGs2vlyC8an9AvUUD
TFfFMsP84S6QSkJmc0qlM4E+0735iRAfnPx83waLpOHR8XeuJC98h+0fl0xDCag7WVdXqjU5Rzrl
9X/pqHcusDxxfkBISOKl8i+NnycTY1eFL0egKGYGB58n1TfFdsMGsA7p6RmkB0JI4h/fg4JEGI5P
aarntLi3MTi81Y0Ug5V/uOm9A/l+xio3wdfxLTOQ7zKOgAd5mytNM35e4Wp6bqwg+mh3b93dsko/
ulKROAcmbiar5Yr0cnKNKDQEJXvgt+jPTS0j9GjvrmLaptggZkNFD50eIvzpeyK0QDNVnHQToJ7I
itV605u6dSDplA5XrQ287YWk7gM0YeOglfJBt7H5IqzEyYpXpAbcI9IouTDWpAxJEexcOUTqAj1h
zu4ExnWa313k7+vrxPN6/5vpPxk8FVJFHXa1lgaCg6LbkpR0gTGKnYszQLz3sq/4aFxoXL8vy+Ef
Q6OIaThTORraqh8CK/3f4xQiR3+ljZ6z7U/XAtBzs7brjf1XxJvXo0oKkk7cDJICH1wp89SdBQbr
6pR/tmdXDUBCk+e6aYZCEBZOamsUsNQZwa96JsOtyfRwoaCmNkR/T/Nb2uFU0Ce/FCymBbkM/4gO
6mhtdi0XIDreREhrpZrF1Ib+Yd20vX3kIq5zvAD729rHxumHiyvFr/GxHghlHFKiJ6VWjsKPGM8M
sU6Ho37HRpSi/0Zj592sWPGhmpYBt5s8EePiw8ZQIqhUGOmRXkbBGyWdh6pLoV6C3tNt6diTe38Q
Hu3BCyvaF93Apk3ThijdGCoy9Pw1oKIJxYzHyMXu3P57sXm7sTsbpTvNcec+kJ33BAhqX3usTAhS
NK4ovQY5S2qECJ3G5UW79luTA0EE8WSki7u6BGJVp2c7Dm7E47jQT/itwBb6as3L94c1XMDB/Qbx
wDIrot7dpNOLiMjOAEkRpnmuk1W3pftIQDVVvpLo3skzZEnCrXnXJZv1VbrLFSKCx19oSKBAZYwQ
i7TAxc431df6Oixl7N0LUSHxGu821k9IP803M0ypZ25IoTIFlCTpT3+1q2ux2WPeNBj8tbyvHnev
nQYMuWVc2nvylnJIwzaHWsDcvHidgd2G44KdUg628/IUhK31Mn0ILEVbsm8CyDCrtcEkOi0+NHGW
g/071pnMIfXqB6zfKRbjKmDWH9WDBLdIy+fifAXLrcVUHWRuek9QfT5zmhgSQfLismKlqUO9a5NS
bqupCYnHoQl5DVIblBw9jbuos5NFgC5t2zUMYK/rcTu+117WWHUi2/ai+Z0LMPazBpOfJb26wpzn
AkPY7DGukg5TQtRLgfVpMClEVe4m3+k1K/poDMN0DOouF/sfR+9+R0x/9Pw30dqeEi3bm5nh47Ax
8vbOnLtJHk8wGTl2VBuV1vXfH4LAHEfoO6KTTu730LXFhQhZEviBCJ65obseyFxUZNJzKii26Ipf
PRoSZeImKQWHWQehvzm88WMXxXyvJ/elWPvINsuTeecPqYfwvj6ZLvLEkLJGRm/09O0tT3MOugMn
w5MuCEQhZaCVEpJSigi5R6dFfWNCGO/inDAUHnpeQRl9+rvWUhglYUN8P6EU1F8HHYKFz/+a4B/a
5MaOyCISgmFghLY0oJgA21ZjJoZ3Ks81oOdN5+ji/TllEJwofZMTwNVzZgHP9iGqgl2Scr5fJszj
KjPPCXgLrqMmbF8FJsiq1/wGxTjixeCJd8unxPvSVYZUif19cuAyFxtE8kdoj04MfvuX+UFaS8O8
N87GqKvwwq5mPT6AyE5awk8V7uMdRbYwvmqBH2LvVnZyzcOaHKYpaCGLs+1CAmuOFCE2WRJR5NsF
vUfQ+DyjSRL5AHRkvnfSXR3gqSitB+5pSr0fZeh7Nm7uqflFpiWLPmdzAk/InnYh7Q7ppCHLniki
95MY7Sj2blV+ZvvgJXNWwA2JPE0cv860FpsMgbYjlxvnublhHvdwkJ/Q3upL8fV1bsXlOJW7v8P0
vChvibE7aAnaUtgm6RQqbSxXdAmIJLU+PPjeVwfnYccO6iDKWGXNHTIvCfRDp36qTUk//NjuKH5t
uPStiHxbfn02oZIFiCg/RAb4FJt1tEQvmkADyuNXPIrfCOxFLT6afXBaZRWBfgxhJN9fWyd6mOFq
48zugmfeXr8RVZQMemE4/L8U1pfbSkDhZXZT8ceP6gW6Mzj1zz4yaxY2ZdZ1cnnn66ubt+H0fLcP
UpoTbmhJCw2G+4vLIfk2TY9YxYqnZ+GpZp6gDMN2eEOQZsbUIIFIaGOD+cIKVWWexLWZBUH/c+tL
GQLa2HGXpg0aF0n7r9i47RrxVE56c/+LMII+Cf2c6rr2qn+be8Uch2jCYgilvrxs4+kx+Em3f9mV
ecb2PuLxNQRaNO0Co+HwDWvJ+oSAoiQ9uIBI6BjN6QzwW+RT74myxLTErv/2Tkbg7+KsfzBSr70v
usYO3w+QQ2GuIR7Pk/w4NoX4wv4UrtKVsAB8+kzwdRwzBD78XSLwoTyDL1nx7Ye0vnR1ZVmnkNAn
+3XZA028MKioTupxHPSshvXialqVL+yvsLCc+L+ua/V5z0EhwJDHBJfdCVPXnhGBbH1h+9woCQMD
LIkJr1VEIYpVuoDF/x3odi+vYYh9/KZNYQvX5Uut5Kgcez+juRTXY/6BsZvVrvs3VbgBEu0SBRCq
F6UwIbnn7O8WkzWLP+gYChsI8c2cvHVo5xDhKXhx2tCMND2j2Mv0Y1PwQDSKpcxYf2EEeGMBMei4
SQ8erJ3/ZARO2C5qHi0MuROohaQqbbYQTkjkxZed09h3WwB4BrwZ+CdPt1UEQLFFNla7+XMM9c3/
QwwcYF/e21sfSBD84hzrRZil+ptjf8qru1aQAkeQQVB4xaFMbLN0SYmQ3Fz4Khxoop1PRLUnCSQB
/FEvZO53mVXNisOv3Xz6vM56m4o1+mqfkIZYIGsNbgEbqbQk+kd80OeJ3XEPT6ofe54AndU9UM82
B13IZkRso/JFgggUEMiMGw7KUb8KH31STpqbOL584Z5gn5ZpScJhYIWskFWIsjg6S8JYmelYNKHu
WQv57+atwfJbpH2CKIyO2c4njvRlhauIWUyTqA/6Z62ou0up+WnMRBy+cwuEHdjgTXoQNP0LXz2b
n1nCa9R0qynLkM/I4KJDpQ1Y+L0AQS55IfGDwJ51HQoqU9guS7YoMJU717KHJNXvBV5Y2KktPOVP
HAkdbmeJUK6VVEjhHdvZRUNsV4aIMCpa16ycwjm98IEbmwLaltjVIamtI1KZf/pr5agccyD1Au/+
HBUxivNfI/ymSZW4/AUpLDovDGRfY0rUN3hQIX70uRZn5ERJOs7lQ2uImp8wVUzdpgaBpeKcx7DX
1Vy+PJ5H8Beq04kNqCZ3eoo/SEVOllNyCLMgR5nmJDWU0TIFh8jS2M4w+C/Z8fpsEI//WjWJ97lr
s0FDFuoPc8EUjfwmOXvPN3cR9uAh7qcDO1Gum1HrYmEMSsJplryoyKKA3AQbqVozigLpXN2AqikD
l0WjDLCZuD4GTcv063vFrFtlVZ8RFajduVS0wEuMT1+ze3q8RM8M8s+HRBdoxQcE7pB91v3RPxPj
uz3upHLDoQr8kTYyQQrNt/LWfCEpqHNcr2zJX6OC+tx13QuOhG24h4LwHE61fx0VSGQ0w65jhRCE
5bXliorLxJOnaGNKO4ZfCKGBLgsXe0+sIOPx4q25bEUDHCzKjbQmcoKhiAqCDHmFBTzcvcZED26m
C+OBHtrtIv90XIiW7btyGzPYDRoY+CFPEAi7At686ozv9zi31LZGF+fO5dNGbLbZTH62alN2ypJS
++2ZXQzR8/UqMj7t6DzIkHeTNX6g4R2kNOrFXq4UPJmCJShmdyEFqWRXlVnvjIc/YjP5aXfrQWGR
rtNCF4MrLCyMy9Z9/PLuS+mVazsGVnFIyAVlEd4TlPu/X/GIjJngiOBiSJLyDCE6rC9Yi86x02kx
I7M1Y8Efpj5H77Fvw/U4X3Km0M47R+0jOpKgFUT+8tmtYY4t2xD4nk7n43ZMpl49ykxfgVs3R3Pq
OkfiVvzl5MtjWEiw3JtcOrJk3kWHitPCRyTQNyMqZDo6vcysUT0WJp6ONRFtlC/pfo8u2EK0ceO6
bAleLimP9BZGkvkm4SzChCIBl98HmBqbllpPVvue0x2LimiIZkovZM7RIpUaNnFQT+DdE0kpJd2G
4W4Y89uYYAaHX7EvBwbewblV7ci2ZF5Cjm4k39PLe6yFqx3mPdQT9UNWJUOEmfYrxjWM8Zi2DrfS
PP9YnzF55mcYa1qUvodIGq4C0O2Yn6f7nS6sqzqs/8+NQynvRJXsv/J26o9nZXc+GdZvtSY2/9/h
Tt+XpwtM9orzo7lF9sNMrwlVROomYR5yBW4ifRKCwK8icSe7fCiQLDymQkiWfOotiK06F4elf3Ke
ZXZN/Xw+/i6DOs6mBuKDPmc73ljS9VY0zQkHiFrFDo2lzB+znVtqL6+g82FKMW4QwoF8+8YcJW86
p8zlUxl8bHFEyOQEBMgsVxwMjfeWWjEfC0zcT66XedTsDQEg2wbFm8y4Jt6DFb68Ed54GxIFt1a6
3eUBvOd0OPWfTTQvV7M+NUdvlCw2alIK6YNqDnH7FGGbRtlPJoDoip/+a80KBXzMJobxupQReTrt
U7MLeDK+vwfXLO58Uo9lAYMMKh6kljPDsdyexS8Jm/KGWMU28DxZhgNSHzjbgfWocD6JoEgKVg0D
oDFk9crb41qyxsOpHTO0WYRPGhVB3EVzgHL0lL5pGlWVfQr0J0e2jMSX92fugJobevh8Se9NGZZp
gVoZaUGIVnJvLmG/UVRgeUVWOt6vq2FFhXq7nQwKzXE7LaEv3AXV3necEcohJCgtcAtoOymL+MVv
+IC6WKv1PHY3Bv+Lp1uwFPdUWtzwxYjqHQkR9SjOtBQX7x1eF6zL0/hAFTR6Y1hET9pEf3lKFaKO
SrxUgdP9nVZBoyE2qm7WGTq51Trjej6pehhNE0jPNc181HMqvr/JHagrGJBB2QTcjEXb6aI6jOQb
HjxXO27m6XWFTd1nvKSpEy8EcOf3tXRukxZ6hr+KGyWjj0aB0hFvOeLlU3CVboNOE3mfb9uhBa8d
yVfsYX+oe6tPqQE1y2KmHDTSEvwUrAgaOJi7LDgg4vRlRfG5c98xAlTEg+FxnnUEhDCaj5UTL+DR
B7bR1CXMCCo4orRx7OyZkQs4yL0e71VQYfEF1MCuEcFqxCuJ+TmYm47sHFQRU3MVmipcCz1lYNQA
2XEyftg2+ieo3A0Z6xR4MvL+XOJidh/kttPbwgfyVskbN2E2vHTzFV3FCV+jDGYm5DgJwgPzyjkz
QyhhdyU6jLsbtwX6Oo36ft5thwwqMqCzZc0pXAj1ORia7wJc69FfudTfcYlPe91A2n5DyyI3MN+O
kcoWhZ/sGFmxls7n5hfhXHFtBazE5X2LLSNDXuWu72o0mmuMMUizz5lQqxFCbUPb7Sx9uo4IaNiI
Bix4otvk//me4RKSS80sbHiOTxONRoapBMn4OEPqCO6Krs6pMT/nE6XqU8C7yf68CsYL+iQg06U2
elr4zTqn13pSggQxWzx/gWIMLgNznmNEfHqctzaWaGiVg8xpSyrtr99s98JP3Cu8ZTrAPMotCQnT
Xl2bK8R30AxxYtT7KnoB2mAeGfGlDhM6ifDH00PFf/rbwGmCKuiOX5SLb34HO3qn4LELNA9GF+74
Mjs5FyYqsvtLbyji55CsKcWHQejhL2jTxJ8QQFPX60s/XPbRINKtd6U92Gms+oH++ok3xZUsIcQO
Pa9KAcIxQR+B6IIXBOKGfzZk2uKFF4DtylFzHuxgMM+ZozdgL0ANpQ6qR+waobzqNUV0q5H8ZtmW
Dz9zvQw7v+hB8Nfl4L+RxUZOAnVfk5uIAeQiCC2Z+dGjzepa+/dlrTRNnClGldwpCPZ4FhLsz0dZ
QCWdsHktcTX3R8C+kj4mrUQvYAlR+Bd/n3bH+SujHEy4teB/mOYEfUh8Jgtlmt4eaThOKua2wpRp
PJVh08v+wWOL++qqbjL8/G1+D3DEWW4tF1xn0ivS9m1OT15f0pE6qLExxYyhgq+mPCazZA642wEP
Jw9V99rUORueV994/bB0/nnUOkgxiUdQrkQyRxz1a0ufa/0uYlLXLIem3xhTqk55ynKcJ2z7bJcZ
evsKVovLR7Bgx5bTFv94TRwmrLJbNhNp7TcffFlU2U5QXDJdzVvVk525HUM12YOa1pOrIN9Mr3XS
yWpFgtDKlA7KS0G/Rxtq43j3nYvOzfIjdkGcemDGf82LUIlxRiCJOsNuQeYDeiOWB4tjnj7CiiiE
lYVR9pjuhNtKYgvx/awrkruo/AYm8Sa2QUt4EQqntCfkbpRMrSVuuFxwS6HGaAf6d3qKWphkk5XR
aiqRPX62GDXROgLf30zol4hujNtlLJbrRBpG6feIJWgfwcMuoLZzZVzbdaCRLPimY9aWoEf5ZzCE
swq5dMmdx60azFwm5uGOTQkrGguLNj3AqSadiPKBe1rPE/59leuudO9HI47cQOa4iEUCUQoZTtJw
vAV1rTyvdTfbMmZPAI2la+9n4JyWWzxyKOidA2EE2Aa8d8L5AWH7R7qmFjVDqtPQDDmGtZzDbe7m
DySddUZ4e9DMu6F1LjPOkmjcBmLawwGWvVZr7t7pk3BCjIGMofcKnHnj+s+dZA2nvBDd6MqA4dCa
6f3wnniQ+5KQOy8eM3YLhQpHjvmnSNwpkALgzXVwIPhqagLB3/rrJkOTEFSactSUZnmQ8m16xYrv
w8uDSTGLi5ShMsTviNbuiuFdF/vDcM2TALYG4QGcPK9IOX1N8njFeOpeQ/4BqU6GJTDOXHL4PfV1
eIkxPxrm1XCT/v5KkjsbiauohaEe0vK9DT/RHsRiPBi+XW+nGeqAGbhwUrTTUbIAttY24i1sFlYs
Gah0OYxL76n/f1bDy0Q7YFjIfxNuKY06kr23BZ7PGdRuhrD79YDh4p9mY5NboKFlG3pSidB4Ouhx
p/gcF1httMftRqC4vNggWKKewGRuC1uuH/zW1IjtEZxpdIdhgqzUOvb2jG3A9MUSB9pZbWIh9uZW
2UXDYJiBZl75XYjqpMUZ62jAZ4U0PcWVrAaABHo1qsDYxoEIAockVNFChk6elniM3XzEVXKOMj/R
g1Z9klaUSW2ikTFwTWAeCyT4xSTJXumpI2IyKo0Jx/Usczsy0/E3OsXpirWNuXX7cEwdsgOTx+q0
iPDV4PTZhNIfZly5FOKzqIGDFX0DTLa1M783opR3fJzV4+VjTaPuqK+BH4fyuQVOwy5GrX/pfQh0
WSUxDlCw/4DHUgGiVqOHrxCxAuF6AbMt7hxnd9ENURFykA802I9KgFb3+UbSlnpHiNHNjpM7DuqX
lQgStwjTvK7M8sYCQEy+/pGVyajiPFN7NyfKpPZA7y3eggKO+yMLX3cevxkm7/dyrKZeu7oo+Pge
Yzhy32iGL80YwppFhT2b9saSALR+X9qrukEkd2/wkr0ikO/g0VNvgTKZtGiiukf/ecmHCIk3LjO8
Q+0gKK/vmsw2DmFnelQQtwa+1UJ8VqWCE+eYF9ycVotUkzHSY7DjQOT5wZo8Zq9b/JUdo8A9nVR7
FkNqXWP5uYbP0lIH3To/3RhyNQoi66/3wzherF4+TZVM5D7oK7p2VsMxxgLW62QLm6Z/FEOsa69Y
zXLtL4uNnfoMShxm0gMhuGjgw+0uZ210A2AiUF9joMoDhn+3VTXbIanSM3RLMY/K6CTodK/NNMGR
zjQ07n7bAh4/4UAduNwNinWjXg2jImReUPMW5podZS76IsyaNfk48fZ6kkQ8Xs7shraLPRtB+RrM
NsiPg7g23q781YwALiCWehA9ZU0xui/eKYk7Jokk6ikZ/OtmuiRY5n7Tgp59yrc19GfM+YSMriY3
F/OlRXxND62lr6GsoIOtL4ax5dw8A6uBiXcYWV9H3rrKwYMH5GGKpVgcNZXqZ1eJuOWNGCv77Tty
16r6NGY+qYf8OjZVpU/sJZgnl6QfPoPQg7gaX/zWfNtWNkvaUfWij3jkXtoli5LIlr+/ZRk5vY4q
27xTlQtx511BJiBSaImIzRvcEQU5gHFaygqtDSczsuXgeGIFCZ5ozeTsvl7nHlUHhEIGVp12C+Id
9jMzZKB9TkHOMRBs+ktvOC0Vj9QrJ55KlC9zVKI6HMHGMUQ51RGnax4cyBulxQOM9uML3u19bura
wk9cxZSJF322jNd8pJm0a+sPXKXNXVCZG10EB6+JOEB44gLJBz4R7PIvO592lQFd9mFdS0W7DKoJ
Dne1tmdf3OrbMgJVtiMyqNKg6BsiYYKxqZtzc5UVFSpTFPJd5xnBjZl+I/FO4i55t4Y0LTCjfgOl
a2+VQIRpI4cabFmRujtlZwL5ANAP72pFshdP3ddrmgNCy0cA3OM49AcTlTM0EW5gVXgbE5UK2gxR
Ei//ktagtXDDCaxOOfodqbnOQhLic1EN/gUhxgsaRmHBAJ3kehk+w4ZdyPB48nZSYuG8nWHJR68g
Ty4XU/iiHjKKDLN5X8aR+0IgZGn5dKwRCUX+piop4aIE2jEyKaBtug3/2h7ZH4VwDOsxBN6ZTSV+
WH9vlUwcvV8wkyUs1ez3fmxQMkxEO0ULa4+8ZF9cKzCw+EDSXTS0zrvf/f5attb4zEjfeK0ZWkXQ
JUFT8zniNQ/CMeBGAoVyisNZDcJ5w9UEI3rbeLnrL/YSRtCIh3l+sk5riH9jnBRAlG1VzhuSXSjE
jC1fM6b38qmnGZqho8wYCKP5BMLgrjo4l68HFxyGcd41h9mAA9iqmtNy62V9PQlNpFM2o5WCiu6M
bCg3BGpsdSo9iL4Js4HTIqG/YkPyxMrZA4h2CA6G8ihUb+3ovzHLegNCPK7Abwf74n1KBuLQY16g
oYYK18uiOOlto9Lh8O8fuQufrvGVRwLKyWJlyIBNFx8IUgUcYsiCn8k6UsLK4GQossf28KzVzrVH
JFO9BC/w/HFfESICNRXBqtmv/HoIrTBY/lYd8BbQK45LD0TBTLH5rVDRXFtvmrfsmVnKT8taGIHA
qHd5zVICi3foqXnYfJuw9oIcDoy3x0MOnb+vj4HBONdkb16jzf9xFEnWaY8boptEFcJt0aBkAVm0
KSrXORTt4Ssoc1/yV7gkpzMi2AK3VKtcZP265zeiqAuVjPztBhlrgrGwJ4KX3xbHCmP0cDlZSFUs
2k4RxoBpuG0sv86vmgH1CT2IYtR+xLhDyNGeIcoccNmcINgLO9IclbgWr8tbQkg/o4m1CBhfdItK
uPzLdzD/VzJU10ghbZplTkOxd5pZWgwES+4+rLnX7xLKFuM+w/tYyHEBncxMprHjMs4/3XrWvAPH
sZGPyidEoWDeTLSJ82fO3Kdbe3fHmnKB3wwim1Q02NhyEWnDBDjDl9MtppSRO+gKZV76X+P9ncoB
Ck26BP3xHyzPtMrS2bvxeFsQAfdb9kmto8Pz3rFuzWpsOgTkD5+IpvNO4tIzbRDxSn483Kfw6S9L
r7J/jgXrMVQDDZRHnzkuroon0riYW9w5bJ4NCkJiFNUY0nrVlelRnpOBXD1VXlALFSKF1ylLqM9k
LmVUWI57FlPejNv1ItrM3udQr531BO3tbfv9C+XGSSCU6/tkmdw8Y+XbJv3ikfLm4nQDLTwKSje1
CFmQpQjWtWhkkA7b5KcUlhlagJ/2tkT8iezRLomzxWGuQdSZ3gQyPuDQUHUUm0hOj2djMnGRt3/B
ouiPrsvZhv9y79LXyskzghmc/buvulxJZOxrgS6AZppwbvumiqYWUip5foaK+MSkDCYsCxKnJBAo
BEh220QQ0kC4MrW6i4uvnGauUIcej9tQTJKGz3A2AgQv2qZDJtU9SjbAruym7r1NsIhMA/0P3qQJ
5k8NXfavoruTHQfp8RqCTAVGlhfDLAkQPolzsDWaJ6Sy0WiBY/yJVL8f1lzoU9SUfa/iiJB9F8cz
P9QV4gXiG3oTr2pBhe5E14Z8mCIFUYZqBTiKfYJZb7Y23xk1KlFtm40+gJ0qQlS1RnTm0G7wtOwh
7pRCLf4DsjbkG5dlTXbZyzIRBIh0LIvRAfGVLaZB2DfhmHpudJ/9B+L1EEiHQNtNGjAzfxrSxpL6
exJx2wglFegt5q8Nx+ru5c2abB28gD9J4FyYkI2dtJMesxwEYR+eRlQAGspEpbFY+hXgXttvPhQ2
MhUerCMlgf1LvNY5NYGYs/ZghY7t88Ne8kNw2zvlhOm51TO3SS7j8wVk1i6Ar+7vACCxOlOlHUey
o2NMYkrZuBsHg5v9+yFf8WEIFuoKZV+PjSra5h4hRtffCLpKE2x4BSMXkA4yCGOZP43+FsqQzTnU
e0Cb3xRDD5wkp504oYfUuD9hkNH/VxXWCIcbJ2a0U8iKVf/OXO4OI/2QkGt0zIlM6MwJZ+Zgi5n+
fcfUDavtJPj7IHbBDtwK6j1OHS5V9ELtHafic6LhlNbV/U0SUoFkqq3b/Nlr+hm/6mR/cook2Yah
2JGcR9TpAc31efRHqyBxuqjMUrKXd7bg42he6xGgA2O1KxmCox2/+8mgKW3gKdgVOAK+RB5rZ+a7
fX3z9AMpy+61DOE+xmSz+c7KCN+aQCDYMEviSJqqTsOw/6ZVPA0IMuAFVzrwteM2T9Hxe8GU3fib
QMCAam8Tuu/ZBK4AYmdNgXDpuCZcQuZNsQrpdfVGxcv/7I0rw+AbtWombVjejz3i1QbZqueGFZHr
l1por02i3mfz9b/8q4P9FGDrkxZlyvFJ1GJNx4w1Hi8TMAT7jYWGB+O1TsIuqpx1ZfeBRGda8IDr
33uW0IF1li5DPam+5wCtJumwOqb6g2BcSjToZ3dGtraOUrpvrsGzzh2v6bAR9jOU95UbvIJY8sas
InTDihbdyEnHfqsqCaP9Xl/yli6z0S32RpjIzCywDmVqXtpxusEcDSoKYFti1Digk6lb9exdmYnG
1RRz7NYPwqI6BrCrncRKB7BpvQ3O42DKieaA+wvWQm+QyTnIm8amq7iWqFoTAL6/LARtY5MXbHWs
L5Teuc9gWTzZ1OPaXpoN74pPdSTYj1TvvRX967BHiyOhOWgCe4AOnjZz3fkNnai3psLSl/0n+2+8
RE2cGkFdp39WBP7FDilqfWoZqFzu9BRl4f9Li1IcyZz5l3WLRXrQ95yPpUuwttH+14qqJrS8ACWC
Bae/3Xrx0lHB9moj1+Cs17K69qTcY4nnCJ4LHHsfRYRQBw8NMuaO0B1XPCBtdXFjqXQDjaZX4sms
GoI2PKDhKcGZ0Tc704722iiPG78R68yn3rAmNaYrm9Rm7D6nTW+GRV8uVK/BFj9rXSfc+2AnA3Qu
2G2pnesAXb27m6FJYDxRJyKasKoLl+HTCN+hHLi1lwn0uLdCvxy0xOO/4ssfE13tqgfCkEw14jqK
0pwAzIQZa+HMCbr6pKD8e1GjZX5zQ1TTPXth/Lm7ZwQPAgNsahOPPm48Y77QguOlHWWQl34aTY94
lg3RBGlOQu5OC4giWGl/eW3t5qRuoOWX4QR4jFzMWu2mxaiAZWXAmOU1Cn1WcYFnCQ5J/IjRwBRF
hC1fMS9NztAuv7nacdPrbQsbpG1sIv4fytsPO4UNQGTOXfR17oxPX7CSju8ab2CvCBefIFEZfnem
bDNtK5w7FpzGu87NtqmTgWIJkhrWCd9xaIaXZ/6MUqaiDSkJNBqMP7ysJf3X1YMih+zv9YiNTFq8
RgqyJ+p5D8I1OWKbjPTqmtuPHTz2n/AWfO/YuJnH2/4+FKXKsi9E++fSMKK/R208/OvwwFUOrZlV
NcPLoSEYsAVLV18hXsOUz7YWRkoiu7QtFXR5Yq9WLNstdDNJ2XnfEVsOF9Gr/H81dMiOuwMOOg0T
nQzzE9ptTw13gxs/rsXffAWkZRrMzCKXhgyPtXqHEKEyTs0BOQDjSihypJyRK1OrFYY64MMCJ9jo
k7AhOX9x0sXMu4EArIXs6lPwCyY8gHrXE2WnLoxI3lg2WfXSj2aTpuFoxdBhIVKC85Jz4hXkUHBs
2H2UpXEpYaRNS8cqVtQKqbLiReJHxNAGH3mCO+7fwQ2VRXKe1ldgacEXn0so60cKwaGrwlvW8z5X
AW3Ljj3dHd3rQ5ic8upkx8tAWhC4adRDy25P+YO6u5DMzQ7s/r8O5HC6uauPJoQH/kW9WuihoXAJ
Vmq3BtEWF4pR70mQXjmemWktxi5egupUTrcZ3vI4k5NgGXUpZ/WUfBPABI4jb9ni5MabBEzYFopI
aBOFHL4ASxRZJM4S7qhOGEVbqPiblIgSoAlABJa968OZBpIUstlA2ptaNZ++vCs1g/Jm0ToSCk96
X8OA0MlhNk/jpfwNd0Az3f/0MRqn5QWYC097d+v8O1HOW50Okf2MIpL8F+9kF+mL4O7QNhqKMs5o
YovQSkS02laCdbUgYm2TZpXBPKAJSKLNNKn2ZRiAYTxj/x2vbY6iZ9tpwRTNz/6G6WHwCd0IWUU9
xQmnX3vmoGjuUteZqo0eXSsrqAsu3zVL4X0hVSFRPvBMjKjHilBKjC0IYelb6Z3NK0/h8PhW72TM
UE1t8DZbhUN0u1a8nfZRD0QB9H9TPUwMl0DAvk4GQOmffaAub4WBbr0shCkX7u+P0tj6r7ExJvII
TIbJ0cozpm1RZJScxaOEtrTy3bOn4IZ6HDbzZxP6BmaePCLODI/LgPjl4yEe36ErH0vmziTpRjps
THc+Ql/chrdvQEx8zSWbJuqjYMEFZkWDd+s2eKfyf3dGtIjcN2dZMtl9ZS8o2yc98RcNPpHCV1fH
8gnmp2iSZz1LJ4jHafUdONX5T1Sx/SJNnoOWv2G7tEnF4pAS9Kw2Qhr/Ir7EQY7qZZoZFoW3+DgX
ybbZ8TU+7+kj5zth70iIe8f73rxo0D1vZ8xjN5Cnyi6sYUopaEh3PKj/s8rcMcsrgRPtNU7GwuMm
ZOda781nZB+Kq8zNwWBvMX/EVMtTtb/TT4xR2OofY9sxYI2MXnbc5n0lmKhQtqBu/EPwCm7p157/
NXR1WWlpUK3/zzB7yzglA/4CeYkR/Hq297HvXVR1mMGl1XmlCK+eHUrx5vrvxkKwN5ZXjxUqwtrS
Cwv7MOlQwu9sBkDOWuCiv0Q5yWwREJBvSGNLqcz0UaJLGPE1r7swJLFFmA1zICTs1axVSfcIbSny
9jmhWxAzE35vh/WW+0eDDs0IvsF7NynvZ7lg8M9NAQ76UT2yfKh4qkQOGxEBMdGicG4TkurEEZtE
DAC+fCxE6fLHzHSv09CoKeQjvF6J7TzBuqyXA2UYsvdVgbrtYPLyqquuv3NGTTPfaLRfwQnslAtu
upo9kmrbRtjVD8V1NiMzj6LN0u56ZxClQo1G9wgWyKl0DTRBqa/A2dFojtWMfWvmJJL8wA6WETYz
Qw09OXhV/nxVZ2EPoUGVTIvceRrPofPiT91eQ6ikVDsiriWoImO64+GzwAQvrXmCUm8AIYQ3Eqvv
8wyIZ+ng381cjGO8kGtyRCz9f96/tuTwTo6FYm7WQ1RWByOOcrfOsF574MPQdyZclyKB10ezX2dg
Fr/er1fm6MA7mN4dn6dAt1mpDNSp3VPb9XHKn8HLgjQPoAdZ7XBq8YIFxXfsJwb/3VjSCfTQLo2X
tvnZk2Rvyg49p2WGvIqGgh3rUTfEI9N0h0djCRGNLrargOwRcnJnpU8w6bxUihKBDLoWWeAP1cGn
dlwaDZutvK25JJbEy1/Zhb2PgigoCBdclRTc3h574XEs3TV3kSDlpZ3mv/At4FmkBMgjC/Wh3au5
VjvOYZdNZjm5CjPsJDwz+DkYZBxDZdBtIeZIJshW9ymEZ2vFXA+eicw9q5JybCwH+8SndaEOBdHc
GEOXJJr/V75EJHFxIWtxfpIaxq9ntckh2KgWGkgsV+UKGLjqQ59ZGs7qmYqM0WwCesCDClL4RZSY
hj213DhVoBhs+PNO/70xTEv7j38f0At4rNKzIMV6KOyTvaMKpQI7Y8GM0i8uwVSX3DyeaqL+gf4u
wbmIdeLGAzy0vJY+2BNuOXSrZK7uapCfDoOwF7UuACsczVbmnExBpgNXgaAM+GjmYpBSJhDmdCYk
QWsESbhqkgM9oPUEF40S7JhDgkdLrVZx55kwGP85/c9JRQ6dTejSVdJzmFqQJwC9fkvFmwPidJ7Y
kizxKB+fNYeCMKulrYZZXmx8P1zQ8EZE97PJausmmJeAiRNQnEaUjmiAhO8ahio97xqJvnq/Z+Uh
FtR9scHg+MDBahr4P568npiX8qDKU/+SDtoC0plcmIQ1srzQsXvrAypduDBYZNmDkwDzTvFNOOJf
cDhTjDSrtsqOlv5KaUswupTS7/488r3inxMPuGzad/GQyBZQS0+5aiJTfbIi7bO7SWP0jnRMiyHg
DibZu5qBRQUf+2JSScnf1DEOBAgYijFx4BSj9095RXAG3W001QvyGX7RNLY34C2HvxuTI4gAlShQ
6Kcg+lY/Iu7r45ScNNGxUA2/hcJM0ssDoBK5lrKmww5UyrR1lWFWziZdPy5Q2bWa5c0C0Va8/gxa
wwkWQMi0Z6c+5Or72bUr3ptz/jJt8Y8W/uVmAagpg4a9nAnJ121MOx1/TqCnumbNORfALAize402
HQZ4/d41m3AnDRp33Oh5/jqQVEmw6vmgLDdEOcH8xbdNXlx9kfdGsu37MVeHuOm013PkNkJdHRxA
JE0uTyXVwqlBB+PPow4+g5oPfNN5vZRTsUpquCdL0yFfayaUBBP9j5XWz7jRRkHZ3ZBFWvB/pA6+
VMhHm71IMGBmPvW3UaoM92ZFedFU/8r0p+DLaF+sSt1SxOTFD/h1NQTuHlAEXy7NhbWUfOHKieg2
jHOg0qVVr5Gho6zlb300OZR7ImJpFdVvztaPzdHNIYXVDRo+UwVJDvmKKaLRZ+hvo+NjWovNIUSy
Sp/smn5Qa3aGxD405mKJhAGawaJEECvwJt3+bGdsp1zA6BCueTnZ7m3EzPT/i3cpxHB4gLAyqzte
UHYQbpLdPXdDhSuiqDV2LI96EvHRpLLFlWBs2KTWOax63aFxoTIvng8MUjPVJ5dmEJKxBjtiNnMf
YsMjTvqBhz6ggfh6EcIwfM7Vilq6npi6GpDlbvYBcjCy1gZSCI7F7tRO50nrKUkUL70/R0hTTINL
K7nBNp1nH4UAiEdmObNlueYDmZMiCuByWj+chHE0UrNTZcyqTb18x58pNMEHkE+FWPJNSur1LCzQ
g/1jbeDm8J+Ur+I2PAU7h6e48dXgtojJVFzWEVhijAwBNd3+IbBi92c5m0NmTYccw8H1GUnIgmD8
P5jJ9xIpsEcK6IPfHZBLID/+/OMwi42QD+CR6vanPx+emMcSOSUWmhF+Vfvr30alkXgy82BqEj8D
WXpddDNX3Ekq6uS/ScOrAqGzVXtJtC+Ky+GfVrPY9B4/u+mKkS6xxb9QW/JozP8evS7xuYzQ9+Pk
sOxDeEHJANVRANwNQh/0nhaybjg9lfHWvK2DHuxq+D0iF1wej0C1KqsQuoQcqfe29wBG3AZmcMud
WU3JoyL30ugbS8BZJYmqyNFGkJqMPDD+9XwrQoaerRw8x0TQuoTlALW4CMSkDhZGNZbKy+RD/lJt
Smbt4ELnpPrj13hIsg1ZHOInkCdwQmvFkh2bVzkGVfhVpKIE0ieJMqAjiYfql04dxEIID1YOcuwk
3qHJpJfx7UWD6GeA1JYYeNAyPItyQH7YU7C5HhcFibXP2IScQ6OKJ+ISVhrX0iNHoEmJnXd7TU1K
sRywknTb7+9CtIvVNdQHMZxvAnN1MmHdSLa/8R2zAiu+9KEmLJIS7NnA7S9mltjhoxMtwmxlMb+q
/8FZbAZKoIgRhSBG4HiQLoxKu4GW9klcbwwR+rKKwXMc3EhWHV28mRt9o3/GNhZfYvUX1phENKKt
gj3quyi8RXOiq06bOvUzhbQNm1QRouPgkWcfrxwM470u5xgAS73TqCyKGLhgrxigpSseN6Y8ZaaE
z/mnEKWMWLLaQ8nP/QsmsnDwD6kH3TVlBsp9yu23JlMRBxO3kMr1BWzzlmu+CC+TtHwBnxPStfO9
Tr0Wtp1v/bsmbMsBFvLaWjmQDglOPgjyKETyQCTMLMhxDCvjba5M25bDuXuUMtDidwT9LaucTk++
bWbQtJlmN+bbNWtWal2neWtFEVtyzL0oeNRBD1Gu3ykojCps/iCTuKC93nAG0hjXnDbNMynMMua8
a4MCrj3S9SMnGQhpBfl0ocbtgJh2C4jo1v7Ko1w0egpdouN9Tn11p4IjUhpOGVHnY3yjUCKD6w6e
KkjIGpOAXn2JGethWLAOfBBpqIJZAydJPVzIgOIyQHA1OScN0pCrEEP58aFNXdDTVXojuLEf+qGn
62u8fNN1/KqIocF0vnhZ8DCnsFPKtN1bSXvmw0MIbNRGpqit8reWYa82vl3Ey6nN00Uzm4ahhRC/
V8ZxmUY9xRtSU/VDrvjjjuiYZ3Fy00O2sF2tdOS3bHcw1sWAlu0XKQWcMDzcxS10+OFFLUsAooUj
R7s3k4YJwQfMwhXptjK9yMTISE1ik4cKGNLgd2DyVFIFjcREx4HkaSSu0SeQ9ACGBvHi1nnr03zr
40+tiVKUSdtgdbD9FYHr6S7LeAeF1satHIkGJbBw8Q+6qkilOg8T6r2zsN5BT6j1E0NGGZeuVSrj
vNbrQTEiYPOm0ZSlNVoSP0tVSdFuuoYCPHFLr/mHt5nsDnEaK9XO/VLrovOTBAurOFYjppjYkS4h
9tKATvAZXHU53NvfPTHBP9xq66TQW0h8ci91tgjhtY+VdQu0wUt9DTa7395nuoFxC6dNCufYl5fa
yPuGt3mwXLpxClR6Fe0B7mH+kh6aJltMRkzuHu7wNlmjeC/SQQAn/A2VgaxWKuJkKBmZXnM455PH
+1butdbtDZ23Yjps2cg/vpsWMV93e3abC29FT1XXLvgRhyGuscp/Ih9PYLkp4TWsZB4pI8b4s7Om
v3IR2CgzrsN9DKQTvxNeWYCnRJy1fiOimW4+KOV3Bhp8an8E22T0XtvP3FrRpyQuAig3Bu7QT7w/
g8lvclOWuT2C9oaoejd9WUveMBnTJBxbIOzAO7hU0/an5xIJhC4aFl+gCIK2C4R9G5jUMA5CN553
i/vRaL6lac8tWp04ExTDRdr3QiKSk/oF5ELV1qJ/Jsv54wXttr17gb+qT9geAkyNEV+BuIYz4p+U
7xijf59pzMRcAFng0HoPad4qJ30go+bscJPgOUEDcpF0Lueb6tg5GZxXogSAjn87fVOeyQnc2IBx
Jwm675lJ/PtMbv+RevDqRseOFsHnw+9dWPkCFgG/XgqDhA2cmGfAFIormgtAxNV/rgrFbEayYAkw
DKYKxglv2C5AtWxKR91tKFFTVky30H8jXtq4t0jH6lNxMpCcClEGLqFwCVQP0UuYYbGOoNFU9yfu
HOBZJcfTqd7yN7E8je8aMC0xCnWpKCIbRSCtwTgcaCjQLLkJi2yBKvUS1FKqsLk6Lb1AVZdjo1w0
AeVCCRGEE0eeJ928WhonYvH0WGuCfdjHcD+WchyMOeoVGEcLDNw2rq2KbaZASVuUxCKWCn8MLgZu
bUNEYbMQXwELrQSwycxaG7Wq9skuT/H8NJFUE2Eta3rkwSbZSbLgrAi0kJLSi4DST7SzYM26zxlP
5fhAfxmRai4beND43BUZn643/E0vh5euJeIcwsfhstA5Vu4Qv8zmVyFcNp4flBTLf5POxGnnGSW1
DlzHVwrrpB7ww8d4uhwMIQ3n9Y9oVIBA0Za3cQmQxsKda1RX+6uoSTHvjQnhYDpGlN/OfIwbs5iI
cEjmYe4zyFIlsRHGkfj7PIuMt5oLZUj7kpYcDFs2wyJ7U7EwyYJcRd/xVQlaxhdQG3V9yMhIeifH
iUoqpmP7Hc0KopbB7pJiA5Gmxge/GX0xLO/CbpyKKMlDus4ZcE+NdGln3CsyrtUDsd+Sj19Jw9di
M5k3JhTe8l7sH4UtfIYsB8RxTeSl+CXjZ1e8uhcY3iUEx4Qt9Ivd93DNt3lKxMpcF9A1YawI1abI
++4IJcJVBxp+UX7EkaVmjpdQIybR/IfjdNTEHuZbbtyxxpS8at9OfCs1FLZaVl4ExiSrFlRYRD5k
codZXK59SAGs+sGbOJjeqZn1eHNpPM7o+Q7yOZbWiAijW+XE9U18juDCjmn6145IISZTt3GRO7g7
Am/2aW3U3wcSzbnyXC086NLKejz3JLfkH+cI1V2FSUAEYmQ1A2HvfEn3cwPPT6xb2oGckvqTUm2j
IrSpxnlmNWVIXXEO2pSSyUH7VIHCu9CJcmdxEhBGy8tZuKxJAA2y0+WzxrWSpJHAwKnNz+YCWPNT
3VhhVZxRliR4eN/QHdCiJXNfp5o0jvvabRrPK/FAZNduxRLnwUEw15qeOSbQGgixcbG4NEHtgol+
WhYNeQEZJfCSfp5kXHYRujHbChFuyDdGHxVD8mMvMUYeVekyfmrmBdLsHrLp7p8LGQia754Ytqn+
hjOygSLvmFzRBtAB4lU9RbUzwwW7TGhXtoRE3zOSCMGTUyVbKxwPpEs+UmniDCNFHVMkD0oPffzO
LI/qL2lGRNiDh9jhgDsVMmfBT6X8FZu//v796IsM1uKlToxUANqgElzK8yzAQKvB3ex1812yy+L5
sUkaXDhWgL5OQFLC82DHyPeH5bUWiczSCbet9OsMlcsC4oWKq/9vczcz0yVuBQ9ZXznHU5dcx8hE
JYIVnCYSfqtQnDa4JjQHuG5txuirMoome/vhbOuVig8c/Gl1f4EPbPNU/MsWPfoKsqmM2iQTYWfG
QZ0M4gbAbguvzqnG0qnAhUEJUcXP49VHMJVhfbzaeBp7+8TcRHr0tMr6KMO+2LZlA6IwNEEwE8LZ
xfRznacgqsaX6+SfSmP99rXP/qiZFzuPJgxxDRL/E25gPlxdoNIUMuCkRVyhHsxQGz6o8VT7Qacq
Kb/R9M3x4102k1rvvPXtFZcS9s1Z82JtwEF0ak+VsgF3fplrazqP+dqAmz0ZLRei0bX9d2MCpqI8
TJCvN8nVoMqs9e0b7TGNdOf8PjtIzk0VFCNTbIA+K6QKzsNY4KMa/2rM6NPfwxoD36V7/O/kOUIU
7aVsjyUmX/lkCC+QsKmoKyi+9iEWh3LFRFZVH0RuE7JIpxkw7k2nbi2Cfj9MJN455m3g/nOgTKJK
VIwsntT/jPWjPQ4ubS9zoXB2PLI3ncmTX0tIpSAB1/cSMPxSjizkMTUj4coub+3mfGmq+jrU87DW
/5AtbuQaySMZdWQjl48S/M01Or61ci2CnlVzJgzWF2vzpFBaQicn3ZchAX2CEKKkl7mvdopeWf4V
D4J9usaPx5YMp3fPNjuhxdJz38wML9V6kdfYJPp+ZEZESUIY6vsdiEL+zGF93/zA1nCcsUW82x/z
MhHoTTc9WLJHJ/9MlZZGqLfnYd9yj8gQB+unT35wlvIpFVQKVzhW32SNRQwkra/pAu1XqTb4mpUE
ymsO7EP4qCDAoXdvvvZtxBpLfN21nGUvk7I8T84/vpSgpvTG9YJMntAC/kHay7nUR/M4pACyHrAY
bwxTg2xF9klLu6fQe9CyJu0F+ZuPWv56l4NRyisOrJ1F2ykySuBo6ROyuPDLuQBPFgGbjJXKf54B
LXaa5viGx/PjuxtprXnxNOh2GiPdgaYFhT3EvjN+CkHLisMz9VTVwfF+jkz9z75YAUpGG6lC5icH
hhndRtf9H1J+QY/xcUQgY8V3rncTRLJioMSKPcVSdG8HUGAO0Ecpdnc6im4ZnruFYIBBG7cqenF0
anRhmMq/x/yBqGVEEs7dA4ilCbMYdzc3FpTuReRPqmTquKOCxQlsVdQcSDy3toyH3caqJ8uPYzBe
NbCddtWrbAWJkBSif3qvAkSgd7FRNYmiv1u87zTOOCAEHB5tqrx4UMeVTo5zSN25tnA2VVUijIVn
7575V3G4TfAM6THp1Kl7Td2BGh1p4xfCAKqA01I6mly+4QogjYJEUFlGXY0IifbsH/NAVSKEDiX0
dK11D3nvNkxX6yhitl0V/oM7f1OMV3WO/lBGINvtVQyBEUN10kMYLfURXIs0ZKVTZQNvyY7KpYVR
opEhSz4jCRsDDdu07VI4aUEX1bNgKV11Z38ZU+5347DzFiOlY+66myCpVB3LsZZTKn+rIgMHsTnw
DAdFMdpynSYAbfISMJb3Ti4WYe2Tb+R653f+2jHCxwjbDDmFmRiBaFFq40V27VEuWgW4IoWOrWhz
lDHYyA6+tK0aWiktt/VH/ZE9Etku7eYEcHvx8F1zyINLyxjHddOIUcBVZeW+qKzEJwAK1t8XDDB2
TJCt/24SOsLFGIm9UKM4hIZtVZwd9ZfkPKsE3mIIIQSZS4j0HM73bL/IOXu/VkAXaihnNYTOX1VC
pCrUimY0MROfiY5kxwn21+jo+526RxXNbHmxTyEAq1VyJM0ls/eSjohyNRQQ8qFMxaWUwx11/CVf
9Nix59TE3tCefSuHoDHZVVUjY3LW9bJVXKSbaXWUk9Uuvg7NXxRj79bIhn3wsPZtzoa9YFcT+7SC
HZqE+S0sw9qL4Q9+i7ngRK1hQcD7sITp3K3R6mjiP+eGk1Aey4l9PoG1GASjPPHvJ1v2XrAfAZ2t
3tLm6SzP2fKniKKBzv14TJDsbNMURWo5PEC4abPrPyb0uk5qwsz0tXSzWGHGSC22HyqL8rSBVYRF
RvmY7tkNWLuzZUA/eFfqaIlJU9kkIcfQKspespc1WAQYDr2z93cZhrifQDmQ6m/LMd+CviUPFAom
T9ekneS1ySvBV1lREKVFx/Z99EHu3XjWPrdBAJNxDolg+rzjwP0RuRaGI4RJ4LWHjNjqyvfjj7AZ
X2ZyFWQGImWngYTRMeccGrL394pR+ZDBV9Oeu5b/of2JZ4CtIdRPMC5grL0ily5YNmKo4NK/9ifF
uK5YpGTgE/vfFbZhmF2uF01vBqmqMQL6hx9RKbbdIMakgXBmGSNTwU16hgwVVyMSWrMl/AyAfwVD
dWSitVT6Uz8ZG9og04uOUhBg1CAs5/wFLiAJnbwoW+woEVblpD5MEQPCCoA4nsGV26Lz0eZVSU4l
rn6xmAkUfcEuEeRpyl+61rR3OlZHPRr+1bH0Q1gjvyPGfW7IWIpfOVtA3vC8d4Ad/oM3fUxcaAnr
SpDSNESxQtCnC9PhADcePLfQEUJrx8VFq9Jt32Jd5rRsOfPHzAgPhFxlfIrrdhLa014NV1a9X5Eo
aFmSlOM6ICsR2Yu8eU/9L9w2xl2k/S/iFSXHYyp7WL+PoyF8pWA4kgGnKm2j+fVxZb2QCYDbfW5p
sfvZ31OZ+jriVMvCfiWTcPpmr66wxycmo/va6WxmdfSp27crtfSUdst7HS2E/fN8T19Io+Gf8g7c
5g8fkhOY9CLmtEIuMkGPJIDX8pbLf1VMObg2bPi8o3zIydO+2q4+FuslHurIb4KlTEG0RnDFh5Id
ktySY73H9IXOU9wxA2Yo26ZgRMPJEz6vW/wnGu13e0mtRAJ6B+pzvDusAEEBBBKuLgKdxoFiwIEk
B1S1e8tbjP0EyiqDUm9b6NwT/GpsCF0LWRSGUVHVUxZzcj0yXLXokzmmihVpJD/9leDU7SNN2Piv
ASlYU2yp+JsUMm1QPeWVp02tocWn+K+sD04Yg/WKHHrsIaXJiwUzkwysVPe4DxoWFZuAKHaSiGT5
ZMswexSxB5rNPkCLFaHpVuz2n8VarsUDIoRrvBqmfcaVq+1wefYMpXHFCKEzrmrQEfHCa8Uofvn7
qi0CGorZM4iOEJ+s5x94EuVzkpmXEDlVcuZDA0zARrS4Dt563hbVoTOkniSECteBGnvc4h/Ia+Dp
lORNzB5KDk6vZQVy6xdzA30zo1PnIK/409e/WU9UDNYhW61QGbl+JMQ8Om/Np8u+9U2bCn0gBpuD
lDSzVE6vJc3TuM6looCj1D1RcLDfNESiNo7KR9/5ViUXiRrd0SI+kXkko3Jz2keCJXE6mgdAoJSi
gvVV/+hlRnXbmNjQYcJv633CVFKJnmfqbV9jr4hEMPSZ1zcWF7FGpiyckA44l2ThQFaVA+YlxcYF
7wS/L3ePQoj+j+1eBnh9q/ixPWMiKKquBVwODeGZVp8F89vy72ARYl74VomOtFvxNgY8lPSIopK1
QthWI1esfeqZmnjYOKfl5R2I9jEukIuiZlJRaXqVQpxPUB71MkPnVSdmGiX0RuYAMKfEGTCdGpeO
ByO1Mv4gy7rDo+MZj4uuPvEUU3tBN6/IJP02zU4aj+wFDfD7SozwvlX+bCa8dF1Or5l4FCygwklk
zGz3MnUc9SsTmIfp5RtbthE1DifcKFl2kT9a3dV0OBG3o3qkE0DmIUXGBOeZnHy5ajf7i1qbisSP
YwNeP4VviNBQd9xOl8Upf1pT1X/szl3J7v9IXTm9GWQzufaqGPqIBDP6g/fKDrrOXF/jY4Qa5hJr
H8P6z6sw93gaBDuvcobvBP/2o+gNfEh87SrW0A045lo2vf8s9Nw9bRSLrSx6OGWZuvFZDWhEWnlS
Fx3++1tFw+iBn6fO4Yq9QpKSatOUO1Lhw3xiKeNCMdPVuvGcrlVSUU5JE8nsLB0Dfd3QovPCL5R+
OMTkECVA8/vHu0G8Cgytll4LcUhaTETT0+JsajlMktunkh6k8l2wFFp+sSAG/pqVanp3jz80Elq6
LCaNONyq91+yIL8Vj8iqnOhCXS69nHM29Dt3ZB/VD/TAI9OIdfqvQnUaRA29VuQpQ3xx7sKpbBuM
44x2+dSWTNwODroHftT9ILeAyurt4Npp26n6zFCtGta57YgSHnkcWjspKQgC71qWmSb/Mkkj94kz
i/hjgVVeeIgXBVUS72gDcg20Cr1/uuOcTW32/uR0SPB4+2WuWTdi1+skpXR3G8lCJ2ry4XjofOQx
SzYTVO/MLqIzJwx0WeCuCzc5Qb1q/SBO1l/DTV8m9XMPB6hs6iTNW3naCB2swerz0S7LVGBbgX++
zDmiFXc1SO4FlpBINh8a9pabpxjNYw9t0Er1MVE3g+OlR00Pt6zJTZFfwn3l8+7ECaZ0QKuH1EIu
TtPqLis4jbvWtkjwliXm4JbfIdm4J7AX79c7eq/7/5czYWT0rowNrstycRH95S6762Ecp03btuBM
AenQCI8n0UouigSntwnyusCu3FOcy9gyc2jSUq/JDChfFO56eVQQNJo3JFFTQyNuS9mNKwxDBx/O
dCNrXfa+Ik1AnPf8mO/ppZ78NPhRS+nPDtu9PoyfVigorWjOvLkKTF+B4vCBlN2TqMMNf2eL7Zme
dT526hLo3jaUNGNzI9KqIG5t2taJDx3c5qQVngMA1ntkNS2x+gIf45OcqETVtr8rOP1zg5GJuQZU
ZypCJOo9Z01FFlPqEMoavyImkX9HlGWYq8vjOjqm/QA6/N5cJRzGgTqLvBZcQf1uAN2UzaS/sAug
pw15ZhPX69IvhUj4z1ZdYHMSK7RrnjIVoYAkcW66tVpqRLcjigtvKYWyto93VWyXk9S8qUQh8FEn
wOQbb7KfRoDRSfjKnRJ++moi/JPzrlVcSXMRmU/i+N1Z8h9Ny6tSCJu4hetMeH4xC4S68s+8515R
D1wE2nxIXN2lMzyC0S3rFRPd+2ER/eCgiMH4dRlB2fQXTO3YzCBhYJybWt5uJSgCVGVY28UPwhL+
3T/IYHJ9oRzXk9FnGWOTqkGKmVFFVW5foXvBNXRtRly/yaLqQAJVF/JN+lCf8HPdfN3nIiR1VmzI
Y2sxP5NtYFvMwXPYRgBroPzzheRjGgCDYZDGiSn/dHtivoYnrqYs8SSeA8Ra1MQau48tZfsCrwft
cQHjvZ5LDHnhXhusSD64R4v+URPqaro7OTuXZdxKapc3hAATxVN5Jhb3CM+EOcslOdN7QNXr4qAX
KaQc9cFEyIYQmZuJRpwsENBnyJrwF96wK1adOpjq67agmUs/s5SzCUb/w7Ohbh46pZIgNx84vJxZ
FdVeBZrHsAOMN5/ujjc6t8hgPMWScPpeN5cxrqYPFg+DrxqQjKZ7VD4ZBCt9nQlebIIe5CVmYmz6
Ai1BRWd4R1lWj0tXf+NyuTLhmsieQJEEDa2xPrE89oVJ8fzKKXAgINKnTtWINpbbiGuBw56jR9FI
rgH/7hofCfvlY662nbUZcR6whiTfFnIVq4pWnPq/m6uO1lAn13FKHnCzIETisBcuNuHjpIHMgvCM
OZj+jVPP7Bzvzo/OtWOwHKW9XitJW1SAgQcryo9DifDCwb8c1c3WDVPkPyOVZa5ZJoDJbv4/eeOZ
cfYvUUPzfce7lEc4sJlT+jg9KfC9lafq7a4Pc41+VA5Y/1S0Hf5YliUmYYStfR7rBdXp0gyBfOOV
oHhJSDz7erMPWX7ybDKhTuMo47q4btV32wjumZ9TYZ6rmfv/Oj+dgXX3RLRbX3oTpoFWQoxVlKyH
eR4eYvPdLPCKVVPZimJnBljgp++WY9Ngz8Jemzovdp9hmm02c0pkGsoPzCtN8avA9iYEaJlhtYam
q6jp6rfy9GbZ/Ysd0qX2yT6/WqFY5A0PFbdDd++bNVFJSoBfVeqZKRqBqV85HT04mwsHf2ors0Sx
LvuKyByc5KOdrk7zzdsfSh93yzzDqbK7z5qTVTzVXa4wyBWoIvdTEfiPe62ol1/5hnBHu1Elo0l3
Ys8a/BiUouH94Ue+EVZtoNn1ocKcsrrdFJbqz6zRL6KL77bavrG70TMe2blavh7uCHjlXUrx+BuY
6J+mo2AJ9R5wu6d6DIA6NcVNv0HxRlBmPFZrxJor3iWMxSmvZyFys3pmXYbY7HQqzz4HG2XMM5nv
8AgN6k/wZNd/Tcd07f96SmkDeBi5mlbKGt2vEfzlfUXLB/q5UMmJyggvtje38Gy2mJA6G9dpr9uZ
Cy2La5fH269w9d5w912kViQ9RF/K/8RRAODmSCyXhzjEhmzy/adOKj09u8NCBhIpjc9RXATLrcOf
g/zeNBJw4QVKmoKwuHXiomtwkR6U+7FFf+3kBStxpZoCSSHJn28Y8wT16TiQigUVphpVMTO0e/mM
t5YIkTw01QyhH9gaJNe4H/hzWkC8x2dpU1Is912+go0qQWDM1EVzjdZYv+5pZVLELsH79PxGddn9
kUqZezY9gJziAZamLdCP3/M1XGy8ARyIimjSfWC6pzRXYsLm7a6/+Alj9+eTWn58mt6Nora55M4J
HSjjhfPO4vqIBXkrQCPu5fWIqcl61RQHeC9+fmuiMZG1Y7Xkjuy6RhNNbjDQCRpjo1/enirKrsmb
0OPNC2tQpAZ7CBxTGowfxiJ0bUeDOoN+BYKhXYj8ZUSQROjV1MEy3bXYATPOrgQ4A4br0+k2lRyD
kXDp5yvH6WHijmVS6wCZnqZyg2dXq7XXCEq1BxDq7ibfqRbUnDobcCsH6rImKPyIWfSJgEal2Yc2
7p59McXaXz6OheKcak3nrzeKWY5Lmbc4NBQL3SUONoEzGlTiPLguT2PvapBH3YfXMriWHr2CANYq
VdzuwEGeLMT0XxwndyBWndqDfrZxbN998yOt7VOP+6OLOcWiX1LM55K+gAj7b+1jXzCL+DcRcPfA
xRO/dKpqrB4OG8p46ALSZmIHWpeG01/nw/5rlqhaAGZ7Q3ubcv1IoXGlErbBx3Q3UB7VGqeNFCF4
BA+e9di9IPMrqLTDs9/sDmG4N4T3+tko+Zaa7eMmpaVNCv4ki2ID7Kdh9cuOuKu2IDN1HpjfPBdv
jjTdZd/4rnprgKVZ8hNDjOsDwamstxXa7dNJ/kdLqkbiYbkL779ghspJPJpwt1aYQJTuPTcfybVI
yTdLtolSdcGtRd0U3sm5Nq6rIAAwnXPVHRiYyZRii+MhnZlSFy2pwGkTjzj3IMWlFuRl1Vlq1hJ4
2jR40/8S2zxCOMSOSsJCikXKYWLJRFn2EJ8ie3YBghK4eXOYxs6z6snoa/lUiMN8hdg+1nf1i1NQ
xQrF5fYdKM2b0Y9HW3alqS6hMccEPXqUT/5Fv0pnKVENgfduRGlZd5K6lI5zbT+E/fYeDNMQzapF
fJa5EsmYv+/8witV6jDYn7RFO51p0CNRpHuTtFrK1wUOTmWh5VaJljjRW9cIt6NYr2mbXPQ1PgRq
IjHUZO3tK+h3zzmIc/3sgUODZZGURL82zSQ9kN3k9Z4PaMqhR4Q56kNa6+Q8f1D7oTic9xMsMRAC
aIcYee6ohoFtQLtzC1fLfWQhQqXScz2hLVTvpKMPB9Y6Keck+6WQWB6j4ioLO4SBCfB58PJzF1Ij
bcRXndjGBq8GQeeO0TAUILSyEQ4NIUrHPNa3gsUDiMSi2Xdj48/QH0pMvQnmYAc39KNVlDGxYOGJ
8h9WeKPd10EYwzlFE3zE5uc4r8d+jYF18YmGMy199CC/UacupwFYDU9QOABZdXipWDKcsizcw+EO
bOcL0U82eoZMLG6Qqa2dAnV1hT4sQjt232IUoHT5FjNhOTMofcHzSoJ31x3Lr3Fo5963EtpQewd4
Q+U4RCzsBAxNdNtvEJnx2PnZkaRhDTqzYup9wm7qoid0cXsy9QwaKsUsjMLGsGRCdsgUfGe6aWeD
+9NBZkL24DPSEGQ3dpdNmJ5HLEJqG95QYrYc1CRZ0ev9tKgDx3pSLFd8syumRkhCRTBzzIQBQ6ed
C693l2LJc0EQ+YgSO8zVt2Or0lDSjYj2IzEOvLUVbCzkLtGYOyVO4hEgLENvs5gVWWviYV951i8B
h9NVWN8kG4L+Z0buEVr04WTyW5d58QOLjlGQXOWZhbbiO30eBVWoBm3fpEyQs8eteBPX3CFSadI/
wuMDmpCdBdFoYIJ79wSs0W86qcKuy0dyU5xPSQnaFSmgOylPUrrcVX/uBjj/cfv/49LXrK4ciYk2
UuQYPlX6hQGpx6X0GLouALmDy+TpG417GkKCmWl95dCFDYw6WsKtqLcl8UjZAeUBSMN0CFFws/jO
VpYL+MsGMdqIE+2PP8GzaYKZ6U+KLYQM+dS2cexb4WS92dtRSBo168vnJUp13AOB0jRHNPvAYAHu
0mIZALb04qWU0w05aNeDQre9ezhSy2jsYBgVPJdteaF2r9OWcLt0UOsVmXqS62AeC5YK962XJkD9
gCpR5C+CL67j5zRvfkpz+k7tcvTrolL6QAAFvpVo+rXjgjsa+nzrZtHUwKiBYhha1EdD7QR0WuTL
1rqo4Uqp0O/ZQGWxUpA6bCIV79DZubqWHxLbSVU4s2LgM0zcP8zJ8AxUApNPGaiU4qXvFyz5dEkC
c9X7nXbEM7aDAJBPaEYM7sM83n6wDLRkrqnki3D0CpjZXWAS54bSc7ee64C9K2FnGAOzsdscrkm2
0NSe8r+/JtNTbwTnm9ZKEJ6BtLJkfHFEftCH6oyXqw+0YWLoXZ8/ksuso9YMNsaBQA9aC3G9iX17
eLW4C0eranPK3feSsghBNUasM0uhpT3j9Eqg1NyeIH4j8b8TZBaQnbMsZlH/wBFVcxGfJXOB6rn+
6rCEkdaZc2wUKX0R3fnOC9qkCwK6C4vneTqZg7eCthr2U+2Nk3Dtd34wsoCkYInvfz2TkqHLouCZ
enocbck8V50WsNUuiEtiMvuN8r0HiMMn2rLYdPFcoq0O0omLz7/ZyNSOQkQmM4yfBHs30nAnXyxY
Cnm4DmhtY0YHBOJrLwj8kwuiP18GBhDlbaBoec8qBAOaSdHCsCI8o1pFNKf4fToO0hKslDYIMUxY
A66BZZk8JcaCAELCEczRvIj03vo/rkdpnKPx9Z7vEKKzeowGbwyfNIef7hzswnbt4UsuuLCzJh2K
2TxuDsJb4yZ9cvZYYaEF74ualG8R2mCdx0A38IaNz/+ynkykn+pEhKgSoEA64690Zrva7uRHo8q4
a7GBYTFU+lth+4OlGbilhrC7Zz2YpwNbWTyT6/2TRJIg6Xe/tpnh9q6/v2xrqAFhrRRtyKLlpfzG
NKQc/IVs8deiSwe3mUdVBnXETCve80gP2BnIEW56/GPLNuIwY9s+IDhGnfbs41mAZ6MEv3xp9iG6
M/b+8hKeXMxKzlk4egdnyrg2ans5jmfalsvUjHqUO7nQG1s5SNA4v2ltye/li/a2PJRfEwdVM83+
YLXzrT8nhsxObKXv41+Uc8vOeBsB2P9WIgdTTSTppp53VaZiL8wxT/yUhDRm/N00jDVorjMEs6Px
Q8R1cIxLcexCAtEy/INRrlsKhbNoi8ckDE+0DOEW8o+wy3usz1XDf/S2ZXxrjvSFPfqwSHgGZjNc
s96nhXKAL6Ia/+tRCu1dk6jG4TVgDSkvyqlGVaihkafAMWP/S0LViKIaM5emVxnlyI0dfUnTsT56
Wug3kZRx1XOcm3t6B8t4EiVZCJpFRTwyzPdkMfYQYsMONBtiPNsW1oUoSCfal4QIUarqZtULQSq/
pKYb5LO2nu2FbLDB4DoNp3ZlklT5xCAhCY3EWg5G8M2SF1eXsL9asryqcpHKWcBL157VyQgTN13W
NQ+nEMm7pHOqB5BBAg9LzCuyGCepqdgx5F73ZcRwuAMc5/94XCQf5rLhBl5hKRZOaNEYrMnuuSnC
YfhRqsoDu9RSo9W9gzv5aI3ibNcnmzrcb4myH0SL38IyNk4dRybdJ6/9No3hT6+WWa1s7/kQrRZt
8Vm0jEaO2R/VdJwTiKgTEoOlpHgFnVt04uIMmKozbgpXvJIeonVuiAiTlTedrbNXqi1s+nAPPniX
rBSresc1tkoHBwRMIeryYJoY9kswjpmRFpwzS1y/LGpdRHxCLdunE5BWH4SrruUbeekBCjTuYGuZ
fW/1GIq6ra8QUAI5I9BKXABU48NMJnIuVYxkx6toQXF94LDLtp8DPeflgRdsOY6nYGhYTlv1l2pq
PjClaPIpE9b6ndCXEpev48Mwb9kV0q1HkVqHVUFgSGKeJcHKWRfQ6afqw8r6ycqfdo0NGP1uAz38
btXnik/FFPfiNj01EQ4E0B6hxRHp29t7w3TSsT0s4lpauT7Vmg7DwJX1FegZxS+LHZ6ZuHVdwzFL
rYpWDi210zvWJOsZHeI9NTAjj2K/n8ZQC6p12bh+WG0g1dMJMKQF/jLLkKSBewAKHyYKTeON97hU
QpCDvmx/NBz0XdKLfJmXMsdSogKPlloNzFDFkCABOSvoVMk2zXAuzM0Q4I5hyl7WV0dA5g5l8Qbc
DUr+8YR8vPlZHrIgJjEzfFtlFSzzzZi3dc7C2mYZagp4M6Ro+1oaCHut5k+OfC6YDzI2AL27roAs
LtZrvLEHzGJXQLamSyxyH3y7bo4D0p6U3vcZ/EwUS3Dqoyjgf62Z+68KgPAzEayCcYFUnKCdm6VJ
MoJj4SvMeFRrrGIthFzG2VM5IdI2IblqWdvA+msL8ehconNr9ZtlHylimW3er4RHaY7AKs9pWnN8
GLI/8vUX9M/fi4XhmXTxuT3fxF/yqfdkP7M83LBr0CuKY8EZ6Y21VuAW0T/SHnc59TAAYLDfERKW
qM/nvPrF9dtrod5D2Qrpfy/djFwZX+f6Fgby7mkcSzbVrYIHCEc1nnw+G9GW55/xzTIKqmMHSq/r
AMWt9QNT94F1u4UfKY1dyM2L0x2tLq3QYk3Y8V0qAEFTAXwr+tbozIYqZcesFtD/3177ItobjQIx
bxUpFA38FdgFI3M/1P1Y74aAoromhsEvlZruM/iPL3tKhjdJA9WEIAIlSoQAGpALWpr8nEKbGPks
x3QAVNa/o9Tr/yTCodIOU5NPAE1syAoEcRp3KArFiRVSGUmit+3V75yj9LTBRBRgD69UELSJDO7U
lea9gIcIoVACkRsC/YWO0Syvww2VGITbVugaUXaQB/dVYUL8flD3TwyVY0zxSQC8eyJ/2OmbUxde
klRLCZS8BSvmGSxlIOxZyAoyvm2MqDyhEfEKvygSavo0PcCL6+xLgp4s8m62/Gtm1QIOyCuDD6dy
cdsypmFWrDV0ySHANfDtanrtZ7wQ5k+6BIBAGnFN8Jn6Be2hQyV8lFKPqE/NRtqgVm9anF9Qckiq
2PR6Ipaw//hdZhgljF+53/C8cRg6XHoVnBuyw/hodtar0F9G+1AoaYt8+fHBiE09KVhmeSNl8Lua
qqY6182C+XZuIYWSHjIGnevF9bEB3drMOKyiGfz5ZImG32nAfZdI6IYxQ8Vp8ljXYWBqXFZyVmO2
40oG36K7IzKNxNvEOPLNi+6w1GZCswGHNj0ghI8IRUH9XKftsxiVIRiY/A2d7x19L9Zg9uQWZppf
KsQSs/rzCeuFKw8Sgq0ccQYLOqUj4l4/4NXk7czBrFRSd+DgnBUbNI24X3duqLwkbpmGajTZEHNV
XckZVJ4oKDLltNpjZSfDzuj2wQA8IijZZX12zmrdJhN7IHK52wZn/jJESxpg79sQhV/hqL6JwzNt
p8kyt4qzKSRPInpnWOLSeFDqcknD3b4cncXdt1+iwVLzWmuFBTLc1/1i7VUg1sUu5ffyeni2xWJr
Ugu4ZbwRvPQg8Fp+LgxmZgrNIWwRQKRwnFhU6peL2J3qkzDQOlbvA2vqoqU4aeRjTtFaKM9t5pmH
+5KRHd0kue5iqZwLOmIHKfZgNItg2TK0RcoesPaH2nUiqCoz05ms4ItrdyLyQnRV6J10pSJRceLJ
DO8Jt7fi2WuXq9/nfPHN0em75slEBero+e2+HGltMQmDUncm1ovqTxNkXlyYGLjJbIh6qoEgJxw1
Eb9gJB8/ufRiZwluxsGbZROVWEuT+aWPyy5AyeUB+LoHsSQi//VqOJchKobyXhOUkCuQH4VUX8Hw
u6Ke4DsZGD6NMXPZy2b2TT+kOYuZ7JAIbinxx/pmVMacm/Q/quyBczj/n6DTTe6y7mwB/9aYFg9F
ZBf+c0HPHDvITGpeXabKoFd+sRHFhGXR8xkMjXDACA1F0tQ12uxGsl7InXFKXyKu7dpBaqcBWYdv
cf53QD4FgZwoMq8QW9tkpkksB0wIVENR+vGv6U9tE0xvTHCmtko1iKOU2a5BaG+SpWanQpF3EN3G
nN8MSizDN0Lr3tFVG/fstPiQGjd4/eAbdLZE5yWSNI5es1MsTnlxmrwxawCjOB719n95cHbw/oZ/
EqLEPaDh9ndkmn86L14bdHnwtN3PR+w13Q8/QceKlcz3gXh3GNS4MKIJoVlqQcSfKlswqntlj+Yc
/pveZxbWhney9W/VCirli0nzkcJpLkiiR2Th6V1KmhAFDe/7OVYBMYeW5LluKGBGobumRe5jZOG8
sg6Rtns2uUGv9WBonMiLI4KzTuiAfmGmR3Zhdkw1T6xaah/glD6heP8SDI2qr5buYhhiEQatUKZj
SDpVRH4YMTVMMZK+Mz9KCYHtVQpS7r6RTPqeNFepUSCa56+owJOBkRiaQOuLfmSZPEqzwyzJpKqo
nwJvap0UFUhDxw+KUTt+CsTU4T0NNQGaaj18KBceYTjHC2h0CJ99nylv8wqKZheXN+Mjgc26pdRb
nc7oHG/jEXP9FE1FmluAmnuHhLhsZua/hjknBi3TtHmuf1v61CXI4nDdveuC3jGMr2usiPZulcXT
6ORLq56hbQid0VyX7AdSVEfpn+QiWCmWo/lylPlylztUhSso1GqPKIIk6OgnKEaznDGvQF+gXgaa
YWbGAyBBIjYKMcEKq2zx9EeZ4ippOq5br8AV+kDT9eMSaAdtXc/UffNemBgL54gKmQ83HjZv/ye6
HUXs0BwBGTFby4bTtFF1Ptt98r++kv4U09SDLxzh12HJDbpbBmkfI5TIEaMNZQbgwD0FglBLHAiN
D9jbS1ShviDBlY1I7TMga0ou5vTK5hBLbIs93ck+qpTHYCgtWynzF2M3uFUpcRGSQr5e6q5wTs3Q
dvR5GpVSHE3UI8Rfjywrdh197JLyZ5K2hSoPuMgJXtH5xvXIPYFy3O7Xn6EisOGks7xNqehheVGu
ZXz1CgDmuaNqff88IQQ6fQc4sL+XgxAeORcxkNUWz9jgLKxfl2s06qYibOArLEEdZRpboeA1C498
9J/bsCSqUvbpIAIbGXqjy5VFx1q87TR47lI5GYkxgyCELH2n2Lk5mfkQz7jGHHSjr1WalctOq2qd
sEaxpIaMaZ7nSzjA1V+OLqUsteOj4l3KBv/+0EOyMax7NQYbO1bNdngmZPNzIqQg4NQud6ZeIhav
QLxN6SljtlSay6vu5tCBIfhKq+KenJiCkxrNnY45iLeqADAQv+LD3IJAM5wewMOFl/4j0htzhEgJ
+/vj/E95Hn9xFOFeiZnnj9LPOGe8Fb8YCuyi55Zcp/ngcQdt5radm7tx+HUNgWuQVjXLmruzQ6c6
ITBaJ0hVERZNFvzzGnal/zjFIQpEb1Y8xaGXLogJY4bvMQAQZx8jXdlZs+eOdDuxedEs9LVpYo/Z
k9PwD4QHGgHYElI1+FhygPtnPl9xgGD16PSPONLf3+ETouuebr/I1Vgyzg4J/3Jz5ZUnXXlFGgEC
y7lG5WmKHVK5oLGVDPV99CBeFMWHuNYWMqzQJgqrXIobgkHEVynOqZpxd6u5Jux2fNeERmF2D3M4
GY17lnRs8PytzDpahVoMiowlqS2jP8gZCa+bNgL65ZOjNQinHEHxeLS5nf+rsNtweBj9twWoSWYL
bak73eUEa983n4Tntckw8q2DmGNQzRgk8xeR7O5wNvfKon3aMbS0tHDZWGRkOOICe7MHh6+ckpmU
ToR9iNDYlTdQ/V9pBbOmeacIxxGe8pVdT4JTCmhp1qUM33d5YcmWRGh+rXki0v7TYt1Y44YYQ3O+
pwgkal1tN3u8V2E6KlYGSPHV1Xj9vnqxSbzJO7+B5uqPlVazZSppxIkLZLS4ZALO025TXAa0e9OO
DH1ERIi5GyTFUitHKyW75poKy9rLdsF+M5O1rsInenT3iQJJECjCRXJm3J3OQMvHp6zO60PBQvlP
IcPOfawfZ9K6px5pmNBYUk5F2W5cCOaSW7up0qnBgmz104IKEwxPNE7W0whdZ9VEzriT3DbmYqvJ
wDhb/11YYvTtVr3G3olWIZZAjnORIQSgfjEvru+lvJYEeJ/ihDhQJwsGsclJW63R3mSKybzInhXA
DOHr+wzv5QIcJim65mdDpO+H6RB05fsnzz8A4yBA/La80Fe5/QedI/Sf/DFm8YO64e36iFExylF1
rXIMG1VKZNpj13+o4fDsZG0RFVcFxIchNOsPI8mm06CgU2ypNnDPNsyvaJrEdYHeAkOxTDXbMJMO
3PpKeLD+inOKncs1aTlY8ytgqAv0Q94BCmQUnKP5MNMc6d73YqkkSsban5/c3g8IKG46pDyQgOrU
hbyMLx8xtUlWNIU/wMJ5rGDC5H1xIGsoOLw2GiTnSTZHoY2Y3FcEhkDVFh7yxIqfPKW+bxUOzQUd
8TFXhXQT/5NSRISWZ+0l/ZsMPTwXtigUu+jyukOF6NiCe+ax9ooXDxRdqFN6PkwopF2t1w/03T4V
7g4r69FmalnQoVwpzJQWhoKpAhQeNc6Dokkz42VE1/i9/WOm8LQPh2BMvN9A+rc3NghB54PlzF9s
ElaRs5blQ9GoAM3Cspd+9a4uvZpQqEmNwZk2IuncSOF0vY3n8diOTecy3lUvuCbOzD5FS5Fnm6KZ
7A20bkvXYxRy8ZTNAuaK9H8ogBUM2TbA/YsaIT+nT0YqbjaCmK5DjHCwDJgp/1a4FFqVyqwXcNTm
gym/fgJP8a8w03Ods3kM2gkuOmA3LbDTpyLpT4Pxmhnj0tCq/+a7APnsXrtqsCdeLnGMtaobunMY
YQhRGMvkuN5GAKy7ed/iW7Xrq4hreoPlp00cTBfhYky08kNDsRx/povgsXPvYwA4Mazd5cnEbH5H
O4ub2bBBTFwMz71hldRIhvC2PtncVPqumpT/v9RJu4/yR6ly+k0UFytZyzTk5zEgW40dLB0A+aO6
yNwOSK71l33R0HJGtzb6YoEDGtmBU7SizipYEhAEQbYXZcMdU73OiKHm6rvAmG2Ry36DtdFGUEuV
xM/kPOA6s+HLQKDEbGsFX2m5Y1l0QhYeVr/qeyxbz6i5TYucXYVKwExbDHIscsM2uF2u+omeXyw9
wLEHxmHoyQ+4WVXArM1NeHdstyr7RkNc6KMZ4txxTs+31eqb49ZSiRSu0GFD5rfO9bNJ30aPPXDk
4SF+Ov4TJKKxHbXEFwgd2V86DftLI/mYMBqcew8UopZtlRhytxac2UCfrS05XYMxz7ME0Oj2wlkm
AdPS6g7FWpBegSJ9qLeWYRgaYgWdUHZPHXE7s3zzS4c5ZNd1zEK6rg5Lui/nsIE7t/KaI3VEfd4d
AC8edZOJE4PNwZ9U700wWTnF14hdL6SjOxO4dlj9++Q8hNbKI125cO2hpbHKpc98utkQjSgx9JN5
EVuc7NJEys/rtiGkOsW0tT+nNkiqIwVtBSqtrUzLyJL5TW3M73yCAPtoPD1SK0TWvxCExd/G/aDT
N5cGsvhIY5JGShcd1PjoZO8ublNxxLzQvlw4Hxelk+XOoUV0vrUtc+e3tK4ABtL9x/rjyKZoM9U2
/GQOlnedb9P9paTR1boXizJefvZusk4PbBzPZfLoyAWu1IzwqOwe4Ih5Z+v7jUubAJ4q4H9Mad27
VoQDQCCvpTp/LGo2NlUKeX+LmHhyFT4NnYX4oKYz1CzO08T95DT2umIKo0dT/EPtZJMZcaOigFht
68eXV/OPTt3685YhLuzR5GtItaIVRKz3rfuWLrqgM5kOeZLpOlRzxgF9AFH2MtBF3qPZwH70h/0U
4STW2igkFrYvo78bBz4aswi+T9ZaodVIzhRZRRNxINHP5KUFlBxS1sQ/4uC6gM0ZeLnlTqBN8ESu
3iZq0kgHZ4hLnD+ji4k1km8dbGxl6Dh9QUD72jysrx99R/sJmStkOO3lYOKmzeZtwmIQzbjWSbdq
N1lbNTUHqyKe6Pc+OnQ7Ww06IXBMIGcJMtPw809dL2hETkYyKDTYp+pm9uA0LMoi2gRnEt4xU8KE
2jlKfIUfn9/pOsAgbNN/ALtqdU/kU/N2xsxjoiFEfWjJNv8i4l04v07cjNNPSWg5MgNMbjOReAON
iVwFuejsOTp6i+OJoIIbPOtcZUBftRC3UWf1uVNsyXYkxTMH6USifo+NHClNzgVSHF+NPKrbQUcb
rkmPGYIcDpejbwnKVRw85kEmRTgxzDVcHCJKq278alaHFa/8fLcwB5b36d8epr4O5djspxnRfEDK
MwMwbjhCil4PZAjwxUfyY6q17+sL2Rfed5doM7k0YO68GoVlf/sYxnrHcTJDjZ0uLfsoROkWRglp
QWWagkNJWY5PbTiypE2VPB81sT+FSvFebRFdoWNJUGUK5CNCORRc+zbE7wkpS6Id3EgTt6YOh96Y
cei3F3tFBRfwR9TAkrPG8heCXtAPRYfH+CMDYZxbfHjpgU4+tRXmHJMM3pM8zQCDDN5pd8D5wE4E
nVtzXUff2OnZIzIwvAdW495J7EFD42uFd93H7ibRxp8L8uac4nVKJAzi0W9PFuPIgPQkdfZS8PCP
da9an9g/jegHfAmGH3/OY6fWlPae4VgmoKnMYB0J5JCuisJoIRMC14q1y9qOOiGVIIqmHZJyYlqC
t5tY9Y+jFW+PgYYCVioE4pmUE/bb/cnH7tK6/Q7faE1UEIZDWID0B0FTMHvi0Ey6uXt3nliEd4a8
t571s0/abX0E0N+SMNJn2G5octw/V5gHycUyXfzBozq40Bztl8rv+QW68/Cg3Gy+yfjsUGMx4P6I
hq9slDmYYEHZqbzFUBBNMQZfSyaVSRZDO2Ulb0E/L8Ywug1fn09X6tqBXkLLNnWPcFv7ZM4fVbub
RaW0t82PTKA9p9TT5JBGCD4zefI9HhIvpCgthJsa6rFoK6Xl9jKHBiNvidaPhfo7pO1ouQFBUmz3
zZQI9MXXp0WKpzcu2WNcBJsO8FsYPe9Z9eOERMSQ1puQSugHJVZRzB6VzlSOTABNykdO41Ug+/KC
W7L7NgdF0TOgkTrNp/zP2QbUsxXou0CDds94ugzwXmJcTfIRzKi1ldDKG6ZKPqLC0sy+X3nA9JNc
/gPPIVD4KfhV8v5rqGgeeJjxkM+tsRUOX0Mcqlz/70v9CiGaiFQ84+sk08817xgnEyg6l0MTaSSJ
K7DNB9QuK89BbWH4BSYP0XpoTt3Wna4Fb9b41Tzaeu67Ke0kx6zwmrlPgiZ419yzklNu8/OAowFv
2CDfuaU/3kdh6YL85uzJyCOS0M5OzE78rNUtESnCb/Hm8G0RCv+rhgxHRZlNllfVXWrz0ppuBzsd
wveo1dCdLTWAXzdGqGyLS2f4LjKo+bt31crVB3TeH1Wg1lF97AoYh4xJJ1O8aXY2ecHVsBDXymw3
AA8PyPFg0H8cw9t189y8aGc5K2Ocx0Lyl42wwkIxPQ8HxrbO+CZ0wQFnFTzJl+OQbBvQqTWSlwg8
cYE9buCS3q9jaWHHHDhi9X8MsCHZuvWd4Qnz8nF2WCwUB996fsYPumwzHJ/D+ifw7qigbAG0bnTj
Aoq/qQoWIuwFSpPnZOOXi+UR9OyBaF4gTqAG+pympkmQbGsppWqxixxjZo/5U9DkTk9yzg4yTB1p
znoHHZ2aYQkkHg5n35e9ydNe4XpwzYEtL8JmIqPKkYh0Vz1EiEv3vzu7UVdeP2ooE6rJPVr9QLzA
CBpgwiomhZPvcqotpCDCSEiSVMo60SJSGd5izaNoNQMOckzXtKMG/mp70L+bhlQdS5ihbjT1jViW
2D8SB2CAO6eM1vJVkyjBfnk/KvC/97Nriy1FboCNKH48ARNwYLC25Z8xulNw9T2NHBmKKx7FrCq+
wZdi0ylWz4QW+n9sgZLE+ut30GoGAIKyG8nz8iH2yDCE4Fm6EL6MJdRrt3SBgP7MXsKtW0r4ZTvA
Am2X8KKjid2i3yK2YHaxGZoM4SXp+eOn3a9DajsNUju7eRxM7UhQdtUTnBQL3H1LdGRGJpFvHaAx
Oh2ekZ7Nk2g3KQD5/wC8DEBNdptXi4NOzyiJ7vFPZr7KO8NKWx2WmA5GhkQTLzIFjE7K0AZQC5TF
wmUqXQZVOAvFOZraQNxNa3FDD04GSNPqwt1viTxnmSV4jOZT5XEtJ7KLeevUjtWNkOKNblrUaRXQ
xK0EHp29eYKDaTC1gSEwc2djUXg6tV61rGQzO2aBdtsmTMVun6Z5+HrmBwQXfbPG3FTaW58zGOog
ODcgGRorKTDbcOnCrBf8GsVbQS/YvkOIjHtouTOG5rBQxfMdSmU9BhdeYIpPArzM40FCObhFzQyH
/5MQqGy/npDEBo4NlarDWNYltsrtLK5uWzp4vDMYjS1TecM0+bG4sXhRTI7cl+eueiEgiQR0Cb0u
8OXQcDFyVSmxoX+G3HFzYHmid7is9bc0H/BmTPjJ6DU7NOXhFYcWMeRuK5EMwcBCrj/8sJ4g/XPk
ZJOkCj8ODciLatUxgkIqUpuH6MIMvpMfylYpLJyi2uiTMGwJqalivHxEoXVsGTGZn51uqHRA7oPo
T5ZrANYI6D4zgCKRU6bRoQruWkTqegYSEYrZ8r9q8i0JUKCiSlrYQyhqf5U0vTKFTGq25JeKiR2F
m/HoBr/l69afKKt7PFlLxloknlapwoZPNcYY3Mgl1Xf9Jyd963JD6c3Z69zedIa93iqjCIO+yiji
4Fb0orm+xMJvvh1m7412pvbstH3W7eyYG5e0f7HA5xMlOaPISiLPE8KXo6W+/3nPP1cTXNinBsp1
XIG3XrS6lO4Bqu2XOsINXiy1j27wf/ZjAIsZ0YHt8APCx3BYDqa2oX/9wOBrWJ2o0Lplhv8sOmfR
0g4+vtLd3oHXiDOxHOeWm75fXlLclDImRZ2BnLZoqxlU+0xWoYzBEN5rH14bZ1XOem86ep7+BAVu
r5jwFEbbIEixVSiG/fjyqUVDbjcnbdGgm6yDX+QlmaAG9XRuaVWrDJ75dp6LKAA097IRLl0somd5
vNk9ZAtnYx2nSjmddwhMtvbKTueYa9FsFfHcxt2+0veKAlzM3JkyIp9LpGrWC1bfUxqJ1X/WwSlT
StZRDQyMFcwLHaQugBeDcI+AM4cnl2bdCiht4MPTuSuCkB2RRiRgF86CFv4j5+Oka6FMzV7fS6aY
7lyeyIsJP9Ixkbv1BmrlT5VON6tqxmrOBn+YXrv9of/2oPCDZGfE/85lL54JSiBgPiSyt2FIOqFp
N0N9hrHAllNAutUNOkEx6plqybzQSOmJtsShc4W8Z/v6mKzbkmljWTWy46ahdkFdvtdX6yf2vd/A
C5ba4zw9aYsjtcnE4yjhEuYKiw2ugq8/pVSQ1xY1bcbiRt5br9+d7MCZwptko6Sq/F/oHPPhDA3b
QgedLh1Jtw3JEY1U25uAMI2OCtIc/Xzc5YxFRc7KJ9hOLqKUZw7TsaqWd7JJzdX9Ov7/Bvqg9g2w
TW+nNyRS7A/4IXaX4d3z3wdmqqj6j4WVfGaWcnj4IyzbFQEPVFGq3bfAb5T06yt7NHsiHzMWHty8
Pdc81fdfpynLCw4H9pLS8AUu8cqhsjX7os1UYxCl/9VPXqwqMIryjQQpDOof0MVMdZb2G8hbRz+X
doPOTC/tUCDLYh/7Qh091JG1PM1Bk1Nqu5xLC1vB1L23H1RH6eZgufOJ7jI1ahCHaRHBH5rAOIq8
luI6Cg5qzHmkwIS2eMXxpNccuzXT5W7PV8OK7ML5LgnvLvZ+PQ5fcvCOrj/SW4i2uQjpc3gVsKSB
maZpjDa24WohaFy24lj2fReBO5XLFy3K7TfZBZ+Nt9dY2n8D6Q8+UtuWOHenoaa7NwPQaFRoaAMT
XL2WoF97dGKpq2Ytnotp95h00Z+sQlX8/OQ0shk26sYRQl3r6w3CUsqSz2mszsKINnpW8YimNzrF
mN9otH42EJI92L4lqjycxcEVmvF8iGJS0rJssSnBvnNrZcYSY4AuVmR7g+DwGJczcoUSJzK1n3wQ
3xn/sgFSDtFDkGwLdXyYWX3klPc2nQ0xk1XlCZgMvmSIVNzS2c49mCK1sZCqzdvzdmNHxSovkc5O
3gswwH5zYvoOye63JMslE6ldwTN8tU2rTgz6+ZofSDuXVelolp51ZX313ldsJ25wmBY6oOxsFKxK
nZ8/Stef144+jgb+PLGf7twEWVz9aja0hJdHs5zQTwsuyNraLQcsK656XmrX5EJnvZvqi6CDcznH
o402oRdx/TjVAHdHmaI9hGA32lW/d9+ujV73c/4qUh32a5NE7bVo8UqBI7/Vh6Kg8z6VwEf4XIWT
6iccWOBwabow0UtE0yOWSwOmab3+FzQcL6W443H41zeWUYrp0D89dE+M5DOKz56otozW/9HxdeoI
BLvtxi4kX4awYsruakeP2PJEg/b/zo+WmPVkreAacp3abqYKhjonIKLpYa6tTJRudq5N4KlJdrtc
nvVQ8XVm7XHjbVX4jjZYR4DTsiwdefvtHtoA/BdLcP1/btlffO2HT0MQ7J7ziDJOxxOxa6NxR2j+
+oRjGsrQ+znyj12rqzCuwS+AjLOWLOZvN6VG5Mut4p5LAZI71VwWvzFc7QuMdJzuJf03jmMN6LJq
Rd0zaW2BAalR73W4sm3LKXLb07Of53YAYv1+AVzq1WcOXQyExRoWn1SDR34TEvUHh8earL3PfZTN
2EPmpXHOT5p8iwbZJOEwsJmajW/FH5WQq3VCwxzBny3gIAqb41T9hyYuEakfs+/cptclwsubXAOT
f+udxUX/nl0Uxc+Kb2eEHJoJhCO3md87QRsezdJbK+JECE48d4YY62eE1gBrOLnfPiVvh/5WrBJm
pySV3COAvixyyLadejUtglCEFlGX4b10JJsGzma3usy2N7P0W3DTxf7Gimf+EyR5R6OVQ7JvWdZK
SP978pBT94SEHhMX5MVqJMASNJjJBX0Lo5Uwo2qcvIE8WtxvPgJl/9hhwBuuUBmOnoWEtJkKoR4p
WxYVt8tTWTDOCaI2XFCFK/GHft2gYUnWvQVgOFEyPFQM2jICPv25mhMxxyp7wW41wjzUfEx4yb91
lFiR/seWFsHOz9kDn373Y63G2+rC9IltYi52katk30rI8XPnSGwJBhawWkdqdU7B377/lm5wg7uu
KDptkXmLOjbiZII/OWXKbxO/VQG/4CC0VU6LCzQq8c2QErHPxAnXjTRltluaRSSPOelElfI4dWf8
hJOVDraVvLPNdJknYVJ3OsF9N3OqBUAH1ojML3TON5Uamjst+d+ikosqCqsl/PkoHVqCIOrUk0oZ
5DOsWoM8ctGPOkw0Ttx7AxgwH8yyX5p9N/vuuLjx5OmDoRgy+nq4XDdtg01X+voz33QVmcUO1/Yv
sRmfnFvn2jPRX71C5Xlcm6iMiiDm4cUEyEaJLm6Ck56DouOx0fYi0Hj1jdjKQFqeF72fONK1ot+W
iqfwPIZVUMti4vap+d0pY35Lz3bGuLvrD3iITh4yCrmjQLn6zYgvuQq/q2VA+cOInx11BvfOU+zw
XmYgB1ziEIkNXRvpVdVPjmAvgKRum2Cj2H5W8GfOFgYdIrfg7r8wNIrUDTYpOlOPwCc7vDGGKmtn
CpNyx6cDGJgLxnSdFuK3O1Qddw8lsKjfBzMuKXMm4dkrAOnwctrJ32tC/gZFLLkdYgXmdocgKURA
aH9B064+qbx6mv0pKRIfiQKiA78KUFh/xEMkW3ZiAtYgyswfLYifrZ6SQbnDsq6+/Fh1RCaqn/BI
eSotuAdhghjl9Au5uNwEmJxu7ZYG/Hy7SFk6bk0rVam+CrHssnoeYXkGMJUcKGRXhfNp7YpwO4kI
hovqKa9ibxtld7R32csmzDdm7FTYveFnVDiYvwJceMn3pimZ1sHUWOk8q/dxbIaZY68xa4+lBB/4
x2Kh6SHs4hrHMMvlNtTBNsa/oqskj7wIhsX/bOwLigfglRfc9XKYAenCwhBytOcEJiUQJ6gF5NIe
IF3hkqQLnmyXRnrMl9yXLYBfiyT8bw9AcQHqiyhsM2YhouHIdTeI4mAKpxrLjN8jE1LNDIJZS1+h
lXvC1Yv03cFIfv+lnf1gbbtP1zDy8It0QuESlEXpboXtTLQZe49DapubnP6SMwloCNDr1/md81cz
3nm9XFu1WhSySrNoJdYN/rAMkH4IbCL9TPNv/d047QSt84tb6AF4qN7T3+aJXrJvYP4zw5HSoolL
3sZ+Sf6cAvJ7TZ4/stG6DNvfYJmriF2uqrHaxbKoSMD/2ofjvgurVCKjszZkYNT5gi2pDE9jzBDZ
xB1UG4rqVS/PgYf53Ze//a5c/RwkXXazp97DlKAnlURY207wum3LOUvRSYM+TiR60vd9esOEExYq
+p3RtGSd4TdCR93sUtAaEfcqlsNNk8r258LvRSEVhAdheEEimjv/gNbLc41jHnaX2W8Pp3y41QD/
cTwQBcjzdOjr4DS7IlU9p+fN/jQ+DODDsWj3Uk8kZDRLBNoXs0JNqG8OtXUY9gVSG5k8sg3FmUF0
q9I8xV3pQYjzX1bv05f0S+2RdryKsiqSJtuQK9hj8knhsk0gkCnhb6FiO0nXDjFPaOdMkZjNGcs7
3+1DI+k7gQZshZVseGTT1xCht9esHxcmwoQQelDTUXPrRRpdkzO3hlSRWwPxQlmMjPhve5gFPV4e
SDVV/jsbqvo689z/8LpnZh7a+8z6HzB78T2WaElOYW2XbZSlnhGfhol5rsAPzfb9omQs06z1rY0G
Xw0BAZDY6DivGufyu34a3CHka5STAkVuLZYs3Be8AyQFF+PxTibavmDYKovSGfX9NXSJ5PGD8m7d
gWKOk5+9iVFwy6i9dECQQlm/H0tiXYBBGXnPmGGIqfY2oMFhOE4JjOPORPzEtKc/bMe5MkyKbxLa
VXIW4pizoXV/3BP4IuaF6WJ/3B2AWhyz3bhehwpUhdGxloEd/NNYBsVnOpWb8XT//AorD17XrZck
8uZ4jGIR6JtGTeAvANZE9KOJP/58+e3hlxFf8unNoBH9G/B9Q6yyrYIX4JJoia9pwW3gjihx8+Cx
uHKn7yVukXqYVDMbYnt6eJGNL9jdZYRA0BkKQG8Cr8IliJcr8pa4PmbVjvMQDJK4IHSHDkjTIr5C
52s0iJwxExgz7UmHwoPBonvvj3+24RKbXDH5MjUcn01IfP4vSpB7FiyMWBB30uZ5Pj9pXtZSDs2T
x6+2vOxtSgh/8xi7Ft7/9lmtuM9IMhQAQROpRkKEjPkvhtgYGTkT47a60AzKSRZShIoLiQvKruiA
ScYZSH9Ct1dWolGkQ6hM7kLEgNP0P57SdKJWAkcVBGIArvn5aNr+HPmpP11ePsaCqTI3ovgDfTig
IKjrQmjjuxi0ypLT2KQCpcFiK2mtaT2H25u6FU4M+HOXyGnIlb3Go3dOcA7YczjR+TEWWHy4NFL9
Epgoi5jd/y00bx5M/RdX8fD3TkOry1Q2iadrMttrLVqL8NtFMpNWQyR98EFXpnBvonvnrDEI+2n3
3x3ZcIl0RS29rfhQbgQvlel5vTLifnDq/szJkcje9NsFJDpjcv7kJZNVydMbCiVBJLr1tHG7d9Ch
T3W5lxJKwaWqAcUTlUifF/E77GoSP/qmZvSYeUawih0FlE/YhupqN/ztcxuZoMNJ14hX9zuxTAdz
J43Jsg697jEMRGQ4IdxJB/cNrjGAzSrCUZ8l97rO7+ngjqXWFWKirtqLdBoG1TxWcYgdqbgWrxgs
XUIsyNTevD9KnFVon2cqNbSEZPbBdN0AcomtbYVzOXTJ2a4hyQy5udSNajqMpkDCanDabaaioxWW
VXT+gGu6emR92/Vt39UUREUG0WsxMLIenAgGf4+lW+bNXzxShuM323wniq3BkW6zcw45Wtdsxtm9
nu0Vv5r5L0JDRg4wEgxBpkvEmFqynAYsXGBzYvfrm9c+RwaGhmM8MUDsvr+HVID92Bm5zSW/1EJa
xxJOJZ6M02WNxM5XD/DJ9NRQSV/Oqoj//kt6rou+cbcmlZCUUOgoRW6FfVWUyANckRdnRNDSVd0G
ETP0wJ6WYDttkN6IICaxh14FR0JAGdsZjz4DasCWZfL/03piNET0Utyjmx9Sgr8F2CwerPwydSDR
KPl2Neme+ssQg65TFe92jwApkx6Q9/BsYbU0n+KNzeu10vT24AcO1qfsuhU/lI/cHPuJVCYSfu+g
s+g02s3mBf1fZ4APDZfyH1NhX9d8iXIbwjmNjVsuSm6oSBd8p3f3AH9gtqZCgtJ2M4uCYLLh+6DT
u7lQBhjwDS3MsHjD1NuVaR2AWFUFuWbz6BhsrkngPfBKPyyycXWffD3vfvtPf0PSXAecP1QZiFE5
sIr33+gTjazHTOJ+cWTLV4U3BTEic/ZDXr6kDb4bUd+L25j/J3xfOjBEo4uYcqTos6xk2FT7QZ/M
oru3uTkmgAZebdpl8N7OfmyJ932e+WEdtFUJpSb43VdTQ1fHfsHpE7Xxo3HXMSUOGhti0fIHmB7n
uZOJgGY9pyf9zqqy+bnUACU12w7sUV7BkCHTAiMQ26Fq7lAqb6RpZ33XwzRvJeNMDzkHCOMJHiqa
83vMtPXHUhtmQuaklY/xsZ4yllEzBwmq/Aor8oGT4mPBqcb0mpRmBbZ8LfR7pTZvGkWcLNqisWpb
sUg7frcVHKfZkIrDh8//Eh1oN6CcXKInTkyNmaGsdgGo/4UW4y8sIu6j/IR8zYx35oC/P7JB01Mu
QNfMeS7Ti6RVp9CRRhSZdvUWFeSw9sgg7VlXnzVy1Sxddk92yiqJYK/Ed/kx0Ui1+3hFn0B2WlaY
fyD0SEAFIri1X/d+QK0/K1ltIyHci16SWBLBiLTkmGQjoSg/L1RGs3slktY18JMBReddczv6ePlu
04tfpi1vv+VLxhz+4Pz7j9KNU1IVOkr2uWDrhUCxCGahIOw8BnFv7VBS2S5QaCAYvAan6Pd97VPh
SY+gM4upCjQUo5zkGeJzFP1GP4o8XGEhyxgmARQBV5836Cj3sN2wqtTGR7CJF4vZJO9t8FR34lo3
mjMF7XUKYJMR2CxE1H4YwLx/0gAYZM2oEzuvhHdyECR8vkDVwKfDKCX4MDKxr3D4eKkpV9rsysZJ
B99WTM/dwPa2stm2N1XnaXTZbTLw5ou70WgbQKYP/+5omXqPyk0tr4uZSTuwf0vKjLS+oWCCDy2T
P6CWwCe9q92fhT8BrDrZDc0cGDnkmM2MeDTvAeIZKjf6J7/uU5OlF4LM16BP4j7wntraSP8DV/MN
WJx9JPUKMKGwiybB63okAfjldv/Us9PYLrHN54svqktQZ2ngrgj8xnaN2pyHx7ONYCZB+spizKJe
JEr8SxvkxhFyZT1fRaBWjNf+JI5+CpHmbmaiJggV6QqDYAbuL3G9B4HB+/h1weQvzYP8wm2Xxb6T
I5wfrqP8pUMe5twOvB2e0HfKYxOujZbiDyFpOfwbVKXb2pUFAjAY4gWFR2cbANP/UhYZltTB0XQL
+iRa28/A4zEoTNC2EmGgjx/4jGib/FgPUCqYUwzvvP27Oau+TPcLGDaT/QOZeZo7jlaZ3S1ItKwn
Xg6qoJvk1ztX2qv37YxmELxhYP813NSLnNHA1llNYMBrPvJ8sFL5q7+BH/0a8LnWFwzJC/h0a8j0
GVdRvkDN1vaLfo+oLTmfN4o2xv5OsxIN6QjT+seem6x5Mj0ZlwLRuCARUsBbDCJ899XJWYxhcFEN
/voT4bHKfUSnttcPQyjfY84UKc+KjzydwhscfBVxjBHOMNhaa1jwIFLTxS8QBiRqr36NDdr8Muor
W+Q4StFw2hXBRYPupi/AvPH3dI8wlQWrFGvplcfKiGNIJPRY0034QE+5b+AxpnHu1i64aFPCrjnF
ZA64sRHnbT4qaiIfBPG1mksx8yBhpK71eSr10IRi+GKqxPAeM70NlE39iMkmye8XOl4HU42tWMTm
nYmeTNpjKm3qxpZevENt6nLaJjD6E6wZZJXcYl9RGM+nMzgkQwiWJ0YiXwS+/qQ0vMs0Vur+iUBQ
MY5N93wahdtJehnCmVnft+19yNtr/CGqUzP+BJ2NGzvDPFN7ujj+M3wzlyHmj+NCAE5Zfb7m811G
aANWC5dxdzBtXZdyopjsCdeUbdhUvBsEHTC3IWorGB6VH2W0ye3bsxaKCwnO1r/18k/1+pZEnUNZ
0/KKz818PaAym7rD8dDQ7zdChlGUzxi39IYCkVrLgy/oyM1UJsdeul1UKijdqLQZVdPKUlTXLvcS
VfbWUeZBzVfB9kbjn6jbdf0fQO7ZafRDfSY71u4oZc4FBk5un7eyI3rTtFrWr2sMhFBS+rP1P56s
7c4R+iop3bSSAdlMj67n8R7huX4J+0kcTbpg5G7ySVB4VSIKJUKOEBab7pQWtEkCo4a4qJWg09oW
gWJDXUZGgr8xDZ7cvrqDul6ync8vVZ9sLEXWOfT1EQo0RJYsJpXE33/KVEdV/lbkmIcfKmCF4NCz
JZid01thFXwadSPdjlYhQxeaa2x0B2dWFnK7kApAOHt4BdeV7VtrSZP19GOIdl84QlthzGMDWff2
8sAD1iHDh3RgivJG+smJS6vlwJjQTHOIHwPAG08nA4MmS9PvLwG1hvafYT1+0D1dAPEP3FAevf0A
+5Isb5LhBqpMILI3/RkAff76dOE46lzEGvw6CqNLC/mY5yxuO63nK2SWoLSTMGFl5CcMXtS0qBwD
N0dPYZtwTHjcjJlb0TPa5SJ+IadBojRxqR9pbpghuiIQg71PBYnO2pH7eAp169CSX8Ef2vprClHO
vgFF0Lc3x/NATPtMQwmq+1Fo2/QRjKj9rWDX/Ox/WYJCCYprewoldMNBGevLlIPRLlkZ5lPIBKjc
Ru4gH/xflIdDbUP6phLJ08jxVb/ZDk11ocB3YHEUAse70mSLWXFMxR96kTGU2e778yqPh3X3rpzP
gNDbO4ITJIaJltJAwqOAa7gexKvBj6UHjNX7rmKS8BlZLwyG0lWU5UdXkYz9bXCQrWh9Eh+8nctS
kvmVjSPpjeLItlDUxhCtU/V6Td/9Rb0hyHP7KuDWS5Oumd58iECzIAO2XdlWwa9f2cRLi80ysy3S
6s3SsKRAclc/xVibAT8y3eE0PrAxscpn7/aOQ6nZfNxeMgnp9P5w5qhiKQb7u7raK7cgKf5oCKWL
Wbg/MqfXNjvRoQ2Y4O/Pu8ntpksE2zJ9iubBsD3/sWUZFfZWglSYTIE+kiVBdt8YzoC8RQZOYUP9
Vk3Cy01+yxhXLxZFFSSWJ5XaHgcD6HseQEl+SDrr73ei6H5SYkhuuXPwUY0SVqhjiPTtqJmiYKST
SHCKVAr4ywUfMHXzfvteGM25gCU5Vag6oc3zAwLbh5KWc02HTYNKdTaN2Z9Aj4hQ6h6wYF0IXA3/
2DzoQeoeneMVTpejf4g5J3fzXFDXMSx9A65qwQcNJ2FOvRDPmf3Yx4BJ7Mvo3KszVJvXDxG+yTto
CnMgogXLiqXqOakn5L49cZA3A9d/dCQip8eQ39Kdp6YCUbHuiKrx1unA1Q9Hiu2JcXQ6R4tviCeX
vrO/4Hl+NkMA23HjhCw8yIY5AweKOVfJbGNL3dMsmYeDY9GcV1Ogen6hwFjwcnq560HNnYE7qiNa
bXahl4pcYpvdTpdP0UMMp/jXo3RYwLrY8wiCiYW7fFgQtcc60bKh50prHTXQnrVX17bnEBVyljYt
8z5Hs6p+ZtsCcETNiEZ+QuvV67TiIe/R8mRK392gr9Tr8sOC8XZ0LQapmhqpjz1M0dgi+4I1ji0x
NolSk9TTcOtPOBjfexQ6qDh90up7ufvPjjagV/TGJ0dX/gxWiLCG1ha8RQz2wuTw9Mi+ZmTuT/ed
k9Ih8l4M80wvrw1TwEZeh5WTTjBE6nBr99ySeeX7tSnmOAyh2k7XBKyyx0y7DFoVL9zdz30dHJsC
xCFBrhkhyjNRMtSm98W8V0Jxjca3nX15NX1FsQxTlgxjMiYdI5VuAJcvEV8Nbu+olqfTkMad6ZB4
IOvdg8onB3s9FEllaTQjrkRjUVnHpcHErFp1h8C3Ttbe6ctKmNLU3muv6LbP1sd/pntoKmnFL0wc
Y5hMNTQlIK6hdWJ1Mj0d2lIIl/vMpZcTFePU23SoNKGhS1hxEYlnsnqibyRd1uFsllSHzR1VrTFh
h5DO5+toSa704PNannY+UGFXKV/LMjGKhvAPvCpxY+0ODwNwPNNnO1nuENrZIMOqd4Le58axdxCu
hSCAZVCcrrs+kLkXen+uGR6CjGy8VcZAQ1wQnN8xdZ45YlcPce7X4185w6NZEwsy67QR4CIs5tZ/
YwMkCMruAarXaxCGZvBzxYu2K6lihqwwbPy+S3XWk+RVV3n/s92//1Rv5zSoyPjqSC7GXKMTDabZ
RiXxlRA2goIFMwq/EGyjG1VN746wQIkQxGDqPNIk7FgRa3gb+mGHlV3m4jiIt8A1FnlvIEYrpEPo
Fx6jW8cc5bgvR8imzEBsEOghwx0agc+bTIx7ezveUnDDa/pe0cNfzBqVoGVPuo8ft3fJmw1boDEU
akdutAuTNaLa/uL0Gj+LaN1awXKrN0Mp73hEubAIUG8FT+mI8K9EHocsVKDraGKLYuNb/jt0oM1R
MO1C/8BYkLBi0hstfR1B0uQz8tnIssHWIhR5ytB79F2Ah+b1L+YcnhdAVKJEtDfihZDaGiRybH/U
bID8kMQlJ2GKJoLPCMkktuaDohqD1VWlC1AQFscMOpOsiJVywS6ULYHZ3uCIlx90bJC0Ak6lfEHt
1hq2oe37xVCa0i9ZGExzvdImSS9J/afi7WO2a42o1hVBocewnl9Ef9a/EM7G2IyhUcOoqQtgqFwu
4uZv4dMcggp5LH5uJzmtTOAn1ZFSIkZ7N7FPNjktgUB9SQ+QdGXqYvn0R3WI04RGLY5k+aVmTpud
ekIy+RMQIGUwpG8Ts70EqhKFiURKrFD0pTxv0VCKrqOgLFqhblyiWuCmKx0GQzOiipCnOB3/fB5e
G9Hj6zIhpC28S2vDeB30dDqVyUM4t4Jn+OE8E/xEeZmBc8ETPDVf0PEtu7DSSULhR/HUmF0MvhjG
GBo0t7rlT1WpWuO+7U9+DHOBxmvsuYYFqDk60l4nAquxn3Miei4RKqQt8eXxRAQ+p/f3VHuE7FpM
eaPrrkzDuH8OFwPzwHmCBdTvL752cNaRjQIEniAN3Q3bFi8homSz6TyDRG4SLhkTFU5XynU5EOzS
Iw2f2Pe96nWD6BNupXeUnu8DC/EJDG5U5NKZ50HcrPSBIO0Yq/W7p+d21tCpToKWmoug80IBNnPI
XQiiFD1VE0ZZH0BXkc5+ivjly2nq8iwSy5+I2SmlXCCNsya5+RSsOgHCso7nMUjjG50Chfjdkzfm
bXpbJ4NrvFu438eu9pyROGMptvhAQj77mYZRPzeMcNL2rsDnZVvsYtYY264GwWMlndYje4qIDsqr
KdGAwb+1iDfRGnOAAaSAsREBmzsbqujMcTbHEyNmsGYAlmzhczvF4CfvW3QA7Hb2mb5oizt+8tiD
lGT4v1nlEU+uHr2GmTcyMJvJ0dxQ//b0dmIy+wOu6ggAu16IwFh10M/O+wxBsTo2t9ujyFvQRwBQ
iKUI41CPX8nn7QiXT2JxaiYiFbIROP8y+osVk990DknchBWL8lFPTD1n5tRqeRGurUe4O9I78g3t
06qX970QvhgjCAL1VDDO3G7zgekbOhNAau/rW+6MzHKOqsDHV0/0rk/+GaSXbR1LTL3AkWYeGiBb
WaITwiJCDjroFLNseBrLqSLyz1oz4YwJOUeIdJSAA8Bs93vtJ+r6+v5DsFNqVE5fdtMhWUCgoO1y
rIbwGYQq7OzImx4DjcxQbDZaicGbpevqZ28NWYt3rHGeQ152d5/OsohDEq4WM944rxUXjj/2ReC0
MRdaMIjGvYBzw2h0KQZE9ZDrOO1Pko/sSUrLC/eDOPvI6YHQWF7ypQdHb0mNwyBzC5XkCGpavRr7
Xkq3GQ0NOZZ1YwT8Aly4iv2ALwtflb2bwVspgkFVfqDckjE9WFVqyrwDhvNZR3JIDdzVgjjXMPOK
35Ylx2fiFCV2+rXzANWdQOHNLBMTvI2nAZcydBC4RgjOYW25j7AxNh7TMgQUacY/8fPelrgA707R
QO1w4CugyGaUiL+g7crqaueGEskECDg2RBUr2NkmZGy8QRJc2LhDbNt13haOZCz0NMprRXyi7QRy
v49W7SL+0z+23gUVoHyqi8/BTs9B9mLFtEVmrJr4Dp1dI3ysrBB43HUjfwZ2LDJ4kPKCE64NFhMM
KHIKdZf/h+Zs8Zbwu43kZnkKa+dqErtdQy55EeS96Lt6JxNjnh65Hg/+3WnSumZNSWeQqK96UJ9I
BLPwVoscqOfPuDMzBx4TuCflNQsm3Qq8FVg3doSHsrFZ8QI3ClKv1DbQsIEXA1xsENrEWfQeD0/C
0rg8GY0/qfWrG2NN3nFA41S83hwAfDppHLUpsCRytXtD9xdmzbs3e1SDuj1VNHTeCGglfyX+oybx
4RzSA3099zlSs4j8jEDiSI2R0R1iH+d7LVMo3xZMYldpD+hr0i8CAX2EzNg4B79qckxUiOAvfmfn
Divs0Kj4fTYrLiGi+Cl279jLNxrOePvSu+O86pm5e9ukA5DfwG1qwhxHRx0yFK9aRC4miSecPgXT
LcFJyMqDKXILX2aRaLa9grP2ypYs22ZOGGOuUiXhLbHL16l6UdLugz/lXI6FvQ5ANHlW0HyZA4Ge
9pyXkmOgarjblbNAy5TSn60G34yXZSEk2emFiikCTa1fotlYS++mPGDVKWTh9bjJ3hWXZ8sFxxNV
GfyzWiZ3oSeCJDHAZ2RtMhrwMvMVIkXlj8zuF5g76n2HQWQvU7zEVwR/dhZQLrA2PgCvtUK3Oczh
g6CkH6Cu+jMz25TYMI5NqnbGTo3jfkxHc7bIod2REHQltUrniuGreAERQU0sF2VKL4SlgjndzG/5
sO7SjKBcrHpKPAu36n67nfx+3xJzgjUX1VD0Mx9umExCBZhNRUxvOPcp75xsaWlg3K2HRS8SVATB
zDgp7uX1ImVeLrVSjKfNAaaATHz+MHDe+JDRVN7LJvgxuo4IhTAB9urEMN3sUd63OEWEMdidn+dx
jDtxVoVAHlhr5Af2CLZ0s2XVCgoQnfQQmvB5rVoybBbgu2w/UqPuGTdPFX5T3/FMl6zeqGLSVeba
xi5BburmjSpI5YQosZUL38xADRdQF+eMV/2istTzMDHDUpMAdaoPNJsHYL97PFjDU+t/juQfTv4h
c7i8KSVH3DWcJRHitVRSAuF5uqwLvzepSRqVRpXLGR0YqzJMurRIs2EgN/gieyW8VH04uXyL3gvT
P31lD2jZULklDmgG56QbcUi2EMGzj1kmPLPTusOU562FDJmEkFPq+CFjs1EZRq+pEfTO3nCad+p7
nC/8nudYCNf55Jj4c9XWYwM2nZ+Yw0anh5m0nCe4yL+gGRd2mYkOgR2oqqBT+AbrNhqZSoRi8yjg
WAVMmR7lXeag/7OayT90S7V2Gs0Wz4krNLYa64P6noSDkQYtJW42LcuTg2rIF0p1QXbcThtMhiaa
fGgxnfhRWHnmSNRVUpyMxYtXhdTnAxLMIsdVN2dg/VejsOnmlL8t43P2Sebd2eHE0RmLVeATo790
7EJG8q4onJYKwhPXMq5+kTV5MmtU91p5u6Cqr9tBTklkyh+HCmSNvapLamG+wvtqX9+lz4LRYb75
UjSLmTG8czEvrbOAIFVYIilYLPWM+NzZbUOuCcxsKq+MJnhz8wYwcMUpsZy6RzDg7HcRaUgVnjOH
53GagbVMiLt120QceXYYn99xC0d5h41gBOuBZZP2eXEufcHnPVBcRT8ubfDGXzeWi3OZ6qe38xez
xFWAiDIOkHSE1BoZfjEP3tCTYSqsNA/AOYZyiW9YKYeowKdCE5BCnlogG0GbLJ7IKwtVmQ4QBqTs
SpVtepaj3qafhF5bC3SMnFfXIy8UeY31Wp3wm1fsJSCFKOPL2VQ3tbSt3vfFFDZZlcNiJzJ51BAW
kfplyGxOYrsSHHi0ooMsL5Q9n3XprWk/opg9UsGJMUYkuDVnA3FpZfWGKhAFeKbdG3NCtc4Ts/rH
4/I4JmVU/JSYf/+BMc0mKl+ogyosg94e08YTMjwQRfNqmxz2HGRhExc4cyZZz/TWdcQHbjoaGc6d
yy3rUsW4ZBrtjqp0AZOOgau42etaUrBO4933REbsCKL1P1asqTYq35MWmsM0SIv8UqHv39vhit0U
vPI86BCfk/R73Bkkbg5nFHWT2+LzyR9MXq9UTnHkq0+RnXACo8/MtfV/wSGuQQp+wzSpf+cM3BQn
EqW+dQByUd/+AFCfuXOtTMunhwZdasmJZs21Shlk8mqiVlhkxG0uTxAQrJOXU6YXOvcAVZzxW4DW
0+tMQY1ktlE+ba6rOn85HAkkfIv9fZjL+5ZL+uXm8UuxqI0VTO9s8AptHxGe7+/5DNU0J+PL4lkI
uJU/Pw49ypqb1DrsfWo52+Bk6lx/y6KWSYSqQ/vyOiCdp5FgiXF5Px05lvFJzjWJhSn9f3YjVMr8
aYThnFUDX/Y8xnpC7FazFOK/dtxDeFywauSMjrT/EQhU2XRZrdILRFa1YaVVUGBu1kp2LIBIQZL/
OWUr1svSxmJuZ+07iI+3AKtWOhvVkMkieB5iaH6694/FZOGkzLiuLp/3MNfOpduEbqTf/uzTx7sF
UTxQiaNSIdpSa2FEIQxlN+KXtYjlr5YVDuZjUo/fQTujKX1GKf+DniFp281+3b0NRsHiZVAgEvHA
eP/ZYzZcrYSwf9V/oRcEM/CX11dED7WH1a2azkpSQ4aIvZ4Gv5tcK9xzoAwnbBDde9vAHN8NF4yL
VH0E3OSsY8vKwSt4F0YdMNbryNzc4kWHqLzm6tO3O91I6dQxe4x01SyhKJXT2KWSsfx8FFYNYmfk
c4r58q2P+dhnbgDWzHJr9p4PMnJK2nSoUDfxZdRn0IwwuuG8X9wScHR9n5eYGuKbBVYsY2sLhH7s
fLORl9Vz9Z1f8RAR7iEHHtUEtZP7bG55P8zB3lAbrbuNZTNmEkXMy7lMN2YENsUoT7akeaVYO7Sz
hfG/4k1AI0A2298NhAWNJ1Y+DkHLRlDfJpaUomYfE0emuSHB9JRShKPxuccu+4uwNUNtKFbhtT62
Kknx0ccyfzhIMoo8xI4iupLDzakrVtLGO9LR6TBxtcI6oQlHJBsIFEnawaycyTbwWq747UUE/27y
TiuojRSCDG9BYK3kVfxEBt+YbLUsMjX38+ZvUvIjq+jsXJpnKnfHZ3K6x7PpCUMHVlwAUM5zFdHS
fc4a0cCbLQ5R6Mgzlfe1zvN7sVc9TKYN/Lz4tA2lPwM+46CKPa9AxxviPRKiLpfmUreO+akLo4ao
jwhUTygVnFVwjl7RwiRsw+oKUpV0Qu7g8ZeF6TY8GpXvgG4Oc1lmgAgdkatmNgMAHsX5Z56wKYep
XoDLSNHmGi0BAIhK51C1FEdvCqjxfGJwAEBMVKuAJNYDJ9eDgfnD9mwUookIxvm1hzb/hPAvOQN0
y5PxTB0OQ6PJJGk3Fd/V95cq5UX7rrpjZ9fR3cxPZRu5C5Olffr8M2gWcTga89FptBYTDRj8dvUv
4xlHnzz/F4L5dfKPEp8weP4dhkbLhxpixk5euKBw7Dr9gjbMUrOS3yJjeYBSlm9b84S8X9zgzayY
FEzwGzFukuDR3yQwdj7VB9thzFQtDAR5jKHF/5f3KmJ6mCnPjR5tm1seMwK4JhDkp6EI2xNLCCtG
HjMhDlpEJ5qyjZ30CTE58D8OfrYAeqy9N57WcrMxjuCW2oyvASRHQH+yqXoEM7ZgZzxk9DliGNbC
KhF5Z/xks91xgIdIhrfds+FA1WSwAENOQORja+uIVdkVh31CNY26AoGN1TiQsdYlEiGjXQ0JaRYn
mB8GTgew4A3xNeCINxBljCXYCmrXjut8HOR+E9hu7aaR1x9sSP9hAMOUJ6E7hkuQjC9V4aj5JGJk
QvuHpMewz3vGwVR2Lk90xoDLkfDkxcusORkS5tSv389sb9S56yH07gLbNbPOCnyELVlODbxNW9UQ
FtKo2SS3mN8jYSPSOP2dXvM98m0u0xTBD6i8Lgc7YswA126ZdOOviICA0Yg1QInPdsOnEbwyari4
WNbX2ssNEbrCIA9hq1Tu6NfCEyAkruv3pPqfua9tbDRRNYooKOddJgZ12P0CWOB5j7JCULXY/udx
LTJiHGhPs8/Z8oJ4GGu8rYth1WZvuv8O6/bJ8klidL6bgDKZEYa1sKaUykQI4YSdcwQrp8d8vNZr
MNMntWr28Pim0459B0aCgw3eY1XM0h/RhxEc3ZQ6d5Qg7KBk0K5u7q9cyUI/XJcKsitKDbTjk3ni
dFZJo4o3Tp9XwymIvjOOPujmiMkQmMCXUb6QaWC40A4Jq+mfshQGb9nUYzswSxHDwohoL274PMOi
CSYZNyVI/4Ex0VRTlEmuMU56d313QB+fPqTsblZJk54SytxwmBLWcoYoZFQEJ4SSypoKGyGrwo6o
gzYZd1xbpNLtmg33zSOWBfqjNHXNr0ym1o11anpMG+Um89bC7M4golt7F7l8riiv5xpBv2civ8Wi
L4y9p5R6VESquNJWQcwrqLgrK4fXHumFz+BPLRObZuhMbBBnYktSE6FC4LyKdZEq5Rh88j4krf/6
Jve8D2YlFEstkbBJ+2pR0uXRPxkDxCYgQg2MLi6/q7wjogxuqt/c2Yqd0ZmW8qe77rCsltnn18CM
MKWCmkmTS0JPrBeGMOaVeKVtwZKzwm6fvAglbKUXmBAzXLiuYYw3mlxksZugmYt/KkYM2Gxz9ccx
fv1yVdEGzcXsKCeDFYAohKn6TzNlmqdGIglps6c03VUAgdc+7oDaDZV0gm77irhiJ0YNRzfL1oIr
59DxdKqVwlghyDa+1JiQMnUxK9XK921Z8nRtmKs0vvrvYMZdhUt0noz3RAukY8IEolADiZ4SGwh6
cudSlVJ7uzvwj4I5w8M8CtEc3rfTm3NGmLv+XvPgQELJdeeIjDd+2r+A7/Y8wJq92slSnDHR9tl1
BHQGYM+UbhVVhSG3/Me67/MrH1wSZ1W2+qN+PtRYgMLObYUJIltzQi329XWDawQdiEpYsAy/cMVB
fSmtBIQPLz6QMO5D/7fLw7kiLml66rRg5RAfRHkdFrsM0uJ+jK0dQki9HGy3lwODZZdcEfM4zPdd
W5fCgrOJaHnMr/WIqJad3lICmomOEWaGPCJSsrfZEgrC+k6gOhOC26uHKoQjm6a+Uk/3iFG2kaPk
EfEsCRbCXF33xMWD02eI89Bo9kyyVW2Qkr7oXII3xzlfHDoegkMXEP2avzbBQ+WUYJ6hVbLOAwgc
xx8VNaU2WKtftsGe62XO31NsdM/IJNPN/abrbRmGVfUlZ1vGDDo2O8bX7XWp53uUO0t+uE8VSxla
P5cYtYHaQDL5xKR/FDfr1lbz7n5LJfHQWouI0Vc5xNECBeax0dx0zhpDkgnJKxInOWeQqHMvgvCu
/al3Ea3YvGmVW7rzwGtgd+N6Ua99NaogJ8e8wn5FlVMH48bVAQQ38oyB8BAQpK6+YyhbLJHJyBlX
hhnYEYMlCG0fDpl2hGkM+Td6ynq2ZJx1gNsHuqhNsilcZMFGeiqP5o8kTnAHYgaooHpbK2m9lGoT
rbVQmi3uSkEkJoj95hPMIFJ5Nvi7RV+211Kr7DnVUEVz4q7h7nH/pjTJ16QVIzjYMGyl3prLZLLP
9y6fo/v3tO1zjpwshgfTouPmQKmjzOZn5+jgagoUpPGCDrtxBEgsaNkp5MlNtmFpJ5B5luTcF1Gq
xXN8gHMB7DcE8mPRnj680Y2ks3ic8OHpzSeil15p2rhShhVvgL2wlYjKLYBv4G6/PeYyKVSK5eVd
onDZio0v9j9BmnpQwAJANk8AQLHOFql7dRSotJnZYyKyzSzefwmsEO+f5LsYcrkr+v53DWcUVAQG
Y9iMYiaw+gL6ymFIH3210od1/cqCp/dZ8Yf98dekQf+zLqC2krCTegzjCalhE2IhHfVKepbD2FD6
vTbYsaEnTbJbpKojM0M0MfQSa1OJ9CztTmsImCoD34efRSvexD9jGUcf6iDqbMwukmwOMGLj8zyr
+g6Vaby+PVfzuDf/h8Z3ONyS2rq6/MKifHZYkqxr6A9gxyYnpfI7kH3tCPMlV8Qmu7FW1ifkhHNF
sDYL8Za+/84SCX+7+w0AWa17a5xCM2ghQ+n/VhjtqmAlljfMVBAwE9IA/qJQdold+Ffct/hFhkdb
4kZkBfxVGNQ5vbXGa2gd3gHCo4SYH+xCWo3jytQTHCMJuu4oz73E5+oGmuUUcqmNNBN5wh2L6KnJ
FfTtteq5/YkdtiIRaADJgZkTklIdCNZDr/KcXw9jtIeV81qTFSiPrUUZrSe9cgqAcBOLU+HTnykP
rOYFaDwpKAxJd7SsqS/gidcwZmt6llcGoA+L1bWbiV935Q8vYKoA+EU/hrTmDwXopSt6y8Nn88+Z
Rev+PJsDIOm+Zhq6z+KkUKq8azjfPnYvZpQZqH1MF5yPtUBZbeqeWIMHO4++B6jqikiNLZrOfENn
YY8lUFv6M4pxZgecdor3+HucBvmmGowTc+HNNsfICcypVYAwsgrkwFkFoAUPFYJunW9aK7WitCJ0
kEZqMOQ4kEf1EEOGrgl8UfpPnPnFLLspwoFuh0HnLLKlyJWZ0/38sV2vKCz8NMXTe+Ii1k8THSMw
H94t7pbg5hUx5I+wGl2emES7PzXynSyBG3dlWm/nes8isVmXtQVyJSFPDlg8kOGr82ifVKj6xbvr
7fAJcd8EY+xRHrv47qmFv3jV+Z7tD76ms0R6KguJ0qs12BkhCtTPnknbNeCjECPh1HQqgvap95f6
QzGjMoQP385NLrC8OXV0+IQl5qQHNXseTklfcmNXAeUSRyQCZhfbvnt75No8NuBekoOLodz6YGDF
dcyGHnhw/YE/iRenVrB9ALNGLv6sIncja3JLpw3YrLKVdFdcGTMrQMJBwWWTgYOQsUUNurqQBj5Y
aY7EZgFCn25PuX2wrIsvcBcim0adRaI6xCHyLq0PIq0ZBjPszXvUdr/V7ekqSYNuJTnkhiynR84u
97c386blR0V6VUcqBkHtxC4h38XJD5oQ5jtxq1YPIsiSIQl3EJ059Xb7Rbafw1ehLdrOs7+fyZ43
s5LVE7NnrzSWcF2JrqJMe92cO7cLlFm0nGGXZ62kyQU0i6+PwNkML4qFUMeaLt8NPq+yCNOZ7JUC
DbOvnqauzF5cGcm8r9moDmvbUgx1N8qJjHqUztwK7EHU1fIVd4FHYYuEkTGqaP7B1mMS0rPKtjx5
e4ft1rq2u+YqXtXq6PC1Qmk5KhRBzsS3oLZo45TjToFH74Ggdna7qDNarvsJ+HayuyZi+Wb2jZ/n
I78yQ1d8y6RGldY7TdpgR/MHIC7OTZnUF8FtPi39GJHsJSTDC/FIpOHaMpJi6vUi4GTCSklFCsXN
h1exxmmSyhneIfLUT8IQ70vASa3btd63xpiKXmPPCE/3ru3WnmxFx8SgrHmN1bqLw+NXrdmsq02Y
bhCkueeiOaqnbasV4YJGh/UQ5/7D0F49+Qn0lhtgBl0IihoSkeqCDIufshhSMcMv/r+tzrSndDkE
1wt/T0zqVBVkg/iH4Q8wGfzAnAwn8tWL3qkee3I/UsCt+zp4QpysMnChT7oWsRWRUscxnNCgO4Xg
CLWMfG6mEkwGzM6HXqs8v9JgXq8CDppwph1QQJoRErIZXz0Gj+NqIc8yzQ+q9PZYOx2n8KQrnN1i
vwTC/Xhn/uh0MaCpTiQ/gGZIFwPOJrnr4dCTkikMPmv3U9/IZEyy+TyP3hTfQh71DGhHsOzrRF42
irxqQLQkn/gtfBnq8zjwKDFWmJZosh5oZf4URETL+SnnY9gsHG8pty9WsUz7zMBOgqtWamJrXmDP
ZVllgw2Ye/Abnrynvqut+rkUHxYhoIrBx8X9Wd90NEEeU3oGxhStsAKhtCAltkKXzcsR7Oss+CAk
0hacIc08/M0WD+ABC+xKIzsA8Sl+D7hWqzs17JDMlsyRHN9r9G81blFpoBdcb/EZFjTdIGOOHcJV
4w3vM4z0bNzgQhuX+658EfCHT/tk04EcM8p1So5z91W09xJayNsiJaiAjPk0LYqZP/tkMPQPdc6K
l4qPa0MkcwVJFIh1y4j0cFO4FXDXSh4Ujy9IMPM5xh/yyG+HLbqToiCgP36mQaZpa6DrZzUWNelK
QjdFKy/iLI5rNnE/jm8lDHDEwNnhTh0Lv/la3WooHQr+UFoJxkrHwcVlf4FjvCZMCmqqyKpY74Zs
xDmzl4gBV9VlHh0aA1AwRNto75fNwaSc2dCA1DJ/L+SsUfDOGpLZrEwGeaJVTAzbxzzEBDbtgjbg
AuC7fpRCwlX7sAvQ4ciWCYkrFcHs5cpCRnZ0tfhCOT0iPESBEzLyp/taK8l+4DoKOqMRsvPqKUMp
ABC9cb6T1gSywj3inYfDWJITU/SQj9zM/38rbFVu4wz34rjMpnUyUHvmNkFdthEavtNYDTc5Pbma
eufwxOgF0XBU/BfnO1MnBZgFBuvAT9Txj9b5FN/Kpnqo2JE1a1CuVy9qncBcS0oSsbX4BFvPNjzg
2PJKpidhfagrirX18LO/hwxodN406sBELGIS+Q6qcJVxCrNzK5smaFdG9+dqamK8pIKSnSK59JJ2
XHlWQiPsF6EeeN2g113OsNYF3go8EUpW5qzLyVxQXOwwucUL62rQHFTAHC9UWDlpDCBUwA9YVxDv
KPfVVW6PeCcuSrEcJ6dcK9Uvy7sJIefJgYDmPC6WqRF6SRVwq0sbuqd+6ACVdYARtqYevtPisZh9
mBfZvXwmewDDAfmjm0rieKnSu3+kP+8sG7Ivo83lwn26HREaVhVJ9TsIrKSP+pHFAC7xVr2+oCYY
e9M9R+riYN1JDOxA/Vne3A3iBa3eUA54YHXD41wDXCacsqpThZLXA/5rEGwqKTPBh7KxMipGzdeu
o20K/R0KnicumkO2Q5jzEcssOH4hiY0KXE17PRz6W4iIMvNHJKHBIsH3LGW99FS6I0STzrGk/zO8
+MwKoSwBSJmonOwldCRIH5kVvegd+vBB/COx8ht85XR8mcomosOjIcRwAcZvKYf9AI+VsuGrslNE
48O5YdYjrxZPSvesiUTgQz41r59x5N5V39s4pEaD01dTmF9MunG0G/IxLyelXwPhaNA/f1JYEZpK
6gD2sRG+XB7M2ohP6fMPglyt7+2mc+nAtS2jdlEbFF6sdf9HlpgLwEl0hUjc5nSo6AGkHCUUQ+FJ
b42in6ESeL/YysjvrW+clKVuV3lutn8mQJ/iHgK3eUG2EKCtIoYZaHK54eod2Rv0P1i8TnhLl74p
2b3a5oB9D9cLWTLdfIfyf42lHjOrvUf9XNHOKG/kjbSOjxQUNG7eMmezQZmyquyUrpbX+6B3oZbz
Q7Y4iSCu0pMMIwHWr4ONsW0YwpuJwnhNfgH8GZdQuhT1tVxJNhYydkXXHUcKdn9T/pR7bzdNe/Gf
jUxG2QaQbUalStcnyDeTik5Uh59LJJg6DNAhQLbf4ARDpxLg7RDji1nSX0Wlhj560MNJbvfwSDEg
3soT5lY+ExEoyJOjAjUpJUVkmte13B06Vqmm//PZfxTUZ791c4zJ1fVftMzvoIWiooyLq08amcCr
Gx9A5QW2oY1kKL3gZlEdkihjw9PJ/XDBSEoY9Vf/Bv+BDGlFujC9konHxqIpnj77efkdjnzyi9ET
Zpwpc9qfuZLoipPL7vGuL6MzUObC/bKEzCFzKfdJ7F4TFv7G0vs8A0ta9EoGgJKqoCcuYUTTkkD/
M75WuoaFXtsD8yC9vLrGHLo/SGIAtI/pB/BlTBOJM1YqeSFrKQ+fup5FShx3iwH3hmKdFVHwD4me
uZchn5kWHOn87K2RSr1Pm+VR9ZuExovHZSb5KuVSaczYwxH2FaqTQuUhchw9C9KFvQTuEsXpq+h9
rFkTlnM/tb2tS4MkVMVc7wgQYoYh7rtVfAdDbyWuZv66XrAMbG+JLRV0NTKRlAomD6Tf3uUmTryn
b15M54oU/u3yMCvpQ4goVDemWF2X33vzYafQ9z8BxF35qnsRk4QS99x7pM8KyVGRNA0YG448a8w2
WWLqJB+oPkbd5wvHvQ/SCqvQoCHJWLLGYiHeioztFgxzF4AhIuRGHdndJaJ9z8SE3vDFc2HDH1ml
FXFvrGD4nnUcpFDOK3HweqhDuee37+dizW3MJLWTnEd5msxv9Oa8rfFpnQ4NeB8sJZEBdjD5YmED
T/W8Q9gvNeE69Axv8GWvQHkYfWlqspPKXZI7WSvB4C50HQ5PY6A5PBXXdKFhn2QPPemH1qvXr678
kvv6vMlw5DkoWhv+K7j3oFF1ahez+4D3ly0l8L23tbf7Hl2L7xCt1qEc16w5Ak7zKTL6c3ROlSqB
is183Q2J9Bob1lycG83yNTuzi3JEydwZ2GKZmZ5gp7DUE+pM3EWWAJxvxOpSTu9QuzWfYscBS6er
N95HojjYVTJBw0BRAtQTWOeK4tbuk3L6cEmOTeXQHn1i/xmpyQdwQZaY+/sT3ArDtkbkeAgtXi8w
RCNtg0EzQPIqG4evVRZmq0sgMGBAS3nuru3n7lMdjpWQhl2IyZDyGfI1BLykcxm0GCaRzBzlFNre
QE9oBT6DBsxRC+w6o+rQtEASE+PgFw4uKoH469LtLs013gRt9Hz4OyEkW7ZSu/qyvF/GEJfEO2np
q5Hr/28MHahLICmQzpDMPPSDUfkZLDmAYKPHdnq+3dZjoll0nw/Th1Q/SuOvTamZqf9jrpYON0Ld
ueqanWfPs2mnSXBW0WNaHYL9PkxHyn4XTCQ2KXQ9nDTr5LgEB6tRLs7luhue91TRlgZdkVaDieGy
xY64VtFDZEz9KIMrF88xsgPXPlasp6/KWIdcHKCTCQ9GdluyvMXmPvEhp8dnMBTINiTS0zdMHvsm
pZOdM5O8ouR/iBU0p98jQry+haYIQuFmlf+ZvNEn5R4QAWoSRGW1QGaGIQuDjDfa/nzjazpt0LqG
n8pIrIKamPPdnwAyzR+TJOFpML1zb+WLGsZPO2x9u/wSKu56n8Xe84U3owizgZiELQqsJK+Nd1lb
sjxkawBq9vRNSpl6v3UV1M0YXagNYoKWZ84qvwoKn+LlsEjT+R0NHHAEHxNWfs8ccsvsx2O21fsh
44IK1iCRsNE02hIst/rL7s2Qw7uMqPSP5aNuK7LWjShOqTfZvtEgLguZcbYeF8ohworV+/YA2xwp
mFwRw9y/60Fh5nh8CyiJ4pHY+9GQ+U88NlB5vBVvTjiBkrcWAAFCu+2QJiGVaITOxHwNnfo5xs3S
OC6Bmlb5Mvho70cbgAdhu04F4mXUOgV0ShUjbI1enas3dexlfLC6b3Co7uyY+lcmdTSpY7ui2wQD
aolxNGv7/meiUGBvyMAXximeGelA+dvOCD9z2+iTRdSfRzTmSOAgbUXDyg8nybPoa605QIPpSfAl
ynI111/idyu9aOrgZcvFdg+Wxg4C5F+TBJcNeBzr11BfjWe4i8y2cAB9c/70Cx4/B5wpQZ9XJJj6
CubQ4t0zMvVolgfJAsPN4lgrxkIiSbpEOSBLeRpzITTSJ6N7W20m78SCf/krkm6Tvol3zS3jKQ2z
7kCSMmwVkk/S/+rBBhh5Lkz9lzbhPS6xShl/rGllXl5/Kn9QOeZ8uv0q/qZW5ImOnUBzAZEqGTik
7OWdn7r3Bjbx3IDaN+25iIB44NX7RatcGC7K54aovFwlxMC6vnxO26paLDwnMp7+nLRZ0muFX6mz
Cjq8wIDziWrIoLfaNvmMot0640Vt2ij7Uz+0Q8ALLODkeOIZuTOeu4trIAF/zD/JDmpJE9Pam5WH
sfHWw6LPSClBWhFkl8sGk/CeYUYBeQvGyJa5rTC+UaSS/rFzyYzQT87BJonxoKCVV9VGz8KOIwMQ
9H1lZNx1SedAo35nsfQq8AcYQeglLOxcxdqHesehsRDZfko7jE4kB25brVEODcvh0kZe1cS01OmU
2ZS15sk2qwMYh9pt4bZ3leB0Q1wXgtwO+EetdXM7j60/YXtap9KQ3KxVtdgsLr8f1i7GMFRnp4Bo
Yf0cA1CUtNXQJd0uY8a1bQfSElWr++cwhAv8n9msoX1WC4KH+awF010xt/gfctDHiUyHSFZ/a679
lPnFU8H7/kkFmvOfYFTKs4MfkeYFxnmKfkvBbKARuldCQL+8ysueBNi4kOztp4V+66aLv1TBunZf
WTFrNaQ/64Wm8GvyeHSK8TF8/DzvbmdDUkDPo0vAXF0y92YsfiEKcvi1iOLdA5WJnMnUx+Y4qNg8
KVDgBT81ueHfets+di0GjjwUVuyQFtrVYEXotqgbRkc0/Pmo14SVfXHAyH17OXw86sh2Dy0SEsve
n2t+Wj6jwyMyXUvCJ5hMOmeb+adpq8aCZnvwFXNRkL7pYySzKvIjoNueVMp09W2a2eZ0fOob5kZD
iDoBhFJN8bi2U2ZTWSWAhlDuhQZhZAZpTrujTMMNp2DbUHqk0HpKrQTv80X1QPdQxiqs20XaAJCS
R94fCjhvxOKINZPsy2M6kVyKT/TEPFfn3OJX7+G+3ZlxLIZiE+V9HE7+7Ym1NnrXQljcgIYf6p/5
bUL/kLAvOSJQU3QT4oSjU4nCXVvXOsvBARk3cpU6SZKgP1wf4uTf/+EeKtu1gBxs0voAMcnJkJzj
eO9U8/q72UY4Ta/b5I+PExQcqovCYGuqL7B8I0zWF2zxgqoGexjGlwRTBzt4qEE/xiGDqHiTsr3n
GfahUrwICfMlCdk+c6S9safQiH+58ll19ULpfNOCJjHwNmZnLs4D6EaD0jDA37Us6hQs4fQolUXd
0MTQlkNzUS4TyzbgwMfj6Xp7eImEKxit6GIQuOtCit6ERGEFEh5Sft2T2+URMSHzFAQ50c8EkQr7
kU+L577a4x0Gi51RG3F2rvWoBYLutI7xzsWESPF3yLCgNTIB8KUSF8PD+n6DvJWDn8c3PJi1aNRv
JoTSaffRGedhA16pGhKt6DCDUt4CMsLwUUGOLji9t4FwK7fNQHgAWeIYHnaBEjRpbKXFg5tqUqIP
69YWYpj1rHjiixs3fZ1aA+JI5fChLtN/M0of8DRZKjhIo6Ftc0/DGTGHnIThEdY24M1veLHLqwlI
gEy2xOvLaYUEbRpdIT61wMoR5ZyCEeiUD+px+ZIiUvLvDqCUPk2r/CksTauQqvaH4xxeWMOhtePb
9Te9KqzksRPoSY6d4c2aGcitFpfMb5vkkKyHF7fYOiQRUYty1PikAJl15/VSOAQEO0a+vFSeX113
GTSe9BQLA+nuhvOmXzkALQBPcyb4IVrdf3ljUIRxMOeZhGrikEGYsvxfSp55OObMxIKC+wOkQxEh
vNwWqbv+pblQGGQdEJMVweQaA6sW2SGeldaqIS0Ie55I017I5leIuQ+sHtoCKg/lf+0G/oPAREWD
lbGfgM+p4rRgHwWdUM0Y508Mtxsq0Bg1wwOi8MP3LdHm4J/IPjgUFDrL9MzKZtnUAgA99hFhFgm0
bCgPMOkBNImAgc91ogU5k4pwIJFDdzINrHIswTUi+o90wAjji3Xv11BJ6/q8MTjuMpUoELC4G7qC
ilo6VdZvQ1iD2dOLpJPYZm+J30CT1vCzKjJKWNRHOPTbY6Z+5w0kcVdit1y2NSi84JiO4qv2/XyZ
3HLyXqSRgMP4GKrpoe9h4dlbTDUniOYkaBcEHIYgX5/6zjmUuodWy/d1vUvNrpsuB81AsUgHTmDi
0eJ+SewFfLrLcjCbsXFbnpSxpfgIhuma2of9uzLRVOGQdjLfeqDGPrgevs1HMhH0vXU8xdWUQafR
lcja2Ps+KJOsak/eDyalyacrPkRJlkfnHeIEepaJ9j2DOA04+oxYSBf7reMi4gdpZev/26zsDV3l
T0BQ0XXUIK2uwdUXmxurk1Qn9a4A7xwt/dYfYyV7BGatY6Ef5NTJ2JRN+Eg364wPb2orvqxvSCb8
BYxyTLha5hkIkNnE+p4qBtGnVGrrYadzr7w9h9UVxpAJNtYNiaPl1d2zx9cfV+rrRyifFsnImM+P
SZpdlWKQY9hgs0kEj749bfICFlKfbTbrxcb8yVOsCNUSAyUodHTrNI+40opam/cMJG9x2DCp4CIs
z7jIyxu2h5Zx+miP6SkQxi5P2FZzENf5TzkIen4Ph3JVgO4vOVbkMzJMeMDsloNxNzWA9yYcxpql
FhOca0FfmjL7ewV55CBgSOwXNRsF0SeGlBacwjOFImcN1DfzUskZWzWz8VrQB4cDEFMNkUL8MpYN
vy6Qu46R40mlp/stXrvNfl9t47hzel02rtONQ3XvyYH6eAGM44KS/XutNXqSGqeVWmQi12P1Qb+K
TbTVx5v04TghvoZAiKIubXySYbgGlHE9LIJTq7HNrW/WMCN6Km8kX4G+L1LZ1Sl/LXPkwqaxKNRM
DH9tMxL4iqbovsV/6OqFuHNd5LmQRZ7VJbYW6jn/dsOA09bSjC9OdCutocBrOVGqlJlr9Mc/P9A/
6asm3YZOLWmFO4WGHttzb+EpowxfP5W013rPBcjJbSJuAioG0k10UXvQUI2l4eg3Ih/RMvrqQvfo
fq0HEa4bk3sXiXUorlvbNjjfgkbthixjSJ6I6v7thwGYhmv3XRpr8dxRQY4sDnR2lrrV9mA0W2+h
m5e1hCqo/H67qKOtmdqTxao9o+hnOhlB7jEAAT18lvOhnATU/qvtMzVKiX3Arwm9f3nRDv3Omw0X
YZ7V7jcJMNCG8jn+7yYcfh6az/gRgzQiRixT33PT3No0QwN6y7o91PwbpABRTZXQ4uMTpDcD73+W
7NqZtcjtmf8zNu0VdfPNgnYMPIVoUB+QbAGDQQ/RaJohseQ7GqUvtcCL95BN5oxXR9uYMjOXT8hx
hEAxaJbUWvlpPy3uP4Vbj0juY9tAgga8Iz5Mgqg+GO57kIPwPM9FQFhN4ilL8lS1Du7V571c+Yah
grQlWB9ejDzvGV20i/Q/Ly5c+l5BwUL12DF7zhcPCKhrxQtFhIGer+Z6Zue6B8Su2OyFFWB+S8gq
+AO/mkPHiXWhc1cDgx1jQRVK26YbzUoJ7NQe4swSyqcQZVqrn67xpbn4X8G7X6kSJCXQcmM3g6X0
x6NatnLgg9jSZ0D0qRTUOJYRRvXKYFI3hXlh7LxuMI3uDmWr+8C7tUMIm+FQdylt1ZHW/lERapTn
2MqKPGHt0I1LUV503bd5/mcn9pZlV6o4Tf2dv4pS9nITVqETI3+wj2mD4zWstiBlEHzWtbuW1k9o
ER9TUdgVoCXR/vud1iCvs5rzJTyLdPH7MA4HTToGe2GgQaiLC4j4HtunCoDjZZ/6DZm9j2iQh9B+
wfl+JZikkwbFO5lY7XoYJARJq0MG1v8nIoYpwBFUVG1vRLD0gBo1v4I4bse5R4pyV7meqO9h3WAe
4qR61LUpcZ8nnTxHM3CnJf1WreEhCENrgKu5NikxbKfv7Rqe+Z7rrUqlTD5FyHjlgkiBCjKH3fsN
Bda58mcj4qNkZg0G4EZaxZRpz0ii/JQWVl2b/2Yk9UniUNjB7e+q8yVGqb4+eLebPOn3Y/+sLclb
enbIYX4FP7vBVBF0LHAba4a57Fv7p80Ky30uaFti+yidyU6pxZm/NEcF0Q5SQxo/NSQfCXuDcWNp
k8ZePSMgbhPIxwGv79e526t9AIL7yuEfH1EzZ7zsuiI2qOvf9xxMrR87aV4rbX6chRZ/DWBUVvYw
37+773IlKpLcAgPOqKfQ7pu2pBPiMduBNT+qlNX3qKI9LZf7OrPgKeY1ySYD8ioOB5pimwX6qo3g
wcnDhAEzka7OVhBdD/dsG8iqQjeasp1PRQdK5XSoCTyROL3FVAJOf5mGpTZ36G+uwsSupxQF4UbH
MVoGYuuPkYbRScIdNbUio+Y4bL+o6cEwpSUvM7vh/A0Lv/g0Q+iZDQfafq/L1+m0m+tRaUJGiMy2
57UOShP9wdq9uDXW5YZKd9FwtRQJWSzCIacWnRf+AkAmcUutZcCmTyv0PpP+KC41WuFMYZ2LiJWg
JRa2u2fk4hPa/mMrySiXJfukj0U4HS+pxp2hP0HQ6KaIo++Fn87hh5axs2QztV+AgS+OQ/a3X+OX
PBMbVXptaqviTPomH4MmiLs6mRZvWnnuZ12itoitcO2MWHbTrkiRXqgu9pB5Xtkpp862smpHAbP8
NX82rI9cHpzWxLHa5UPYdcek7ZzqHVwVJa8ZyuwWaYDKjnuITD4pzNLlmgRzxtk4vlljDRmWS0NX
tFKvL1YCdg1SLHVy+8wHqf1NxdBcS/9Bf5O/dWZvKmEJ5V5R9a3/thb8LJnl983FNPoc+froc5YE
JXiw860V9hjwvH3jy3nSsZU8yPI2ysy1OjvGv4KVBpx+xG4P3o7vjgMO6Eof+zKxPyNwsqL9LHBV
e6h/JUIYEu9Jl29nGNNEcj3u5F6XmMCIuP4VT8cdiE/CEVqRI7Tvm1KFR0BYZxuAwCU909wy8LnB
N108fS9whmzr31IZ203kWsCjv7dSs28T6qkwzjFmYBhZXch420fyRYH1/Wj2hvgATTegcKwYtiOp
R/4FIH3o82JE81stE8/o4Edcnp63PATyh+HDsES9P6PY4VEwVYALIz/CPAfK2+L5oeXssWMVp0tu
3x1TuTCN5TzcGzP35NX9skwsFC22G+xG+qREC6bUSktVPyrO04ma+Pt5DCWRtImu/lqaq+WuAU97
bAU5+oT4Sw6JZKvh0XEDeP9HIvlJXhDf9KTZ6qZOooJKpAPNgwGGmB+YZy2+Sqt+uqJPWeLFHrHI
4h8l7pCvwHUnWwm6CE0tuzCKXT8phuWUQdE9Jyg+UN5Mhcu0j20B8/nlm7VjF1L7KB6MiXWwNWfM
8SkTd4o/JbqhZ1sM5ESAqdLKofdvvN6Wp9qBFbhb5EAg8P+n/w2EqcjWFBM3Q+WG8gW9fkCe9Odt
jenqqvHztPr+77U0SY4qtg/bOavEuiwNsMq77kobUHmwUtJdN0PSgzLpPqaV+w9b5QN4JFA2bjK9
1qXXs2tJs3lSbiIQnh6AVyoH0hcuzl7lrmT0RL1CuDTg/BeFiqneCuOBmoYnL4Gvhwax+zXzuqnJ
lMV5gjj5Hu27dkZK46eg1hR1Vmapo1zIOEGHb7teHs2ZuzaNpl5/wQ2RXOd5abyfNdizKOshdJ8o
Or1Jn+IFpNSGlv7w0Vh+Q6HT+fK9llXEFvCsZp0bqrKo4kLCaaDL0CSUbwvNjj34iB3TQjeCPi1l
DszZ8Pnx2Us0sXlENfOUJ4WlXLczUjKhkAhAA5AVZYQCtuZkZRpVRzso314/0rDoxnOnndEPKi3B
SrE/2BJIUj3tqnPaD/+5P1+Rbu86KEV40vtGdzZ9eB5OzzpCI35+K3LvDNFbSJ1yoMIk6h0CSqKz
VSAF4YEsaS/txwRpmC8NCIW3P5NUjMf4PgbDbMsfHxFM1PdCX/fhLndm/Y7zqEo/yXfCI8CZz8/7
5Al2GWZcJb5UVlR+Eu1c65Z3GT5P3T1RJmqhuThA4P65eB7HdDWFLi/x5exkfuknrkAkDkfIU9bA
smtdiW0q88UCl7TuQ7H77jCSf5yEPmY8NyfRnTihgtj/i/fx9el7QnVYfJtQkGKmbA6xUmC7k1Vn
GN6R0F0pM8vmrA021iCDshI1h98gn7W5czCSGF0G+XQO+QUHvi7vGngqd/j7loCf3dakHHuZueG2
UDivyu8sx7VwOfg9AG5D+FeuQprcdd8VmLHJs+oERjundM7nUS5rQCGFJY2Cj8bdKOOGSWScLPS4
E/rXdHcgLBsKc/uHLyfk0NsqsBMM4R0Ymax+cQmZxAAa1KRhbHTKLMKMTxxHSeN8UCcpX2lzrT/9
fk9sdBaExk8ct9ndVlcr3FeWvF+YuDXPiebqllDW9y8HvuIjkQAeQAqsDrZA6bm3rTxKJmsXUwS/
QMXSKncESIxpIuF78gzMs0S0I1Yy6YR/FfpqqoZny54ciUbv6tcoC4xdPcFKiBjPXxTxB60Kw6z9
LkW883BrfhKqDhzszlsV385FOJhG2gQ9yrYAEB+W1w6KLt/i2sgY54PCHNqkcOkfn9BmCWM84bwv
4Dy7V/ooi4qUAOtURj06RK8/hc3YBJGK+l8RAoJfr2QpkuiXLr+DYpySI5z5O0uB62HpzHFp4AsB
+HZTA8falhotAyHUl2qj6qYw240nRL5n+mUN/nCajXju0tu7ikzXeI4+36R7r+clwzu/09dB0Hd8
cCL493DzAAU4tz9ZHNfuVyn/gPBicfc6TuUodYzRxTm8iuUUNy63rwe1dEamEMT0N3p0GVVXCrMR
LLOF1yCeiLXEwuWaSs4J7PmI6Uwggo64EDzEqrAsduChOdqSXMJJ7/PirplHtvZO0/4MaE+uwVmV
0a+H1oDJ0qDwC2I5M2oBJYvpvzaYkGkHShtRDzP/glU6PxfCRYpic4hqmwJlKlp6hNK7S0LGQKLf
q6LW7gkuGLV/tUDgveBJ/uAor/trf4oy+9qWrIoHHGtBVnfxxj4Yf+pnQLfe0oun6ubr+2VtUVcM
xY0/7ktrSDPi9zIQlhmIGC46kJOOh2HLxdLKuy42Rffv4J0l/ysd8GaOuYrDxRlB5yVzqGDQdiLD
Dzzvp23/IdiTz82LriliWRlSTfQP4TWm+9W7OmzTmJppOJKZ9HRWTwt8LzXOIzJOvHaqHYRVu6vS
PY8m7Q2b+wLTZwdDYEOM+4lo/AKEZ1QxBnJzc+imOOTcQCfmmjGNa6ss/TnxuJknOVYtfLN6kDoz
VTKX6oBPGQSefRwaRXNsg//7kEmadcgBZfHwvUPNWx0D78ncRqOQlWnHeQD6WTFsS9lWgOrps/hN
NrW1tuN5d7MQDzMUFC2L2A3kYzC8YrRBCBRkuGREnWeYF2NqVTpLQyAoW4AMP3CRZSLQvYCSmgJA
pLVqxagiXoL8t8dQSMXdH1DnFCq/13WztnZHypODF83eGQLxxi6bfM3xUF3m8iRB7+oCi0pRcVct
vtqAKDXfqi31WTE6/2oKy1Fu35rTofCJ7NOJt18SaclNYveLpCYVdjl50x/bDbeuMgR7qMsi34La
02P47PgL9wXantg2vtNrusRYtOARti2LK6eeG2+IIa2AtsR1sJfOmEGsBRG9Mr52S+yFm8EOCWRp
J2q6YBgrscUTRb5OP6bz3JkKTG+KZtBm6KT9L1HiEAKlDf/ndF7jG3IKla6QK690R/mBVFFqTXtz
OBmiF9A+aRsCaOlHhalI8kygRjZH/Pt38g9UA4BQQRJSwbJeW+D8CySG47tXgKFhuWd3ic9fMVu5
omFs/VanySFUCxrneKdJr2yc8e8yOMzRK+Ry9G7qpVWLJvtlC3H8YR98Bpn3/YFbMJ6vzpJyWXxI
VDky/dWhKSo22+REFh0a/fuFpRVzMzBS8ubuXZQ2Z9UZYKs6jFk/PP1oJCEI66iIm4sa5M1hCqYR
q7SCv6Q4Y1Jd2ifplcQRPfz+fIHw3sQKVcPhz57jlSlEtgn2J8BklO3q4co/cEMuayqpJnMrcZ1J
BA4m/WJZj4cEHqLJamRqxtQqE6RxXuD9dDsy7VDwLxfxFZ+Ag0W1YLMgrWSefgDKN/68cGpjz8he
3S/tPXcQDl0KQcF47gm1eJyTQX3YJFbnR9OK0sBVUzkL4rsUsCOIcl1v7DejZx9anHDyG4M6M8iW
e80b9N0d/2aoT8+flVAFzBrdRZ0dNKIWZK8MwXHhgrLbbd8hywnn7fLO6+5s+qrewyvRzzh+DCiw
0M+5dgDPquNlryVO7DwgrVUgSF42XWTn0PJbgNxybWob/IKR5UVwoob7BqbPFNxxPKj0lq/sZSnz
SLQcwESXcMG/tADFhgIT2fRmIzswePzGVNWtw9HNzxULX6JPu3VeicIpCsgDYOu7Buzo/EMik+6+
nA3LNpsVnMGVtyR1AXFpO3X6g0U/LCCadI6wuaLg8RvYoQiFNolLAFKKYzfsSdTZ2bee9pxE7SBM
ElrhcmFfv+vjmNhgUcLst4Cbv/Ds6OmGwYqa7CcdxtsXgKPIVUv+AZrIa8OFQUo2XDiEOMbNFu6M
Jsu8J3ymQYRD3mW21Rs0R6DZ/1d/+M4Gp0TFx6RZrUkeoVruTyjq8FT9YgwFEiRZlZhErl9CxFW8
Hkf7QNGcG+QU68MpDdSnR8LC+e1P6eRORJSS4BVRKhEIs/Ka90tFicnNOpMJfXVjB+5VOthxZh25
dkbJASd4q9bXS0hrwt1Kf+IwDmERSDbj5g920SVE55kC7KmwQiwrXmLDBCGL3hZE8rskeyhl+iIZ
1ZPDHk4N75e0cxg3YKvu8fShKdYDfrO2w9biYzMbE8kHfd3W65IFYA2jH7rEb1ilc1lph9elF41d
wqqBMEcTLa3xDCxKrYKqcL7C6KWKxN7FUMT4776RVK8prJtoJ197COZ9ij4RzVyUODwj0lprqyx3
WzLf5oX1Bjxh5DgwqWLavkS46FN9M3C325st8leU3NPmYi7LEmKlkNDDu6jlGlZg+WV8dI4cXuJb
vPwfpD3gbrJmHdCfQzomR/f8a3br+W/k8W1ufAkNfmgQlL66BUSM3RT81f5kb4YKcpK5VaBU2aT3
I2IwtpK7whHQqLAYtoWObm2JrusdH4bt1+ei7kaVSWOHBGp9sjFb0R5P2O8PblVnxzIrznmznwQ9
tY1TiZ3kZC44YSHnNZj3gCkp/YGaE5J/MzJBfqo3P7ODxtujlHx0LLsq5cxkn2ZD4/LtKSzOfCR2
+NCUuQyEEM7iSU9V06AUZiyv3yuRtQKdr0PaiivYOsNo9KvcxznDqMmTFog3tt8GOxHa55PD2I7Z
9tBBePIAnv7FIkB+XWNSSqIAdvJCSL3EuKhIbdmO1VHhN0Av3mTVVRyPRhTrwJpPM0YDSttSv6qF
3jLT3SFvcs0hd3qEr1VLBfkAvFZFtTwRbCn56fm1X9jJCnH8Bt7UcPT2pOdaNdGW5RL40H9iGINb
5Mt57ivX5DzGGpl9Quk36hIYqbDi4p9GlkNIa80rfO+VfCyLMfcYNI8T+p7wX9EEcIAPq4Ry8k0Y
eTgSZeM385t+WAuot9NxmvNTVlrqwhRZLU2xiIRVQF3FZkrOHMkv1BFPM5TpbG0q1oLr2aR2OTSq
WdAHcD0cJI2IEYjw0t9igxKqFO6ZUpw5r7Ba2O6Wj8W03wURo5qj+yXgOHHzfDfCiZCD97Gy45Qz
SgGH4TBIXQakI5b2gX7F4rw96/buDWJ0Kl9nNU7Xca1rQvFf/pUHUwbmmDDI0Qc8sjuVUKFlgZRH
au9LKMLqIi8hw/dAqfEu4C0ZfWGqBtPDxh+ENRVFdtPWcemKEyei1D+HRrnqL7V9ZjXLTaThi6iA
8rWbS8Z8Sl5D7VF9c1AYmW2xd1fdCGs0bx0Ue+Nx0UMiXAFGwsdDbAb0hb7G1XLNCJ5g1nL9pMRc
r++Fq7b24tZaeZkRYE83x1AUiaeug3uSbXWYhpuNLoLLCOrQ0pZbLe7DiT49N9uEZR0K4XHJcNgS
JjJuAlTbWHjCiWQxNQopz9JT54HJiHlWdyldVWbzGkPxsDP2Ma5SHtEjIxpPoq3y3J7PU6xGzohq
0+Wd5qmYyd4rBjdBwLarbqZV/QsmwHk5cA6EOC5boMgWCs5FWYWzRXvi94T8wOMF5144eIkf4bzH
JiJEIenSxdh4v0TyGMAZ9IjjIVMWDsO0aYPziP29PgsLKeggkAzZJJEAO1EHBbutznNjrRD4ZEAk
cBHFZu8CD2DIgtji+dG4mBpQd15/l2jAgyHNrpHghgbEc1ekytBH4F8ozAjSlBtMzk83vp9/u77V
zVkIg0BAy+8/nW9kR25qgR1pE4r+LviKtUzbwTDVLiQWvCDjaEhJyRHrEDPpYoO+f1igYQvoXazA
e7SOHm7mboNvkHZ+n5doMaFkHa5tazAC03qz538UZQIAmhSLg5k0oc4AQhcNPKZvkNh0394WxU9c
jXXTNTTOPwOSg97sEBM8MKacNZIW0UP0Bkjo8RLuFnvX9ohE2sq9fWg6OCZF3YVP95AZ6HJMuV6b
WVhr+dSQkmsrt56TO9t9/YXBedVW8rjfUYcIpQ95pNNbZLbQHGeCmQnYRzxbBU0UOIC5R6hHyIEf
r+RorCdmsujd8xQZb1V+EWS9hBwbqnJub2Ym/gUC/tSwp0bAmMb9g+diTZCQrl+Vn4q7mS5YmM8u
SVOAvCMMe1aOLyCFn2RSbV5EjmsnDNUZ9sQ7lgTpnnJzd2oXTgp5k3VcoCdRlM+nKf4SLIM3gMUi
3WDbK4NJ7h7769F8csycaxYVPtTl6rhtDq5Xu3uSXu5UrD2miUqz2QwRVjPBzfrklsnVPLd2jGih
Sc1ZQqfJWwQwSNFHazqI3074PWRd1byW0I49cHMI5Dz7S7TrcoHAy4SLA4NBv+xReiwisauSE3Po
xluCBXmfgBme0qH2bQn7qyvcV11KTcUb5lh+8uRpE7binLUpFTgr447Sg1Y1KpDiUDxmTXP5egLm
3+nsjTz8whIjuHbPNH8xDk823nfIon4yxGOsy1SbK9rOeF/ZKRvrwhAxTLDWQCf/Ogcx3SAHS0qm
qbCEGVN3wRQKOcXLQ6P1fdj51MsJR0D4VZKrxgyjuxS6ptfuZk6CFyts8gVYWcJ/J50AY7dlcZ0N
y5QWMO/72v/hU/jWRtCU2ttmwzu/2FB4yZwLK20srihBfscvL8FOUNyFmefP80H6QbghUY/oZQj5
Ig3BMIMU9vXPieWr04B2mXBNOebuV6tnx6baQ935C4bNe9tNfxRTiWdiZgrtq/rv8GHifCpsv4kN
RwMjR5SthAPTch8gxjT+Z3nH5ND0aHeepW5lzspTdWsGyJohIHorPaD6XqMjwxqvhDTIhJQJGw9g
IOCtCasFBasrXHyWxJA/ucXZQvALqKt6mlsNBgXU8JSUUrZX/a8si86RiFrwPZzG9DK+9H8SSeIi
H3WyQqeCKzfhBNO7SigWS2ea5evvF4z/XRw5/yjgYTSKXkE3sOeplWaGMdLI/s3Vu8pPzwN3rvCB
hScgU24QqdQvlHbKTt7DmYSdFO8EAHC8leeC2J3JqSyIYowj1Em8UtCJeHunqQ6ZzyIl2rI+zuDn
O3UYfJIR79mvoL6L3Y0qsFDlHmgyqb5Q88o10zh66s6m5yf18k1hCtB/sVRXVkACskiMqfKUCihk
sYe7grNk9ukb8EyWFDp52BKcC7XSdPvQKMCmq561//4ST/OHq67I/Qrl/sa1uAwaVUassJcEZDtA
c0imPq/n5nA4cTQUJJtSLwiQQaYNPI5r0Bl6s9e7TNnfdvBBlJuUyvxy2zhI/DGWATZGZJY4WI2s
jAnHqov9xd1XhI+Ryg9dNFgX5XoEfrB0j3uxGrcMuQ1Zg8y8ZNJ1mVK6VWfzaa60YoFb8KQbHapc
Asit2Fqv9I/a0PlostA5Cb6OPR9eX/XeqcG1k9eXJpV09smZyH63X86GlKfNPDXQXISHhFTOeHc2
6xU8BIrmQMjRVrE0+dYpnY2Fe3JpW5rIPHp9UO1EUiYiMhHtvAwz7IEpyS3Rz6VPeCQRiPsP5LCa
xmtWJt7qEeJE8ibovrKDtknfDbfw+sM1IIpClPX0fYctQ3GmpleURIdvMYQ7uQB454uydjRgUFAG
9TEES3yi0UbzfSRQA8hr9/FQz2GuGvO/fShDPGUZmiuaA3Tcl+SN7pTzhqOGuUwQtMIuKumEV05m
crz81qB5jQSTVoqgpKjznpEDyqtSMSGTZJK4gilOGJgLkFvZThA7X5i4s3ulbcsIZ0OUttTroam2
JhkKq3SPXgDLb/k/eRbOFGTEsy6nZ1KIHUe7KbgC9y53wwxAR3jRFNy5FxtIbZge19XQEudnsApT
4Hj4ZgP9Lwv20UZFAw+tyOI/W8OosPOojhqHD7QccLf1J1JpznDjnIUn0ghf5uP4o962J3AZZseS
CuKJPa+pHPUY1t3ccdV/HtNKpj9gosypCs59NJoTHVKxTugb5pcGkOvwM71eE6q/Z976of1RL/Nr
H340mVaqz83f/bFwto9m0UUDbQPFzqmcqT2aSq7cLolj7ltWEC5r1FOl5KZaMQ/Hh96esv7YzPNZ
M58MMVFGKgFQ+At1nFV5Zz2pr0dGoRJCekpebmET6Rn5mUvN53kESFYqDXlCfRZl2QeBG/HHUqkk
Ye2j7FHh8w1++U4S4a5wolHPr/YgDe5De3WLrVgFf5CuNj00C3Bm/U5PQUbhHcOEIyz+KpDB/mV8
zEstFGMdzNgHKYu/lUqzXiF7YZGoSZPnF9bX3BEVsvsZpsk8YK2MJroVxncqZCniwsTQDY+Uxf9o
+IrbR1WcKuWwRWBvJsvDv3V3DucIZjHp8INHMVUArzbX8SohVXxFp5McfnIM1X33WtsOf5RE9YWo
Qg9pNQgvsTQN14/1k7mpi/oXfT6Wdp/+5BjD3K0KUww1bOifzHWDGLNKwYbxD+e6WHaRhvu88ABp
kEt1t33nM3tmnIUoGwdBDas5fWzeaHGNmYELAn6YM5jq5EWZfJPeW9/+OTXBHzbfL83/xicRpT8+
G1URUJATblPnNrMsdkv/QP+7f5OtU+2otbABiCH86PbUKvPUYQjtm+w+HLhngxTyY6PKdkfZaeyw
Ej7zvXgonqxLz1HgTPN/3odn2BEHjq4zXa538dkAHA7jubczMiFJ+cD8vicAQ6n5EI4DPh6frBaa
IGwXxiIBgaep6Hxya6T20luWJBTNGLICr3K+rTiOW32tJdc7zV7jAME+v1K/qAjlu8M7/34yFXBK
FSj5uJ24TzGYDHi9JRC8RhihAHJ3Hn5WFbg4bhXQfplCdwNmFwZnjSpBQVfv/Hfo2By1JU7mu1JR
TuZj0/PsR+Q/T4t6+uCrnaENwwnpqaaKln8tAf8kvZlVnAC8tEVaHYIr277XDJ+DsDcT3qvL16Rl
mJZHhhf25EM/Rr+EF1Agmgn8bPnuS9kduc2hNxMenvfasa3vouNWvPbR69I8/fK2GBm6ZM7PtdNo
dlvsAtTTd/JbCu6yDRBlS3rP65B1PUsKzFitnmwjCy2WV2cpJLxS6CP93Ryu6IMq3qQvN28rRSk5
oQUVACtYRfFIj8OL/jJ8y6GfUnc98vkuU5xQuadd9/38j322Z66G5+AO6Iy1AAo+micQh/mFwIGi
xqGGBndsR2/OQGdBWT0q6gw1qDVmNygc7A68sciTyypZjNIoiZriUjO/C1NwS4hEnxc3q4uKfJLD
OGibAVgzxEgC+eh4aiSNvgKCbQKUrBucm/o/Nk0PHBtucd24XKluhvThvf5uQyZ615SiOCIVEnas
O39wmKUb89PIvuV4sRCjpgIArEFEud5HL+Z+7EQmApymzR8yENpqRAb3jcEqgQr2gedJz4CVxjLM
KYQcj2o3ZnviijMgYIiP2Z7M+J6/oLva6GYjDB/KzB9tEfPjaIHB+ZnZ3BxV0HPGbXx8tdqv/Prt
ep2yu51FvufATnT5cdI+kSYy+wgq3n6vc7T45u/57Xk5GnCsDJEPca5Nvg57Su5l4+j7L/BEEO72
rUEVni9jtZ838cfr9Pot8bOgonv2VU75v2SEBId3gNjgEntbL4NxqvE0HBQe+jYtM1HMKmd3Apok
4ZFVgfcyrjLFzJK1Jab33UvOM9PiICQXt3ZYDYNnygVHf7TpG9OxDiDDrdb1oycFvD7IIUKf1lof
hhkwDPrc+C+ExUtyJyWjeFKn9ncbe3vXQXR7eIyhuqB2WXSk8TGU4DfobzIiCtq3kU8wHe8C3QGo
oh6LVriTJu1+GpJMoTRZS10hPHSOYrj1D6cUItrPBRlg+B2nFrrfjJoD6fK9pElTEES3OIa0wTA0
jpqe9t+DtEU9Mgfgja4AjqhZxjkOS0WsWWcZCSTcIu6DShh+Hrl2muc+ELV+u3ySxEfCH3N+3pVV
PvmT+xkblDQkd4ChDpLAbHvllDc9i9KDl+zvsINcAUIkE6RnxYKKp17TpPeiNGcTLEy1L5BQ/Yyr
bESXvsRX8LzM8lpwshrC76/yw0yo/+y20UGcU/+2DbfIJrKopxpEg9skdUl2v7A4/uxm+/mek/Jm
sZEMIHi72GZWdlu+ec6YZvl5oLIp+8hqNMMvmFRTygHiLzz2Qyymjd7lPodx1xEhnspROZc3Bt0K
tLl6AtN678Im4HF+Rqho+b70hsyKKbgkqgmgDCUEbiGo7sI1rYZ5rIBXV4kbzATnoqb1U+l6FNPf
/Is14EMYUL5qhIT9Nz7d/wcOoa/c+CV5zsUmyfgrBbc+pEysSuGDNOZZK0F97CA1mjt08J7G6AVG
AY5lqBhke+afEeGWVxajJKF6POQnGz3lMvdTb/CTzNdoKmVDBr85YIZb9b07aVrrf0RNEPqObgeN
B9F1Lwr4L9vk+uBCo3xhLmowTcPPeVJV4lf0eJp7P8WxlLl7fuTYC9Cou2aPrQIbZSVsV4HR997b
s9qalO3qGRbsVYW4WXg3OZngiVbEb6fsVBws8XuqEip0EW4alkHtSikInt4DM8G5Tc9g51xiBD/h
v3s50gho6Kzcli49zfqvmKx0Vt4gZpyFuk4AE1TTSRO6fRR5tjEjLGbuOKJDYAxP2NBtJPUJ84qQ
RSLJIgn9qRtt3DuzOnzwuGgeVndvACZNDkXF1Js5iDXLgxkveWblBmoPMxOwQkqKe077nRn/q/t0
yUIHTgtbzLU9pRg4fq4W1VfcVy4G4+rCtCyB5I9QMBCap2oAyJjdcYUX92tQGbL1GrkE+krGpnBt
zkzPzB3O4mmbCb+AQflR3r0HEu1trow4nGhknLAUqwcrqVvh5UZVqy7d9RPdOqztC6y0LuOdCCL2
/BGsb1L8pcM6bxO48nQV5itKjVNN3G3iHq/kT3jTfLk4A+vOAUyIUGPvMDnGLvKtCJFA21MZ4R0e
VkGvmYIr+AfkRVUKM2hb5beO7hLSd+sBEjCOrG3D4qi4kxtKAQe1X1cIpim+cvG5kaYaHK/9aDMV
jM75vfRsVrwZYKmnmVcrmwBoV+IG942CKqdclexpxD6Czp3ub/in4cFfIsUI6THeCmXud8nnORqT
SbIJy9x+u82I2viz19vx4oT2Y+q+vaOWGZ+42ToCH+2029DWyv3TBEq6nHpMF8zeuFEHAvm1Q/hx
GQ6HkU0t4h5kDToEg5kErVjsNt+juxXsJUWPYEQ2+Hr6iNcfPTvaByWvgc6nD0OxcAKnQ92Uq6r/
YdYLjQjmOlWdVs1Fd5/TW51PZjgDxzWl9x+ox5AxQgWniSJ8Y4kLQ6w0ivqKqy61TCwZpKo33rHx
ZuWieoTkz4LF0LUQdwpJg2v4En9LoN3tGardprakdKOSXrIRMZs564TmO8PPrh4Obtsp/QqfeqEp
yWfI1qldkmZIFfO9dEfzIDwPfxE3qEJhVs3W563jufsh+IURC1G8vO4JgaP1voHVCbSIXh/deMly
m/oCIvpns6u0oZ51+zJBr7BiPkfxkYqNmIrg8unQRBdelb1JFlwYId71k3OLas8HGHOkf/R9PzQk
Zq5UkJrRnoryQ89sYv8ND1raSE3aI6sCuef6wRnOhsSUng+XHRkzLmgW6EE3V/s7zOCP9YSZSQ4v
Vo55hRfOqHRJjKPjUVyQ+kKhK1e5H/pDTSyHXPpahmXt3//ov/3Mr6HKfEQxA/XFZ7Dg8tep/9Lr
1Mc6xnyd9i9GVw7SP94loPPkYvp1EHNZWTHWH5azkFiAqXNwg6FWong3RIlSjiiWgzVY+61NzR6r
jX7UQJPBrOCNM4OYvgr+uMxExyBY7SS2+fcd8WhwpYRAgdqfAwXC9WvNIvzqAauX+vBZ5I1FXyU6
cJZXVAYSd8PrX1X8LMIN610r2dJw/ALqhQSbG9XQJoNcKQh0y4ThxE9gbPM0l1SaNcE3U0PSfhdS
ZaCxCn+xRDMKvUJp6O0zvp84/3adV26qOYVTOo/+HreHRVCZt3D9eSIH/wuWsobEUuZy99Wk6kr+
o0Oh5HMhpYFK2Mt824jieH3q5uzMICiFWsgNiCQ4jtpjcJSLRB3DoKirsbq5XBmMr5PBR4LD5PT0
evOEeJkGqa1QIG1F1nBz24tuJPhcw6O6kU7oIz8+eJxMuNxAIVR9j8uId6uwCvFPuO57tmJnZuT3
SxkoPm0npTRBTLJLAIf4O1SRVDy9AQaiHZw7LjjUqeqcpSPUCbvXm2xibGiCiA7FDj56NELpe7zB
Dpb5IFVa4w4opUatvM4XT3Kzh8nPndX0mQyEcBvETYlh8cVpWjBBTE7eMsImMG4D67pNuWi5ZXA/
JrnfHDxbXjSl6RiOrfBpy43nO1XEjTChCIoeEb7iAsGJ2Yp0Tv1+Wwx6mXvvsj7jya0HUwFuHc7K
NWbPPIUmmPvDc5OcGWZOVnJJfbSpjYm8FF8xSTY4t2JTsuKYhDO6c61X+nkl5F8lKtRs94WpzlDX
6Md44Z8b2gH5paTj5z9+5ptZlLow525WxtM3sJQ81NnT4GVigj4aq6yza5ZhOgw+IKQW4uGWAuy1
n9mH0EhuSgoPy0/nkQppPZ75Ca90dpuL7+CO3P0fJB6X7q9KpiwOX3PxzkT8jH0RWoMDgdTqDncz
ULKB5QXev1JmxJZKrAyHJM6gW4yKwOrmFA1a7KcNVp3FVAbPHz4w/QXH9pq53tJS7KSM4t4YqlgI
VAXXcubbWSNeDQ2wlUT1u+xjpciTtN8fPHQoQ7NuAjiQayZaZUMhoPAWpL9Oc+3TGsl3haIk7DqC
UBsvVlnDxd2DhM4tP6BRbZKf8AhUP7KMufjDnrs4BXVnerp3CiijasY9Nq2iqkFzUPlBjnEZm6Nc
5qIgPSTKLhCgvf+1WcqJdcjqv5QUZDfX1nJy9fwvoFWLrbKbTciOWbnYF2NaFXx8x9uH8RhB3K0X
z/97+Yimh9FzrHOKMDc+841rbjC26c7bxh3xWG0KCOlOlQi0w7L24bg0l3QcPY0YXxtyNu+Zj1nl
GSpOtlEqy6kDEpsrQYF3NOmT2j+T1Tg92ij00iqzW68ErfrmfVaVDeQuKBYFgxZFzt4xL/w18BIk
EiQLtDOZ8ySg7SjrbV69YpEe+8a5XeI9K1EHjOEa01S0AkuoPITzO3srQiQTtPKiTSFKuwkPUId8
5mBCG7tB/pQGH+ZN7+vYO2SeB6wB1l+Khae2T8A4NmLM1WLgMlKJLu1BnXrAbfvynaxOMMIv9OoA
1HpqXKilC6JD96QLoPTNQoBpV7do9hPYZlS/gB6lYFy6YOwgOxGoREtLFmxxKzNvLgicRE7zCU1D
S5ibfMKnVQD5ZpD8VLv6F+RYcdyeARBVc7Z8ck7j14kRm/aPD95IDwKAh3T1lj3PGDNNGqDcqqSl
1idUXkXmTD7GZmS44UgHuKgp/KvH5MEhLXhEkhsPupVYpgnUFUyMNxXG/2dwv6VvGDZUxlNOz2gj
X+p+Zs/HivmnvJyO4X4S65qRp1im+8wiaw/saodTkjY2KEk0lterd593hwauA4RUVoNYIb/KS5iY
sHG7Ravox0zTNVFjhZAA68BCiv/kkK62XTVbp+pV6xJrcHOdnqGrmU01Lod1XsYR21dhMyFCW3Gv
c+R9Uv0tm7VBmzXFH2rwrdCrdXhigKogECqZEUa+bjSkTqO7Uh45aNFtmztuEa0M8RVTjhErtXIZ
wm/V/NgZtbw/+Ge92e33LFfQkpA8LthrnUmTDp9TClQr+pS4x1ru5wT41p3eP1HYeUawCW6453iO
AVfTSr3vXuVPaYNkaNhrBmOd4gU3430/YHeLRVDYIiSqva7E+oSM0xOhowbb7baXqSzZYJyzKizr
6baJXAxo1+23rZ2GhBK7fICbgB8wJSPUf+CJWJRjoVwpF1eZxhFlIebRoKl0RmKGPQGqzadA2UBH
nrSmqAbAnGTR29GRe5HxglMmEZOhud5awBZeqDEWRr2eFpFGq87rt1EkmZWsWs3RaagNC/JTzrca
1aM9PsBc+Jq1O2Za6JDMmZvwtC8+g8VCdT9/lrWv6ebtqc+boVyTnvo9NmDIbV8CLTmBwobbFLNJ
cct5phS0VjIAsM1ZKRS6nqe061ur/WwmTxeuHHOBswIZx6zTUo1RuWI65+pvYMGM3Ekat4Sfumuv
Ad/NSS9Hkbcl+mqcCi32M6r6APbnf6+bnoJktGuzVkG7sxHbwtxfh15Riw3LI+XWpPbIXcm1Svs1
QVWXgMcdMYr7FWD2vThcCJXe8ZVeTbzd2pRQBkChRqYzDDcc0hUdhyJuWiwMAkWrfki1y25sV9c7
645KJ374i1Tj5nekO0Kd7Oo+aPOD0FpxVRFWqrVAFFyXqaNjpfmn2qaka6clDi/cmUcx5MClWpyz
mFh7a0EcbX1JgO2qR/ERF3QqfNi3DOE3zUGy68Edv9f7wjlCq3jln7LgByIkhugYEgYsNM0I6IaC
vaYooKdws4cwho4U+kI4fAMR4y18kZK7JnfZMwaHLRwpBG3lKFbyshUiRslsZ88SyfKESrd3dmq9
8LohUy6bMXfUHi52YlBeACeu3ttTqPWHPYh9yWy/Ioi57K+oA3s793WOjYX1gakx3VCK8wpuxzif
yl50GxN713alOawpRdgqkDzqXrqrshbRxCE1kcVMXPjylw4Lu9oTU003ZlgV91ajQyreuB9pmYF6
2ynVaawSvxCUaw6MxJU/A2qc80wGcnDUvrmMW9vRxlEq/WED4Lxz3+N55FRdlKVXDqbxTHhGHAhP
fDLgTLWl1sVr4RPa9Vt3H5krp+9BoHT8L7kX9B6zaU/GYePnhJzrd8ryE2GH3auFDM/cCIyFxzmC
rwJOX172Xh9p1VzFOBRv/YnJO0rp+PmvBh00iULLx6GsXVtMvpiTA0ly5Qul3nNBEdGdcggdYFCa
or+QZx4iOJRPZJ1dq3wmgXDAHpSSxSHTWe1+qf4Kbv5t1kdql5g0hK/5sQWuD+C+zFskNndu47K2
EPDOg5IAcblEid0PHoJFSD5+Gwmzhp5Q3mpA/oiI11g6rOFlRaQ0GpUxj+3gSauseaF8wjmqLmPe
JSRtr9JYre57MUii18KoMv2Rl0DU1HM516SaAcu9YmMLzj+SNEEdfYff7vU3zbndtb2soNFtPV08
+6ssIo/qO3dkIFZG0N1ndXqGOB6P+GW6Iy4jhWzTb0eGiVRGdRXQ7K6dtkvHfWEE9hpNHCwCVTRa
PlzyeFsPLCGBMwXYqe4OBzynuwg+/yoOnIAXBWnNH4XnK78P0s0AakioMYy/c6THqmfsmKUZi3ZS
2srGUVIpB/81n0HeGmc5Zk8BNRISWOUI5YB39T5C9pYwRCBoxNw9vmoc/bN/ffJz6AUFnjVY14b0
MajmlCeubPdBWfPB4aPXj8B3oP367wde6mHikq8kWuVvnwOxmnm59xemsEF0Jhh93iH6YUrdsFFH
mx6NcIW7OwYe2OvV0DxzQJMLte1O10OZjoHRVvp1opl5ewQIztEmC5l/2xgt2FhSNaAYFiFgOmhb
SpuvHhtUG9Mk2WCx9GHxfmwj4t5mzyqvLE1tMVyG8V3aRYWCNchuCu1Ti95QurpNhe8NemJRivvC
74Lkke+W7cxsFmJ4xoqonBWwPxMd9BVddAXzi4t7UeL+raPrNpjtE/5lYcqOgSIudjEGsXpUYJzY
sUr6TLTyxUcHwTSk2ce23dYg8Bmdvf2ZPnK4a2LsYiGu05oCTjD/IWB2rlf19FiT31rG9rKwEQZJ
rgPRx76uyN3J60FxwlDkLPtWanA0a7+lOndsY5KLLqBuFsSSarJPzFmJWME1PTWTTD7iXgyTzSov
lFIR7d3gvKxX+7JJrkKIRXIx33rbXP7YVipidnZ4x7j+YqRKYgWHdPZ5ID6kx5DndCPEKPmFus0C
ZhVmB5H/fvOlDo6Qc2yxSutuGJXMSnpofUuBEpwwyvv2oEK9nnB4zCbykCsAj26kPseTXT3P+ghz
/DcfaGQns82siMP1As38SzzlHZFrVhxdH2xNOz6FA3PyP+/ypLnKUr+jX92dFtkANVXQlBqt7Sef
jBOXu9WbopRjBE4vy/Y2tqkiy2AVz2PajCPF3LiDWoh6glqjwnZlneR3/eOHkqDOj8dzBcRgjYht
wUq8VnjbuXHTqk/iaSvckNHQvQlwttOBREXdgcfnpe7Wy2MfkK3cjGU/pcjRdO2H//uk54Tg5I1E
YB+4wZeM8hmJwlBFJwJF/e9/EZrgUUzDhZ4Em+XXJtCT9CwMozzb8nsjsSeocVl+5OPqqNAM18UZ
AMYhqhn7zI70bx92lKgukg6Vx6t4W12oG+1UnWyu3StBRcz0+3hUHx+Ms+5eYJw6cbFGpwm7p9Hq
Ed9trTULnXe/wTiekpVMWSnwPcsq6deF1pDcyiocj1J7/pYemsEdhojyzplncqOHlqj6SqKGqk4S
R/BSTOB+m8McLZEY0SA6wlY0s2AhJEUjnVIinRF2glL7CSVy6JaFPhjAfbFraJcB9nrFCSOHGsD2
yghhCTpD43OafHGzWKISGmko8lSFYF/xTVtD2cxU2pS3R3O4405t7ET4aXlEZblH3mvy7nFFYuoY
B4GeQ0AjKKc+/wHxDKKLJUiuMMA4da9F7e9Spz9gq59INz5VhpixMBA8Io/uotlzMhcQTqnp5ngn
YhD7xlsbTpgmkagOHIMOIRxn7hT4m67qcyd8oG6eY1ewjCxrf+ao/ECiQxMx7UzfS5+waWcG45JS
w779LPSXzqmjgGmEQQV2pNEknK/oKGGn7GMd4LV0iH2S89+zpVP9VU+97bBooyREMjrvNRk3ohAl
bkXGo6j52a8WfwiGHuUFsZy9Vj6hGN2e4UU/+xJ3VnQfx523G2kdNaI5r3crHcLoH07sgdgHSg6S
sZR5FH3IS2VK2yALXa6nqnslbyxtLtUvz3oXxMH5qkUiB2Z0+DBV2Tuo20VArbAMtbOjUAU1ciQt
xrrvyMxbi22EOT6KmQ3XTAZUpoufjOuW0uT3Dh3kWFLjLIpDsmao4OIs1C4K08PsIg2Q+t41tjIr
TkDM+mYlB7gDZaEggLwBnYXrZOIj/Q4AnXeJNEKgYWmoU9bmxAAKeSg0BCXgnp6kFOBY4FuhhQ9A
t8vL1BQ5j8nCTgJT4AOFolpUMOW2JAQ7XVVgclo+RauLmE7rN23Uc3gbtcncviNXC2jT+inpm+YW
I4IaUX6FWfb89olgOG04SwOdU6MAwJzCQ/rCXSDjyJeIBUjxVSf2qeDkcsPsBdaOg0AO5KnNyTOs
nPW41B3++8NsziKzqv5S481Tao7ET7OG7muGjJp5+ZGx6TjhluEklBMbWmR/TdAjngEu3vji+K1n
NNKOhJKYLdh/Kj+/y9uObgnOcLmoE/BeXjHuH9+CWX2F/+y/X/YH6VpnrdI4pU8BFqtgihf/OGbw
s21JTcFDtCjzhCE3+4+YjNy1sMBTW4p+rbaDrvaGj5xiHljAJl7dUFCjFgDCVgRJjGFFdXgb1kMT
+C56VUBvV2F+I4DJyZ/b72lsta21zkDlMhs5ECYsYR9bYNYaMukfMgu7MzXpOgoUlhFFDwm3r73G
RwY6iTShgL3hl9IbDDUIu5XFyM09VCgrMxx3OkNWX6/Q3wubCXbufWpIVA+UolPzx+nPJA90Jd/T
p8YMJ46+yJ9IzvWnRarvphtA9A2ZHeHMPOThwLQybyi7jMdXN6bk+LCg+Q1gCrGPUCtD12pdhDcr
42jsDre5KzdMZDcFlOm4gg1Cy5/hEW/9HbF5NJBbcFLTJA0Fxa2Ve2VLRFLDfUPXWiJIDrDC9/aB
Rr+rGfOq2y/qsHzeaDlxxjWT4LXMjFdFgblTe9iHSzD4CDZvLYRolUuO7Izy2o2Pw9knWZCGdzRg
Htbgc9o/6JAq1klD+xn1tNJaXBx8M8V491LBZqEGLvRMv+ftJvGyMaIF7Mspt61jqalJiJdGQQTD
aWcA+tM6Pnz7LE0IXpolDMPql7XecNmKKNyOT5lpFNqXI5uTMcy68ruBQbtRCYG1kbwLYoxNBdkD
FYaDRg8aceqHV8NmeY280gH1XZ8EoeRnC9GM3INE1MMWKdu2EjODc/bfEJFBxkX9/eDkN/UNMP0K
NLZSBjz7JI/acPNg9l49I3IjEOFs0JUw+R1irdjDieh6XIPMuWBr8leqDw1AC8moEOzJ1g47FV+j
Q6vadp2HWTZgzKFMrzpke9d+rXbRSOICoOKgaNpj1DBzh0h6Ud1HmO/4N8GT1pJfr1nWP96gAy+S
zwS1IHAnXqo4u+RUk4dqRXd+Zug2L7FJUioB/K4EaB/PsA+Hfn652HTQZf2X36IByk6UpeTk6hue
goajluwBmdCbK9NS3QcfznRqIW+salHFzIGTXWXDjLuhFPQ+9VUtcKuhn+wPmylFKy5ybwHCGHfH
1zBZfbwJM5C4LYT/ZL+D9uWRHJyrW9KcXLucBbjP0FQszKnz1A785dBSnqZzIZnsMZfdPHdN7W+C
sV5WjbanQv0Os1uklFXl4sAEXDEA+MIRRcHa/QH9W+NWuaTUy//eUtdQZUOVA78PA/eEyD7w6CrE
67r1Z74YbytJjQPLBG+a3ToXKe+XFTzvhOFGzSYi2I5Ogipwy7BFVjofIlwzmlMajaM6tj1TwaEx
kPBYAGSdimah2TQj6Cjt0Qe8q3y8MihWiImkFcIFQ4aoCHcgWkKQQBbckfy4OSz0BO/vhUwDSPNE
UAUU/QQbvAdj/Wqm1vlJl0nIKDenQhjg0Y5bfNpLPq/SE65wh0rXGnJNR8HS8LCPc9+F6/QJD8OC
0nXGZujl/jlW6t153xWl6LHYJCsJENgTZv2TAD0HKEoHq6EvNgMZyNumwKMr3J0h5eYskLwKgtHX
g1kgFHsvffdQzTj/tN3sA03YNw8HhIzn61dKcH1iwYtMLmvI0pVavHZaWeLEMYfP2Jc4CHBBYk/x
kFH1p40PwCZ41lOPFspp06isSjASsWJkY7gJAsCBaH4tOyKzq2Phv9lhHe0d0xxfp2aqWWm6qeRR
d7KNzbuz5gwUk+uXM8eBJflFMCudruseb82EJVSR8oZIuY/m/xRTwyL8xUdbMzqGPqNCZUZ+/QVc
9CSqGhk4yOJpCCV82t+PZhEtCnt287K3Fo+MH9oyurdpFGG0Z3e4xaRbxcRl6GB/qvnh5jNd/yRw
i0m2w+FCBOBSxkWgcT6NCfdIh8bHI6pFXX7V58Xp+S6SXF88IT9F6dRftJMcaogS7LGBdXea3hzh
E1qtpmpx9Js2srIrZQj7pbUpOKoJsONlSN666lKV3angE27MBF+2sx5QHGK1CJ2DylPuvhYbp0s8
X6OJdF1eSzJBeHWqxhwjSnorhX09aUVkZw9MDvgZ5P1aZ8K1R9HuYNHr3kMdgaV2LSCQTfaaSyel
rI4quRlO4yzasCW4hH4+xNTVDvrCWnGv9KTvDvjGQrqZGy098Nd3ejvKFur/iHcqUudBpj0dLCIk
yG7KN+rporwGxnII88qrSqnA4izjkXtqRwOMVhCuCHsXwa99g+Jm5SY2cmd9V7k1vxpC/fPCAxch
7nbmcy9DTzYzK6NnRftvRGsBsE/0PHTLymM2DbO+LU5X9sN1MRZRb7TnguD81HbjRG3VThfvtD9K
JWC/XCe3emw9dKr57SvtldwI/Euvz0pGBxjCPO4PllNIR9LPyZxz0DFfsWUd+/U90MQrnUJld/zI
ftrQbz/PrYzew4AA1bR7Fjlt+6+T1XSQCBFpbXMMV6tuTomuMvUHll/u/Q5muVOX+xkdcfxpGZdX
dlVIK9A5cUJWsQgYYBraIrGKaJfTxoQ3HzWGLATe2tGkJDauP2xbqWIoh1EHhOq3oYI5bLXvo1TS
APGBG85joQhYAfIMYI81e791ZTfSLSjKsWZvd0wnb0S4CoA8+fGcqbU2ZP4Mw1uSl/wZ1upK2rPO
3gLizx6PY+1U9/6F/fxtjcOjalpLvZ07ur0MdFuSpBh8LdgtJGebrrrGfIp15WeBdlQMK/8H9QyV
8n26rm9spPz29NQuY9xXdxqkyXCTWFUFcOu+ji8MoIPYzGP5miiKiXi1hodtoknCRYpVaUNdqbgz
qfkwZAUWPnJluecCo+y5uuFVJzOrFkN+Vz8HQ2+SKRTrcTwRHLDKdFasAtW/nCi3Q/MzPjoQ1mi4
xVpeR2bTshC2kbLUC24jKwP+7B4YzoxdbfC4cVuINB5qbclmueAkFgd8bCv7R60FCrX6aNKAABms
Nu/SZria2NRlWq5MHwH9wpSIdOQwHEXuxdi+jBIReHz+LxHisXUy3xdeAoOuyQQCq6KCs2z04Tsb
A2s6uKGSBIaje5PDkc+EiSs+pXZ8jD5S1X5qUEilEK35wePET5Oddr7KZxlXC+ufBWrBJ/RfM1Yb
kH6o2I0SJYVuEpbSmO+hAB+oQkS6sTBjx4fyD+WRhMnq5U7tA5Lnpxalt49F8ARpBtor2+IiP8CB
2ltAqBFCxHtaGEovGn01Skgdl+p58yGKdcm6z0T79K8RwsMwUVvVjJlWKkxVxAGyeg46KxRGjlB4
VNvKIIxUtDqri0ziD5awpNmqhGzcByJTyjKSBAHbMg1LGxVu7FYs+rkXRy7Zq/IjIa7PxZS1r1oT
/ICCCg1iI5UpnWpqRBvO+SIxGAL9VqLd176qDBYX+54qOQwhzahA874nhNsqXBoWLCJkviqipnQC
Ev1E8ihK/xE1ydmmrdFgpAxmDTdu5xR6fPQIARiZnK+o7PF8IydhtFDw46Cr/SbKpmRUhgTo7LU7
CeP6orPL13jQDJZ/kWQDdYYKnl2c6qLO2kwGzTqNme2sKTYvm3jy/vhv8ln1WliJbwpRgNLaV7U/
Mo7iD9fjB0rO+Cgmi7LVKbXUccCCaL7taVtaJO6OJgmL2EgBgWlg4SpqnzE2iEmvbyIVAj2QKJLB
YAnoqWyAhzfl6tnJhgz/fbzQpK9xVPapvwyzPOuCloXhLW9yFfF836Wf6aJd72yt74GsMDMbDhvG
ZpPrsN+koIWFQWSDudw3pIV/zCqauvvOej6i6so+KrYeAL0ku3Ol783a63zPKZOnTlEZx9LpWXpd
WSlpaXW/T70BYKwDlGohbvOGJArQc6c2fcMna1c+nt3FgpihoZ2TG16wOEDdNe4YmE4ctQ3p7RUV
guhVpIngud9TZZD+RpKvb83ir3ogFtHs405mewKaizNn1YPi3t90mhWLVAPGTaBpU7Yv0Pw27p3m
tih2dd7CgjtOVJs582Tx3zwmUNc3xDtU2SfKeTkE3nQ/ufuXp5vKEEzA9NTqq4zNUNzvY7y5vTB9
PQ2S8/gm9vMTxOQg/GpXqazTHf6plqiqMNPIdkBlF4a3qoje1M5oT4e9oAmxXa/CkgjxSvA/+22c
KoroxzoT25EMjUbAKly5eE6ULo9n0NdEWH1Mv3sYsC2vW/cYk33VzOGEAoYZVOHEh71geoLHnsci
8q41CIh+S2rcgK9k4UWulj+nppWn2dlglvXbqEbsR0V4ulSsXbhADezJCTE5V3dqS3LqtwDDaR1X
5+wiPSf01bthmJO+JcEw5Kb5wT1mUKZXK7dq/XWsFqtrw676Ka8b3SxEkLlOhCe1SZCGXkGHijrk
VRkn44sq3H/OCoLFcfY8xWAFRKUEKf01F+R1DjX4rCNYio9QgsDo9i4tShDT6Ohk1gWDT3IysyxU
rqeCZbm1mYIs0xGrUA3XvtjkIKQbePYFV9scjNBBOj8+02ZEDtgmDOpDPm5UgTvstEXKahtEkfXd
q1wbivWWN3yuaIXqHGY6zTZf69i69860k9lk2RNYqrf3o/SerAFg6XpCcz6mNwhqy3H5JMsk3jEa
cL8qiaUJiex71/b21k4gQrUWzVkqYRHAPaW/lkEG7I8N0pB4QYXwVXw8T0Bdp67m9aZyBwQrjVus
ZgpqKJhM2JrQVGv8gGRu5JzPAcv3ZdCAXhMPDgoU+9IgeWWZj//gYEAGSpV+KW7rA1LT7mHi952j
OLG63zmPXSBppGFDcEuNQ1KQQYuizTRK2ayQ1xmIBLcytbX1DJzaxpVoe1oVtPxzhsNUzXWGlgtZ
QE01Rgy/S6gJcXP6rqpR8m5LXlRfM4eU5G+AMa/hyz8F8KvY4kYDiVNXA/a2KPeVYdlLO1Vvcm80
iIkKkBVXLKhrepTE7+TYR7q1HXZLvM/8DYkfAzDTkB3be6aZ8nvBpMWRl5Pa4DqUv7LJDvMJd66r
a0nJQVaRemSEZzPe7hx5T3WV3MOw3+/0YcE9IVb4fj3MqC/EGCDqaQo4Jg8eT2T7Uri14VVlm2vJ
/ruknL1oN4MOVrAfTjWeKqiD8KI7ztvurs6vZflCCaxH9rdDio2KxkR6Ic9bRLN3RwkNVUhOe8ZX
LoTegQZYCGYlYBHgLYtsbEeBCshHxJHB03SKdawct+3vfuTnOYBdD+T9RTeg1dVLN10UTGXPfRpf
yRpXhTSDMwZHI8aRa1yTz96Ncsnj1zx+ZO03q3U4ZA+VRGBKNfOxTuuD6emo7HbXCz1TyoX2T5V+
a80BNGthqS/3SpZxsfjo6k+nZskFDYm43t2w1lA/ZYLi4AtKgT8UuEDJX9qY6+bLQ5zPzYCTKOKd
zHK2nlfpevyiaYfFXLJw388+ZTfgbjlHneYKAFZT9UXV0pfqGeQE87AF1s4lFkuyrOIsBk/Z6Q3J
6z3YpStWv8G7YV+ji+lJEndLloNy4mpWvFeImKrLOcG/uQED+uYj/kIJfBEBKiZhljqBWd3+ld36
ZVKE/j6ZFXXhok0rmSxfCQTczzdpb4Y4gZaLwUGtv/sJsZhGoYwbGrNPKETeaKaqcKQk3h/TzFDm
4mGLLEW31xQT4x2G2WXevhm0T7nVyLsvUToEp4TJ9YDRsWkRPrAq6OLEHn8QAXmcsqm2O84npXTk
C68/BTs+zeFyKz2YINQ2ld37lsY59EDvhvsl7+BV6x64Aol0YxlJ215CZ9Avcwq5VfvQq35GM77g
Bz/CO1XnkzC4WxgOr4xBEBckHU2Vp3jbjdtSS1Fei6eU/7XwwGWZhqqSDz3U0nbV+PZKYMVn6hH+
ymHc4e1zDD9ok/pKyHB0VD9ZzhN4+PEXJo1AEuky+TyqdIphiWBnZkIibNu67bwUIjAzEIKztoF3
I5iPZHL7P8k6dIJbnJwRcops4GjV3bwHpntpkI/kxA2CPUADQaq5YEkvdzHm+S2ue9OC8FUNauCG
Ect/rEGy3JQTxlvzYcZ9AJS2qD37WafwkJJFqkHCWM8LDWGveZdrt+AcivhGBn2pFZPvn2uI9WSG
LAWnUWEHeAfHsJuFVb9EfTcd6T95lCrsgTdZ8QRrnSbVdOpcZyZBN7JW/swHNqsu079gKQj1gynp
tkUgRCatBHuNMqSM5fhiUGe8mvUsHrjc7cRFa0dwPWHKU8XbRBnsdXGmRxWtnz5TcSKgadMErVR7
5ecuJ2vvoZ5IwxZ9v/ja+w7YQt1pxoB+FQsk+ZxvHr6CY34e2g17h1jCBOeWxZuDWoQktpGp3TVc
WFmvBGt5FJJhMntcwiFsVeGqi0/AFg6GFXTuooXlSqlBkfj9r+zU6P+uiXWGs7Ue3wZxxKE7ykvD
ElZjYJ4vyi+AliF3AStZ1SXNmzKd3kQgvenh3e3r1Q5SpXB/HKWYQUu4Qp1jswumH8/6wKexCR/t
K5kCC1kA33B5FRHkmvTAaKZTO5d9+yLjb8PE862jxmDjMAij8ZS7G/VKCOu021/4dht8W9VuCksz
5pY28E4xKL7yrsPqg9LnPuhDIQHgG3eeOzlYW5Vx0eqR92ybCTLboZhENMxnJP6tp7eeyS8hTJfB
Yc0SlKurVTQxiaWwk8atlP9QJrzumgW0ayfbMmmaRqk5Zm+eYEhy9fRIY1KN0FVnaxu1PIOZYU5b
eov/ik1WBhKZma8eGcbfvnYDxluFu+hsN3RqSoMwkzKBYagMgW+D+8vIKTZcX9Cjfhj16XQG3zm8
6GmWZs1yCsQo+q/YnMVzv6+ct+x1nJKmPTQyyWcYRePv42YH6b/Qk42LFjOxW29oU2SnmJDTnsnt
QyOLowFW5LVOgXF5ejPCtyKrFBmcY4MdhyjR4pO+LJ0t6SnN0RokcKK1/ATkpCMv4zGmcHU35k/U
gVtX+lDhif3aW+9baYUDJnlPWGZBR8NRrrIp9LO/H9WPZ+QNddHWk74GzMbKKBwx1myXBxQ8ZOx/
JO4vvx+Zf0zaM9pUasXJ9nYq2iMe6L+Dk3+YG3gyVCeNmse8OIZtsSUhOH70r1Bef832hmORZ6k5
Y99uxO3GVjeR/Z5zfEbcXjfQVqiNBSHYIkafvMze7YUSIl3sunCjHWup1ZiGti5d8x857PderklA
3IB+b+dWpOeJDgRIjF6wEyZn+Xd/nmYU1+LJQtLrYCFP/j+bk5a3uCTNIsUULe3PUGGmlnqku8Wm
IR+v1Vz8MWhr6eC+SdSvqJDIZhNuVZKXY0VmRExn3NayRNOPvRfLGetX+4JWaS2ZQuI1u6dimJ1F
LpjHDA1XChn1CLrOtAnodkY01OKl+WwwwqO4dAjT7OdddoZ7f224/jz1Da9DFIMTCwco/kS2bmfn
lgCGYF1uRrP1C2EbzK/gtXzqxQWNDVL59xKpKTLwxWKgdL6g11bIRT09f9YnLN5zBKWQEL8YN3uy
e3ao47cAobztDMwBkLueSJAx8ECb6IjSNq5qnPR7RSBMrq8RXKGegmg1BKp9Op2CGCJg8R5miAMm
zW+c2ImTtYwkx3ZXXVWvR8VPC5EtH3CvQk6NPTLKRFAWcQkB+OaPZfkxmNBG++7xk2FOBXKLJukj
e2U+xeFMZlzUhtwXcvbTY4v0IwVUj4lTqjPEWV80qO1djZrEssxQnPPHYSla3a07Uem4uCzORtt1
CzEVxgJMf5HSRX3AsIPRfPBvJ+CISMhiQtwvYludHSsiP0ae/ULou5XO1lR0D/hF4XKfNzo61PYy
9GDC31NDFALjsBeTC7RB72EpkWlocFfx8Za+2gFVXNwOrTIj2oEydOXZoWweudDjbDtaHPZJuwTs
gTW+z4vchvQmNs74M3ZRhqTBcpAYJ+XQL005ibPQ1gidAIBHn78ZhFEnx1U0sQQfH8q7KK0vuZhb
rBMbutb338i+X38PChnzFgsF7ZcBccxZkX8F/TK95aMHbGhGkiHUhrj35AtKAxVsHIzkI3l40j3h
xM6AgJCE3saCrbRUd+5Imkr0KWo5ANANPam7oczsDGou7+aVEfsDP4O3jl2DUNhu199LOh97H/3t
/mAt7OMvLSSmiDF4FHdWGTqLESqgn9DQge+LgLOzQUmC7h9b8KwQ3hTP3zXkrCXP7MOtuUV7Xn5x
6/ehikcCNN98k1SYCgAXf/l8ZmNRjlIU2L8CTvJjEn6ODifZ3rRRtyKBoEbP0rO4zHjEsizWuJLk
m2F7YeMEXDDFKmoop9bZHumfxfHRWxg6aU3SkM5RyphpCZkmxqTwSIBqUBeMpkl2u30KgNPox/O1
bq86eTc/ahzbW12oA00f3MLmvQCGfBtKDcaMR4KoTcOP+Yohm8JyCRNbO5s7SYSiu5Pu5MQZ1pIB
S6yL+r7jeYywbbw28RlAEUHOM0IrqE3NkC0+vrq5F5Jq5bU1W97k/BWoe0Pof1AbKcB55VOygrF/
q29XSiLzOqWxh7FshoyvsXUihjnZIIMqiYnJ/MAd+Xm3cu5zKrzcWnnzyrE+t6f2nLOWDa0S9S9W
gyWtumTzo9ebPd2OGHXYsQjNQe3cPFz5jB10phNG/opEfx9Vp491Vaw60lFd53ePyyML+jG3zKCv
pfUQ4CACFmXr/eIfrloXEyIjsWJXYWvUu9QLlnn9J1dOWlDu2T4wyuKaofAyD7qmxawBQ1fN5AG8
x8FAFOGiCVZDfiK0OD05K/wgeQg2Ft04qWV4TkTLrvQ1cOdL7bIkB0KBxNVfmmanXrQTXUhRNqOn
sjcwSbUxU2LrpQfFCgtAenSsoGUGlfwK9o+kShZh4sUH+vgITr72ikVm0LcIBlyHo5HRhTsE81xC
JCNNt72zGhJ7rXUSVktkghTiIkdgyiBAX2QrCx87sXduIvAdoz1shrKI9lty+18l+9PK+R6vC0RL
9MtsYdglHAFZRF/5ilRXzYvCLI0fLE3139LLmUKPmuxPTZS+fxCwt6mU6M3DlTbS5GibHu3e3opE
X6PheQszhcQtm91ndXlOvdl056ZY/YjtnDsKj37RjENY3Enjpk9gMzkh18SRSghfUYfAZapqzjtS
y9wL20Xaz9NHzvOMWvKfo/6fz3B5Lwngi7FmXenlzZZhcwLErplAKpD/rP4jNusfUwWWvOdrgj9k
VYVbEmvsEvVdXUg2Q80pPdunDE8+n5bJVT5Xk+leMS3acRnLuBnnHhOCq1v6HiAjYgCdxvsnec5i
nitB4HiAdoG2FLHuHK9xpqZW/57nXqR12AT2JskbK7W/6nvW4P88X3oa7G9SQTzPVJvP9pac23tG
01L7cwGrT33QgUYeDpqO086xYCO1AhFKiqTsmZh5Nlu63HiYOWJjNpiAA9+EII1d6hmts7JFNEWL
rZ322LNG9hxc5Q3kXLyFGa+9bTEkqxwgZg6XoY+Svm30mb/EvKwq1dTtS4Rc/qNEprU/QSFU/Kdc
sS9JWLqvHJNLRGQ0uQmFzuchqh5rJhztX5Zqm/EJNzlHZ8bMc4moLux/qrlszL1ii1IWi9bYV+IC
tv9Ivxo2nuOnY3KJBRAO2tW1O4+ym39mTZNQSRonJgTgJBooHto13sjQB1MnKSTe0CGcJ5AUUCmd
Q6/CQ9RrH3BlWSQWuPi22YUdbsPvizSC0jiEXteMJdEUt2QzcdTeBcCaqqfPFxyjTiAnNWSnLLyX
WwnV/pHrHzJBTLGMIh7lvRW8KbrCpkOj9tz3HumQBEoXEqMEN/zXpO6ME5+xJy/JYIQY7gjC0PUV
xkrcpbet7DxJulKEinn1W28+XoEmwc6j+dH2GmWMpwoOzD/1sH2rDtODcQ2opxJIW7E0NQhyps2s
yXCjxLbH6srEBDdQ0evf5Uvi3MW0V4iwiU6/9UuZpAYOG1H9lYK7PayzmIZiWnhBA0QUA633qH8r
0z8slMhLzIBYAMpn01Y7k9/9lhLmodNMlWuKip6p1+x3BqzJROIMZ1Pg2KzsDkqVIMkNq6U+ZKC5
WNeiepP7tDiKriBW1ZbVP1NUOrvFEMPRNFqIrmePLwWzkqbNlHPoJrWwGFVfMds/z8iV6cqSy8ND
e3SEhlG2hzzslJhs5KNOqq9wz5ymPnuowWaSjuM+y2rnWjb2/+6NjDcRMrau/Tg8h2AgAL5Mh4ou
Z4vklWt1MtnWlTSdFdkiZWx8E8EXjIC0pWkOcxZghoNiQRNj5BLX8eSRaSuTpBA/Ul20DIWge4jr
MdGWbvmdNltvZloYCqs4vKZViwSXIJbJ+JbFCBYoABR3kVsk1ybTaq8iC73YRdEbz1y7j4M99OrZ
N5xV/AtnGK3Hty/OkOHS+kvv29BVzxMYV/4J913mEvI1nmmUGHfEAxMPkxFRUoNFl9gtEL9FZJ7k
0RiJrpqnpy5w5Kfv21HZupxrUgrjs9KUBeMYwd47c9pEDduhguNUbAuGou15GHvyteJme+4RIYaK
PZzgU6wd7zoeZuNpXwOkYA102SjOZPjyF9PKRxfA/pbBYIFD4MNTJReeY/Wi4AYKQuB30jyFaQCw
LHA6MOJc8kXbReRAEFazu9h8HMZP6AToq6Q1r7O05q90cNDS7EKHu2qWbtJLXyv6jzScjhsB+f9R
Rek+RqQdjLllqtU6L2aXc0kzAzxFmoVS83yjXS2qWrpmPVaPooYH3v71G9o00o+2Q+8iicrMYM+u
XkK1iFb59rcfxDv78dHSQDeYkAnw0R7/OfcI3LabUEymN2iewNk2gy3guHskA0hsanK7axuZtkXU
NFFGrqHBzxLkVAjCUpOCaAD5V8KGPDMVNeHu+hF2reNrvxFADK/0T8EuQSyo4Jofx1ZqlvI+FfEQ
Q7pe3yK+0jSxnm/8/JhYmubVLFesH0rKvAy5gnC8z0caB6tDSKpWeE/cLAbsopg5UuYRWn/78I7H
yhC2FDNgmcxpTvnCNRNEzlG+xc5MT5NheNtYt9xQ7MDqHcSM7kVqlwM83sdAS7NVXP1ekyOz4rgB
yJAkcfxsSPPqQy86M1gpPeT3N6chCu8CkNN98Ce29F6UmvrfoTTgkS3BHzcaTazY+YGQ+eZJluwp
bgeRIcV/qjL47Bbm2NDE/P6nQh0CFVvZBRrHbktNqswjslh6NPcHgFjQCDOT0chmIeo25duG63vL
gAD8byJuM/P2ky8/OLxdCnl5U+CIvjFFxvssZJw/l+xhLFHVsns3DQHGijqDNv3E6GSr5B+UU0xE
LUnRjqw2GNNKsIBwqZu8c4xlIe55JCIK04BNmh8y61Hz3U6S9R1tDpj0AyUXceUZEmY7S3gx0d9h
D9sZOaGXvEjAdZdvBOYz5YJ0eqgylfcciBIRdezt1tUGpTR4m0VBg7h26FsnYH3sPhYUXT6Rq8BC
X0rKxhJ349chL8gLfYxGzUvCWWDDBNZ3qEmr6AcGRtfGRo5q7+JBjRDDDPVNLqf96jFtyS9IUE+h
PEP8SmnXSbn+3N+kvicrR7HK+9ewVMa18gwxFfCqM4Fv2LYMqnhNHhGmMLOBRimuWGcO4eZdI3K9
0iJ5gqmHjzonUjAeWTE0cQD/x8BErvhNatOJzUkX0kMBuoRZzB7WL0pQ9a/jwAM1DIfMj/ghpQOp
nQoRZcDZsM2Paqi2BY47o7wGQfJAUMcjrZ5SJ0kEClYRpKBVL4vNxJpMqm8kYcTWa+d4mb9s2wmU
hYkAMtAC8+/p4k/huDm+sWD1pmEmk/oHv2u2AczKOXOaFlOe49591FiH64VFPDvi9V0eu3UBq+Kn
kh5SiHEI7topX9UiA/CicCk5HeQC3byG+mQ/YNUQqxbcZcWUkWewq6SrZM+2XQbqfW1EpQdJIqb8
eFcQsgGTyH1iWgjo/opDA6um6hpzZZnsjZcYmEk9JgXDE8AIGok16Y/2Y0t2xjmy9kNp2JDcylTh
UHG3CG1n4+qrIY0s5PUGs6JHUt09fPvQIJqOrLMm/+qJn1tLB3fpnIeeF3OBVJt3JIJUQPHrYt5B
nz55RmDeazRo3x70DGWvb0RegVRCMMVpXC9n1y7133aZJlo11e6uaMAK7tS46BK9McIrDsBTD07i
keZTv810162cE6qluynemnloIOF2SZIDuJszR8Yv5qGbBMUxMkNKbdbbP6YCeLnWZZHha0X5yTID
9frvdeLc1Wqx5ITic40v6toSRiDoPC0O5X7EK+D2wNL4Vr3MM1FBYkWz0MBDmoz/avUzI4Odh/YR
xJTBvvKRESKLWjzm0Fn3ZwUSTtQWfuo+/+O6jnkoTQBGx3sKKkFspP2/jBZROY0kvOiX9iAp6N4d
wR9+74ebCDs4AX89ayvIL/I6V7cH0IpeIgpbOYZgVgh0XI9ICKsi3nYTO0e9b7fKiy/rq7okQbTh
AJ2ImOZtTHV5CSanHl6ImfwMhtEg10jXJdg9zTmmHywL04LkPaXP1czpMneZQRfYjTTHMEXwwREN
7bXyJDdA1RBWMBAk2sqKd0efmUMeRvhTfU1VE3I4yKDFcliLbU07h+IeDSz71Mp39CkpHCo87J9s
cjOs6Yo6yVAsfHBS25kjP6uljlLoLPJ2y9eoLYt4/hY8Kq2QY2d18uor//Zj+vgsr8Gc4jG7DyY9
Fctdoqv/r24+/sp1njdonbiTSzvM8Vs1JM8rrSmbWt/OKQ5KAJYUu4USBhpa8Iv6ThRITXyTYO8T
iGXBfU6FPfEhBQmO4scw6qUrmdDl029sUY2VhdnKkNnzgXhzyCXRhr4EBUDXuRmTvp004WDIEGlo
dzWqiEgearseeOzZFxAgVjrJl2UJmtBDBZfHsU9DbCsbv1yaeASaCblhDTUopRcsAkln7LGNpERf
3ZMJVEBfdIIgdktWP+iMrhwV/Dk7K/TRl35guijsy23+OePnQQ9FSKD5GItLqNrs/5TaIh3XKo6x
Dz7cLoSSmNARa0GoaQa0morueohu0fCe25f7Mrxr0jbfImreUWDjY6k/2rVTENk5hHYfE9zWQCy+
2EGqgI2jJc5L05y2z/QFPY37B/7kkvLbWh22vb6F5ThI7ajwXfhcgSI6OUdLBm1KG6W8fz6OearL
OooY9SIYxNTifYIT0ljvw7J3Xqi2fcfHZbYSENoq+zpLHnL/Hdef8QR9j43zb4pklK0a580Uv4Gq
CDn1ij6DT/vvKz/EQ4n8c08GoXuqcIY5oZMzpdBvSmshdAh3wD36MLquG0KGTnh9q8Mn5Gubps8+
KJ+JljdB9EuI2pShQ0ousT+jMuswC2EBlsoCyl9kNzVnud1voBzNpcuo2beszvtzENWdVj+LDKvu
6INVXDRtdW5SJ3EFY8hVNzJoAsy5fzlFqcqfGZ8f/MA+ydaM9fQVZ3Ukh48vslkdPP/xlIYP3g2a
vSG+RHcr5drubZvC20Tq7PYFUm12Xyo6njiEKrv48pxNyB94f/Uc3xqkYWvdeSm7XaP1NJqir37P
oLpucmKzU2jWuk0aMT7TjdarnZ/mf9p/Yo7eRIHhq0esaA5Sz7Ce206edQwYjMSHmS8R/5yGmLH3
uEkAheQesgydSvL5Jsbs9km7WFjmO2BHWUKfpkJaprdSgIvDfpDf2tSnDDw3tTujCV9DDb2N7Y2H
8okxHz8E/5+RFaQW1L5AYqDMInTy0ar3Z6fVYrpRiJFmuVvMLwzUUXjTNTAD5g5BvmTmOsMb2URv
8GnZf9T0kfyx2i5oZFJbjsVlzqSNmG8N3voAdL8vaxjW4UYdHb92JYT7riwRNXo8Awgfag4xVSSu
8ftJ4Bir2fcaDvUmwHDApG6T+xjWUr7+/frYBYhqA02emcGhLozMbaxbJhbJ7eVSWcigG0r0kXsN
S1awww2MsU7v05MtyN5zmRv9WgoF4+M6Bqeg9FXjRB1jtY19ZodfxBIXorQjtiLmGfYS4RnZjX0x
BsZkKSYskBeJEvkF1Or0tcV9gmsiv+saR/nkm3TYh/rIOwG7Ohyy44zAZSEmhiHK1AjwCi+GD9Ou
FC8u67e6fKXewYw3PQ48ASJHS6zJfEZi5oBzkcbBqvJtMQY9oo12eEcMmhHT3ctP6W7r/kaSjmAW
SOFHzypZtV7xzjEhpotIrgaLyyuCxvsP1AHlKZAtWUcXmVxdFVAGPhFP5W9Xk7GsgLFW+1zkZjvr
/I2ZZ6jws5dVrAclYVuWK5oBWqY6XEWFxvipcDX7rPYfh/6j6nUDsZk719si0hgda897Pj836nEf
V2hEqHM8QrVVmklDPobyWIoPZe+1f8ftJFLv17cQqtZbdw6hFQpVvareGNUE5jLp4J/2AZ24Lr/6
dgA64sq0XnTZ/cQR/lgfo5/il7LY1++WMDNqGdWITtOyiKWX/FTqgGYAQpY20sLc8THe4nVMY0o3
aXIVdXBKyYUup1vjkgInXoOuvyZznTwwv6LlPjxrASo99XVy6Qk7G5MEKNJsIWKUoU6r5Npgabf7
kgtmUxfw0b56ePLqOEKYBJuDChd/TYie3hEj60YIWYXaRd0LaNO9ZT8GNPfNwFHhOcgC1xJZ4plL
7qpbDOnspnfLbVYBJS/f2Vz3SEAJRgACeKyaBhJ7NdxIToK5cj+XN+BsZXfJGya1+5jspo4ZU4g+
qiLaVvTEla0ndY22Rtb05h2/e2LaAnx0mIbJjE44PKtx5hcBN1+jvj6hfLH/ioUxLOVfZx3BZBRJ
g0r/XljBqnMOtAo5GH+fXUxU90YDf9uuORIvJpxjvhe3/w0C/oh4gZ+GI/3oleTu1ptfSnjHEho8
3t8Tb1KQxQXbjvW7q/luztGNJRj+gRB3GBMErCxko7IN+BCHpVzXDBj2HCKZDLnM2E+BsBoh5SkB
qbibc3WXnKPd5rTW5HELaLI9jQsTbJ8v3eW+tA/wZETPhLYIcGRJedBXg3CXkAXJYUZbOm6vQ2eh
WhYV3hxVehaTA3eZ5OPObjPnWwnevHSx5aRy+uYHb25djHhIUzA0rbBzPWDb8VWiucjjKkD790Oe
uYy39p1Y3D/uITfw0WfkMvuxn3i2QfR6nyHg6CKYnBZYU0x0E0l4eF0EkEyy0DVNuWIdg/tmGID0
iCqBKUXMLGT1ZcIW3TjzRheKByd5/bWZ1n3t/4Meqa0tUhRTKBnfTOBI4aB10wKEJ0j9K3C+0X+O
Hm3NCbf5RdFKS+jY/y0Lk58Tpea6c+U+DahfJ0Rx4FPa+mLAbTEmlLXHWIUBVDUtYPyo+/Jsddyb
Lwm6yq2QpJBx/U7rL/ha0HFJbsAymkYc4imEL2m33AUpOrghAPxZt3+VvBcEYplLVRvx6dyfRV6m
k//BCBwAtT61bR5xMqhRaq1OjiAQd8nEMVK4WXFh8Fnd1bUm46QfIeO+oC3NHfNgsUWdsxDhTCFP
zra7epk0/+3T1YMvi/JsGT5SP2dCK+s3AT6RHOWHULWmEblrjBP7fjNRqjdKjMhP+Yl2MymVGo4/
vB49NfjY+9P+U6rzLTG+ISZVuGbj8mQfiFmsKIF6HyHhrfqgdNUGf5W1WFvQ3qMY1yoSmlnQSBgR
Mp9nHwyQdWVcQJz79uVfkFdkBsB2i2MmmeF4W6qu4t24WIzNakMlIgsXwU4UsNsAKi52riNFeL88
c0yf90uZWz3chHZSQY6MciX+o3tqfEXcXu2IlKqTv7p6gJoj/vFvMTx4e7gHHnBNzmE4xF95TBfs
A+xPS51j0BRcj0snCN7u/UZvLOoKvcsgVliJ1xxpPIG3WaqYVKrj9+2JVv3/Zai6QmtUgK/bVLgf
X8M1M7nz3TZsG23rA8O99hNVs3eGX4uCXyaeyQmVphvuF2kQfY/1/nPV3cEI9IP9AWnVUEClLRJZ
/cTYVok7MRkc3AGfkDiOU3RmDjVigITru7KGf9U5ylfldN3d6YH7pk8/FehesIZTkZfOQUzggGXB
Wz7x/Iw91bAhzWzq+6SKWh6LpuvdukuCsWsmzRwm+35alewUluzx7HYUNOKaARI9lR7r6RP/SXXM
QU01kIVf0mQvcUAWvAd7AwEVcvrTQP3n9sxxNyhwHkU0Fj0Euau07Ulcb+VVToqRdl5/JKPwM4Eh
aQ9/+LNynB0KhGR28fqoTNi0HsS0Cm7NlLWA0M+b292ZAC5WGnzYWBHk/KBapKbSZzz+HUre7GF9
yJpSj3YxfWprP240pAmIim6nx9EPyD25XcTS9DLVsnHyt38TjUUqMPbB1i1rZFc5nRkbPbNeBZd4
ozxZRbC9LGImzz0M/m33zk0ibbnPXHcoshULwbgMDWswKDh+NkoJJ7p3qi56Z5aD1YYa9g6x/Q6f
aqhzxmfN55q46MuyGA+K2eQ2YiWatk42cDVoHndfPQV+hU382N+Z+TNHPul6eMWTwo/BtSuIdarr
OxfYXxWgMESYUu18uCf5JC7CCAaaMa655aHfuP80jHwJ5yJwwNu53TmiP7hLuVpaFUmr6PPNLfSG
oRWzvzrYED/2+/azqGdD4Bi3GIPcvwPifnf4/jetKeSJvllhtE3btU3uJG0LbMV6jsDTFyI6mpa0
NwU4nN9AiBfKkQ2KQMHruZ/xWCt+FFf80beE5DQ+ESRW0WhdrDPmsJez50LO6VD2bt5GJBB6FRzS
3VGiUYYGKUho4mcRodjB+0esuzb6rpXLi36cZAxhFxo3c6X3ZZH7DYKGTz5nfba7iHL45MHHvJZa
i0kjeFyEbcND91USDi305xrrDg9ilXJOnrqdjVzUGG64S/xZ/rp2NgLgLgLVKyS4TZwMDnWUIwSj
s+ysstuQEGhP8y/e7AML0A827mgpugSvhJrhAla/Y7T8dzLweP4OSXD11O8SdKbBLsAA8ZJNGZcU
lpnxid7uLkQpL2f2wD7iJjplF/Ur4c7BgnrGtmqv4eQDTXZ8wTgFHuRIrWbkBXYJk4GgjbGJLxqN
vrsJmO4NHHRuG1+Q9Gz2vgUnNEUIE/AYgVxKrvsdEib+mmfIR3h+AqnV4O6M7RzeYAC2seCFbmcS
FzACV/iRZ6h9Lp7MOZanoyD+C6Use5DDR7zVMalsivxNuCcWCxJ1PA8+W41olRNThvnZRrv/q7Dc
pn9a8gUebWea5kPJFdflhyCROpGjrDyLc/jQ20774bxjc0UlA7pPiVEVXWcFg3npfPBhxF8GErRK
9DJomjk+3d8rE7I2XzeMPt0joCjeDITR/z57cG1oF2KCNLaOyhWqqdxV8dRY1yz6oWOCfbjO9l3Z
N3MjPvq0WCRKx5Tw4OJVKXZu5yFHkWDkdkbpMEBcvM7cKuFsbBnTDlJA5Le6AWmfpGg8HevojFUL
on8kGjh+UmevKwgwbbdfbz2fP1ZYKcgByc3gc1r03gFcNChz1dncB0XdPYAWnrqJ6WvB/skkrNCH
W8jypx1DkYBzbeUMJ/h4NwHqzZ5qjAqV8PdsJ2wr54I7/LUUk/CEyEUmdoMJgfIkzJpyrAMEGJRY
19XY8TCKNkIN9hUD6kUvxvqg51MdFFysMD2gbVUxq5/Xr28QwT+58ScpWYBW9MYtvY/t8m07KZUA
gcRN6c9mxbdQVPP6IZuydtzzX0v3eVDcb+d6yBF6W3Nykx0S1blVJ4SREvtiXB11Mf2AzvKxcfCz
QTt9gz0ZfVVExr2hXBzhi+eu3wBYRL5q5e4oJbxuXmfLE9T9u3Okyc3rMz7sfYsHKj23o30DmKUS
0mfo9noWPPOydnWE4Tv17JEkZsruaSiA0B5GkUAr9thBBv19GxedwFO5vbymCJikS5oZJaQcbx7E
HFcZ4EHWGf9Tm9tcmW7KLym6vv2Hx0ZJ+dAO3PLXgN8Zdy70lap4Xsr/m1dBF625EVtjzwnKgFOE
RT+66VKOJgZ7jOy5GrK2QvWsZZwSvqlX0HZ5HrfiueZpaVQEz93F8vZn91o9Q1CJJah8jFbySqoa
fJI0o+JbtokcWdtg5NSSkDSk+XOe9lF13d92ZpAJrR6ygpoRU7LVAR0Qr5pE6hQJBo1NM+0GOU/9
717eA6zUJiYzpI36K+QhebkHt1bAehdqWuPnPG+GkYi4J/foecLv05DP2PyxKsNjX2748ys5eN4s
hIk7axYQIIgE5IuijB1QmXBcXPeNyXvtc/OB1Bc9k1S4FXPJeujM04+q6/8QHW3zLsYm+wnJXkte
Kj5QSivrJThA/5a6g0dj/mjADQaUbToglHpGevp3v02UEKEgNQ+aovvy36HUv/z3qqzsBZk/9M7U
f7H3U9hGXBFDfGEwK+zUBtB2P2K30lMf2KveBWLDPk5G2wj27KZ39YAZvmXCfOIrw9r5mNZBskP8
uxI1ZRNIUiLIokJ5txH7kE37BMlQoiJeclBWFcQAb/80SNcFxc1b9lUQGjzc/lHgbt8ZJ5cN0tuF
/YB1BvspVFc8y2AkcZeao1Qkku8PA9tLKHH/pT6lA618resEfJir96+JAJVsfJ/S0TRMlb1gNnXf
Z4mA3QeUcvf/a729IqjPUlrMzrgilSqAiuNNcSIrIoY5k9RmZgOnAgmVWwxaks52OQwpq6lXLYk9
7rkNn8AK/UCSkYzk+BUSL0uZLnWFkGDf486dqL7AmDHmqJgv6lyiJs1yd+XjoBXYGBARepMCG/Cz
ksUwYxGAtlkHykCtFdn3H/aubaRdC5nSsc85OiTz4X+a1t7+SVKc6gMpwGgMOo7aLREr0gQldnIo
h2wVcuHOCajeZ7ujMzvRCq2AGdKPSCJ3JAPye5BQ09SAo50PcgdIl1KplwFqvHMT59qvdJCMiiQm
rdFJ54cl8vtk2XIFfKijrkV+OxVZSMNhsZb95TGxbRCIL3z0nuIiB1wbjxmOpnDlrSROpvRWPR3t
X3nboACf1I9Hi+5GLy9Pmkzq9PoO7/V2QYzZutqXh1DGyz2swGpcfZFNuJkJ4k7OmCsB+a+XuKXo
kiirTTWspDUzl2E/WfRrxnNAvHzjvUpBlXzekaZ93TsEFrFNC4TTbpZo5baD3S2kWyCdcuQDC7v0
z6RChWFkU7PMeUi9yR6bkAZMI/cXHk/9eFCXQCGtQ/xWhLYfiaK4vCmL9X3qw08H4bn00CucqMEc
DNZuSFo8CACP7VHGuZIXPQwKVVub+4x/49RF7xRooRB9g7+YvzxmAlV+zKsVbWeQRlB8LL6X28Z/
T38Or70XHhljbgDTJEo67uaD6YokaEkDj4gCB7R/UFeivLWHlpWD0Fn9bVu08S0+VtTwRUadkgQ5
wLxRclRH+voeotAwIrRQ5LA1exNV1jZ69y3oBVb0M1au5aueoqS/fNIsPrk2fGugtUO/i5pteVgq
W89aeDl+by0koFa+QUyjtZLPdkAKMXUKLUy18iy3lthdAxQz4z56JIQqJATf5iazbCzJihOvSTnr
AoIkyWgqLjPx/ILBnR9cvf2i/3jw8O3wzgJu/7HvDzn4JyTRUjlja8nr/nc+ajFzTqf2flB168bc
ZThOMP++7O+KBmw3pViJiyltoIbD38bTokatnNPKQEqDWj14WZj5tebma5wHgRBv6QcA38B8UZcU
RHRCZDxxeRD256RDkDV8A1UlSg3xgCZFn+hCS6Vf1cjuIuubb5XyM061bXphgMa8KONRFjWRDzvj
ASiBCFzN14b29pyrV9e+lPtiosnTIM7gNY6nNUm5KTxSPSwAy0TO/2ROAti0USsS1Wd4yA7nHq2V
lu1gAJ6wyxTvEi4w5oXJ+V6S9z0XjNabn9ozHw7LlhByXVSEJh2ZS5fAz9XBwHFsKR5bwRi4PJ/3
FGBnpeHhO6iSfkr8wZMmmGnm0KF1dWt/mHuXzr9+mte28DvGYb0xi1P9FKiOm4ei/c2B5NkEpvuK
fyyx7ldheG5gDLSrhB7TJ+9Nn51zXRjeBiKnVzOhvrUoGUG7gUh7Zjg/5WGrM0NywrVQolgYm60U
KxahNoE8ax2EHMVng1ZACLUYPe3Swf4VMdbHxigrTrqWU9tOdgdLzbaoaowRvAev0Px4+uOpoPeT
60ViGhxHsndNkkhpOldaO9gHooqhacm49PGFZVlJqfTViXEmTg8SYj9wk4GIG5aA0vUG9c7II3in
SiUtE1mvT/ghZyaORe8kCDdrkdL6gu+DfsIEHL2lqC4iEmfYHpTJJ1HwIo8B4D7vr0GCs2fQ4/wk
LP12FM0MSAWazoSZ/jFT1j14g1jnqZp+YKIKbXTlDBRzlIwyZjaUyOeCZ9F0oaCh3Dtp6Hj5grb3
DhloP5AOySm4ynoNc9D5VMyFgC2ANpyjZg4Iy7NuUDN/YIFTXU8xjtmTouiDp8pJPGwFPdqAJS5U
UZfppMNMqw0n1pp+O1PckeNRA5AkMZ+iL2y1dlewvi70zLxw+29ArrSeQ+XnpxldqlR4aW9xE6go
CR1jVYQfNNoVzTkCKYoJbTe/V8ELiTkC/yUYIuXe8pZKCJSITGYbsgpbOIIinJWdrlihXn8sAqbj
gipr5EVt5EQWGCxd6hN6Y0nb2hgLKkh9hwr2VaaoOc0uyodjGREUQx7Z/TCl3QWqQT3T9upUP3X1
umrCIP3/y9+zbbSQWIpS5d+geu56r+1h8Fenas97d8vifGpUdD/eOfcB6zxemRL2Gr+ar7WuQ+/6
xxuYECLlyt9m7aBGgmLabkerwOG7zVaxdsqfngPddjmqXmxuf9LLoYiPTTLyqQ4Era7vPkBsMmyZ
ug55u/1/f45qQIztYloKyeVOezdpZo2plBMoZuod4VTmQu3XZPcNqwW6vcx1zcYI7TWSZ89srhaj
VtH3IfiEjxJKi8W9qMYCV7dymHFQ0tn1gVHRhuo9pEeWxuOHFPT/XRLua2ZVo6KJ2jtcR3EDTtMb
Z+15oPAQO6NvNWOhXKoHZy2L5pKH5PcUg51ZRpCKCzHaUwHA8KYofX3IWNgsdgseaZxU34gfsC1L
tkQShnVFPGrxP973OT4GG/nne2keZTy10S6ITUJpLc7R/nx+TtSomavLkhYsnKEkKePXeDc5ju8R
bRFK7GebTimsAhyhQ39sC5/GMcqBkiiAScYr5Acr0UFo343KaHO+hTXKs16SFTP1JZQCq4jqo9iV
JwvXk5R0gDmEBkNZGEMETOkNoFT+vyWdTYWBKHeeqr1/9/rRB6sLLOTkDSe+kJj9DaZbdgkaekxb
K9TpUOiTG6SBINjbZ59upY/sWYizPC41ufwVLyfOmwiYy9Log6FQYg8/HAJJu5yxwcXHwfxGrqzf
gyRolTnNaHegTzKSCLuZBd82nhiOA1tWuVnKWRXbiu0mwzcJ/LZE9+mrRUgAJgZJbwpJcckLczYB
FJR5QM0CPqeMhWkimUG94bOYTaSqQTJ/RiUan0VRMM1cTiJBPqG1JI02w6OcekcxgrPyKmK8MdjA
vIecIqcWyY/1GUbNSnyGCHRuwAAZvEg2RrPdzOW8xNcYBQ0T9ZWP+fuEkDWBd/sShD86Slx0vuIT
X1RcdVTDhKDoaIKMzHwJ6b0QdtBjU8H3GryH1WKlLc4x8g7fRV9mlZNOFCw2fHcLyt6WLUs8jYNV
/iqJkGViCIVJmWrOo/OJ/RzFm2TreZ3WTqGuZX0z98C4hOv+mgSJ6j6+AmJeGh4FAY1/SUTUPO8c
IJAlHRQ3qFoC3hds+AEtUkIrOHxlQJXqo7FM+NjsjO2eL4s6h1WDOAqh6nDJ3BtROVy+VrlKsMCM
Q3Qlt/lBKZKUBQtg9GDdYhwyZQ2GqeteBR7XC68pWzorIooVdsKfGnENSdG8waDzFtZ3pgJqAnge
g+Rv4oJaJq3d0Wigep39660ZG0chdp6rQhoWDyKS1HN+B6LNG6lFO6om/+xdO/peoZwGYUgSRMHm
OJPcoBarlVkjTtH39mVgFpzLg3u7TxHwbEd5lZpbhOyLqV8hUmxzhaT4M1dlBz9lQYypKommhVXF
37NVAAuNK6edHUhEytw1Drx++qZ5F95cDIO8OEOEn07WGxNSAbVQ8nJoSRyIvwM7PD/HuAmW2QTs
ed4giy8iXsexDyx8CzD3yuyaFiHnHGUVCLKWUJJtBuz8UrMARXUegPwRHhCzFz7FykMdPt3Xdkil
PEkypPI1IOu6IW20c+Y9rgrMWQ3GQlqyWHWxOIm2ZW5Y/MmMWog3DMpUkCe/SJT3DgVEgQ8TXZ4W
1us0A/rTZBXprncRsza81X+yjYSg3jfzUPDiXCSkGZEvYP700EInxPbs36llQrk8+SN/gi/TJxI4
lXwR2h6RDCIqBqpTKnz8eq6usioaCf0RUX5XKGqExWKWeZaQjEKsMdD40ASkBvoLyPDkneMn33vE
hLL6PsGc2c8S0KRopx3LbRc8dSl3UwJRL5jT6QnQ67CuMeEZVAd0qUAIliN51GueCg/dQJkObEkP
WKDiJKiFQAS5bsX+s6xjJO87WX8By8bHy3oHSKr7h41b0RkGVB/+kenO0jFlXOcuj0QAij2QsfvU
qJy+/e/aW5jaQGZxQhBfSQFFY0XZoK423LDDelmI6mNg0LSJRzpApDuR2wQ3xuSZFRlsEEgOApXX
rWEImbUT/S1JKA8HhRThYvCb1gI7ERB+Y/sfad2n2+tg21I4hKA876CvolLGeg4aoOOwzKZS1Fdm
fiYCGD8n/7ecMFBJRxJ2HJT8A9D4hWYh7rKvY08r28PjD6ePfckJ84FdkTJ+tse6LjnV+HBDNofq
2Zip28fKVfMcI/GaQ59Zet9dnx2kOQFw5+MqvptJHLsDrMJBgz3OKro6Ak/rZyJGU0KVnSHKLJOi
brexgX189w072Nbxn443XjFXGogV1wUlDx/mDtjPKzvwE4NiNNkFelTWm8uanrILYdq+Xuiv0Ihu
FOTiaQjjOn8z+kAo/9JhgHr+zn4Rwcb5qmw7m4o1BZlOxc2BgBkZ2qODZswIUxgrpvDyQMd6cUbx
spl68F1sUM3Cfryv+H8+MuAzK9DgXER3B4RLHEhoCKK+JUk+cQLXywFq2GuxOTBlokFqRvSuQup8
yi6BFuA/I5xVK+VubSiwz4shDQDmxjAsE3AmpsBBpeCnHKEazNse/Bf1qyTUtWaPB3SqLFP0JDjW
Uo5+uDfon96FPWUvmeCu0CM8wlnf7S2wBHU8SPDMJj0JkDHe5wMeZRlc5m+q03Komre9B4wkIEnK
LFvk24eX6Oh3ioIETR6rVlMMr2eZhMb4a9zwQNZm58h11y8sP1BAdyJe7zZLDVxh4yW++HjzLEvK
I2B9VoO980bHdWZ6OsrcMirEZUnmilj3uaxsRQQaoGJXmrx6eBfRvPIwbIZDAPAW4emWigj2tUud
TfrVkp3LOa/eeAhzphuf7xDqRX8hxbz7QQr0ZwYQXgHOspdaZFmYMN8xjdGOelFhcOSfeEnaX3kQ
IiremOpd3UHf1a+IprWfctSllTBAQhW8Fg0F9DDp1mn4b9qsE9TYhFzEofsHWEQRyMFm9iQRonTr
K0i72eySD3goCR7rpyI7EfNVdHGHgqh5tWpAfPp1jEHH9fIf2nxp2hpXzi3uqwxtaBHr7FgHTEtx
3AlutxtaLQT0oPMv46QvR1qRZvNaloMIeeH8l0Yk1xkd5zh3GEKzyqcCxSvhCJfxrY3EaewkUOcd
S8axFl9AlbWp26YXCwPkNJeGwG8oVGPlPBMAJwjirmoElP+w68yv7aEAmR3jUytDaFkZgGYtQDTB
kBYC9RYM/TeIcRmPxnXDIhRY63CO3BSnfKcJ04fpXrVna4OydTlz0kSPOcGJ3MOV5/tHStKNiSSc
NXakCQs71p4MEhl5HkmoDTRRF+Vgl6rnDxDFJqc3jOxzlzIxhZkSZVP4iwFPb8LMQYPL9Z6XUx8P
Q1OJ5M0uxjWn7XiDVQ+kDl1PXOTCxeABdFGvAt5WDM1+KCnPfHwkjfmRQpoPGxwuT6TLPLmF4lQ6
NTdoKFnvYfOnb0lwwExYSIIjaySFoyMq5PaMHa7u0/PwqTqH8hJFSyAbN6rkqAyCh/tXJZyS+cqs
XGsAGaWXnRLsXuDjE6E4O+NAKThICmRidZtPtpSKxXh8B9FS4nN9OfltKZFhlaKVaq29Wds2zEFC
W3ftgc6OaK/YCNbLLE4RXgHdQHp0YpMYkihFU9R1TuUnUGkQDQDjWgnIX9yUXKRkN1gl0k7lszS6
Bz7HBjiNOta8MuzTaohawAQgPZETfUfwX8xuiOGWlgjRYbVOUUuj3QcDpJxwqaOVFShosGyRIN3f
VyfRRdycpiPBEk8ShCK5YFu4yWVq5shizuwDh12lGclJvi9RrJu/DPENDhWE5dWSAGCE5/PHRwbs
cCkjHDVqgbq507vTPec4UDf8KZ1yGCjN68cmh/gX90Ms0F4ZrveU7P7XUXEh1jwFrrs4EIZ48249
DL4/kZ/x1ZSvTx2bdtwisv5C8IhflthlvvLdJk4qP60BXCl21Iia3Pz43WD5K7L2FwEUd+qFDYy4
8DxPnuFy53Grtr/bQeeDKbK1RW2AF22J6EAkJw38jwjfm4Lq0MDSLrc67Kv4QD0J2XQuuvp5rTs+
BJWXl8cmtLPs8XdsjVbMqil3QcUWZIvO+cvtRIZpfGMaetMWFh04hEHrcDy4eGn2BNQw5b5eK8vO
0Lb4BIyNuCwYJ26O2WqRwa+f2K4NMIRUCMrS4TcTt5v1jjmYtockLuvOpcMeBn8n5KJR9D2jxspz
C36PpvkvZO7dBLGbgvbhUOVC6uwkopkOJI8AjdB/rRr3Ip1VsCHnxeepjRTkhrQekPupcXwLi6qU
BJIhE+isCP0orv6TQH/VB9e5SAULJyRZHp/8Rm+eAvOVwS0121teYcd3w/Ri7G8Q9g8+hQSlZHSq
FmSnTB9aXKuDCinNB0CRSueSn3nV0+dyt+ABabTj2cxnpGe8edFnLD6N37hq9p/2EeOq084hGuqN
AYu3rRP8NxXbG34LGomQ2U45YCWX6zoxjJglLAVqV09Zh9YBuWcL4JSyIBGULUggE6N9Sf98jtIb
YF1YVB0wGDD0veKEckXARVgT+urBlRMe4JUhc9o7Gzl5goOBMPEqbb0KUPyJ3IaC7UNVrmEZUeYY
NHTDwQyfJKeJCHirrp0+aOYb0hIcSO733noJsXUJwKODSxx5wV5iR3jzejWFOiQ1tq90fLsHYu5t
wGeJfr7837cEcQGv609jGYfbZgvtQEObfNjk8V1dPdTg22irbT4VPGz28bVZmPtI4S8jSiYGhrgZ
11L5dzczroOYu5DTItpdpfyyTyBt6j11uCA8vJqu3K82kk2ytWE8jcMUqfdfUBeeJo/Dry1soJSo
VIZDg2RyskPgBHEFHe38Je3bP7SRekLKNSUvosWqopeBiAeaCZSZ6x5BivVQU32pzsKcNAy4wsMU
6fhpP+AteNInIyGmyAYwbKL5t3+7DOySG/dsgy7PjxxPsQkjkp5FYL3O1PqOMf64kHOSnp9AjsRO
GNK6cpkGvsewEplXkgrBozQzMv/rYSQqP8CNYasvhU5ghM9FpwEuNIFdL9Mg6Wg/3wi5+Bfy9jHU
W4QFKbtntGcQVSN5GTmjfM+shtI6dNdleen1XsKfMlvF+c+1hfanZWKv5qr0gRUVccteNLTBC/uc
qAjO3vOQs5l0JayNV59408VwWQcTVn4ZAzfSeYVKacbzg92nTpRqOe9OZetSDAl8Uwb0NnjWZPu1
eRco9UOLW0U1wZExiC7TLO4QfNM12ppaIvrTJaJQqKbxFfe3SJDhKONWtga0hJiOcCps668rfKnc
24jXd5dEWsWyxHUbeiM1AF+N8IcaSxKD6HaDCsuN/lIKErZ2/JPmm+wwlRPb0Q5Tp0aaG3s0FmyP
h0PXtzTj9O5G9Oj9/2LmkE+igW/0s788S4DygDMDltS8/ZnVNzL+H/9SMVc+J74+FfBTRHwioKMz
OiAHZr/kwwd66CB44uAP9ZdH5c29YpBLwnMdeYFr5do+Avx8WZx38XqOC0N93uFYVjz4jCnBNlgi
rLPCdI/oh+MWiFTqY3BfOEZgsEUlmCsYQAi7NYT0/dHqvdCDN64fIt3mJ7PmzQEpFsrc2orvPD6r
64+xqou94eYhjKzu6VHvw+IfrN7q/vYtszzxnL2x9vNa0Tkvib9QYU97s1JhmrgYgW6zyqsYn0fx
50Qc4mtMha2boZ1VvpEY+ou2J8Zz6bqVRwtaPTtmxUACrsz+YiYIgRnshbeh6NHmqHSZbiXGP3Nn
Hsx3T/nJZGa5JPmHAHgvnyIS2CgIRR9/bYcFKF5JsJs9qsAker95+7h2cmZsmfh2CpG2Y+w6H4DM
sU2gY7OZzBG5r5C+GYwnGJ6VkKbZbUaTTNK98DseBNmobHw/pcoZKgvfADUD+FghBBK0mDdgvXP4
XUg2OYbfpFf8NfAZYuATc/gF17oFpNW+XtVLv0Xkl7GQoHyFsdFFaBWCCCNEd5ixQAdY3KWWGR0x
CikYLKSWZqwlsThHZ7l5t4miNiS/88CmS52Y0oLadiBllCWtfZEVPhTqb/tmYVDjmHufmU9mKdOD
tfFGcLvrAfIiOgoXcD0jG7vQM+qUgjVn+DPnd0wPXw7cJ/PdtIQZkxUoE5E2rTR9/vCdDsBBnWY2
KthlMQEuATL7sJV0bRt9Rw2OcCGlcdVG5/iDwd3ciVScNZxXC/SKmv6Vq5BkyrT62qvPrY9o/FUN
GHIfxTcLaWq+RE6sjuriN2o0qBmH/2CFF9P2idb88QYzD9yw3fP54WEv5HTz1DKANPyXy1QlSx9a
DaQPqQZnPWnviSJwWNjIZXPfBh3pBbrdh9KDV0HyEqy/eBqjwwGrfSgSLOhrdUEbocfLHbNoNPwx
LftMwcLJWUA+2OC4BVfJi46sZ4C23VjO4pA4S1L+AW6yQncbssJC3NqTB0s392tvXmVq8WrlOpvn
JAESqy1lrycVYpWPxgjrC4zcwEMmBNnaGCs63Gykxb89D9iYkLzm9J2JEXp8qlT9qZ1B9cyUsdZx
Bp883C2LW1CxqY4yU59qJvlkGQorQ9nrWj2MEVYNmY3dvlIqp5ULKuT6Qu15sVA8JbYzO7eauaIQ
y8z5kOQy06QIEYfAiD/qwDgQw3PwQxqxFZTfw+nD0u3FPHe0KGv67jqK3E8tMAQyCIz+bZYHQnbc
fbOaxO4xZXUw94A20i+zZwhjuNXIn5E7MSGz8VCUDj3ZbYI0Y7XGblenguP2prGnUvERNjdgyMnC
MKbu94WdU5FuJT+8l4WykbEZ0h8h97OOashmwNd09nGHliW8UHoxhKSiE3g7CnkNYTwd9l9aUOo6
PeA7TW/WGRF0Jw8bZn2v1KYytnjXwWB1K0QfcFZric4WLZx7jY7GUrcF5h3es+ckXznQauXqaxfS
bHI5LDCKeQSyKgyYgZgQla5eVspMRkTfZaIBvq1+dFSqwBcjja+EveFJFFFt2Y+7GEoABlAZUSj6
T4GtGV6zqNPgQHabCZLNPsPFMCcSa0HuJhxzWpUi15yCJNDSXsm4paABxyxFGwr2xWdvIQ4p7Wkr
hvXG8bVSjsPBh3ttp8v3IqQ+cOwVWbdy/2TI9ce17RRBLTfXf/dw+YrtzskngN0inBFDHYNi7E+3
5cnlxcgip23aQxXAij9jwR5jn0SO47tHNRUFXvvEgfP9uVNFg1atKd40B7BNWeAaz+btulSfvXgZ
n6X7Eq/Epq/7s4FdAQYWnqH8buld8WqSxT4eFv2da37iULGU/PCNGn55Tj/aeBZJeQuFSDHOqQA9
enCPLbPdzE2XjLQk+yuBtEdwV1wqsUkSkwwQwOg2BHRgljqv6H4PknqK7CWQXuP5Ts5I341AEpMi
+o2UZN+MtYl3AzOO/QE7Nqm44BszbtSp+R++OC0HwSnsYALYUTwMkXhxdoKHZsB8tXTCtGYBp4RB
BgY4PyWQgM1ShXbRrQ6ehJz0kzmGVYVhQAe4gSUGLbExkYjnd8ZzvFeK5WF3BQP/JnTtK73SjVjP
pUe2u7JULCn2bMdU+ZVdhSZ593CJSWxI5alnzTTZ3dVkaFz7LZ2u+o02D9GNNVGPSvVH7BRPkT6B
Hab1nuEz6GoHRVfahs/I+QjGyyvMiNALQecpRg7k68EC2O4VfEZcSi8LZyhnIpGV2wzkugmJwlpC
3WA6ML27pbWCo0MxV8z2Pd2jZs95MDvb0Dbzu4TL389jNVPhVhHCiPyXXoOava6mGoEAoEuEKUrU
imCnnspGlE6eC5afahbHoHME0wHjDTPo6Ka8S5kG0pZJF9Y6YrseVWdkKLA4PXcYHbaDjWDcrkn5
1p3hk1Gm7O+yxmGno0E0QiPmRY1SucAKc9nuNI1YeAEupqpugQJryir3we03uOIM0Bcw7HGczvNx
CRxpJl/i7oJYYJt4mqqekbfQ3JmWs4VE6gP4d6y4kI8eN8jppbT4G5k5Oxwl0KTGfn9GCT3reSNr
i5VKZChyhIYMPJqMwrZ/MdM3wIKKy+mhxvBfQQNyVU5T8xx4+dLVpZ74JhX71AhiWqK4hI9wF29o
QHG+PIKumfUJWw4UDEQ7WR/G4+TL1HFEcaQ/W7ub9LY22jg72dx7cZyZKPTB7Z9m+wvgkcuPYHZg
HkzpzG+FkoL8PM662+Ug0ZvC1u3eypes28aN6E3rdwTjQALND6zqS8UYS9f7zU04A49GVB3zSq9d
ggo3bhRUZ22MEIFOf1Q3PtWwF1HYY4kTJkF3ejjP5xLAP92sJm696cgGnZFzHlSmyxLDijBu4Q2d
lVBpbUiY68/kfLwDT7pvMafw80u3OPaMQHwibbWe+uYKxlcNql9IGQ761/okYn6gW2Sd/jm/vQhY
q0LvzeY5l87gUJHe3qPabQWQookNH7KANocsmNNsp1X1Y6A821PQHqdJsD5vrLrW0tc+d1YQntbM
at0dtfvA7IjVqN7Ichbby6xWwTtlnNP8gxOMZsod1mzjsq4pYtRWdwd5Jh/672j0wNgfaC8yDsms
dgIWdRrpuBv1ZdVFJmsQiT+/vJ9Y/B3JiFFIz8y+TZs7V2kKXvbf0BJnm/+GfNDPiqFniL5Z5r0g
Y9fOWVP57bXRMgPUTNmA1ey1xeM1UbyNKqXp5fHpinwVKmpH9kmDxMNAtjGvPQGJGhl/wwmXXpgd
AzyplZKgIVkwUVL1BzJwQjbKdrF6IbbUBkzVeoH5fBQbjptVIrqqxiG6nXfbgJM880MISm6gYgci
O2jcDGwER0cMh/8kSAYa85LObKQNAclezu0YEVGtGEN6/+dWzVgAegn8o5+DxJQHsKkzSLX1x3cp
wk4QedUKK+3HYf5/Vm+fQnS2Ib+ZkGoYR3VaCu14sLv0bN1VswchjpV/lwMC7vZENFhzdy+/+SOS
ouhGI+paKVaOuZh6NlC4CmlwnpdClnwri23ifbaHIep9JeYVMf5CNPYdI30GeK2p0HbWPrNZPdEG
MliLzIqfOz+YWbw0gZy6NfbEjq82oghyT9thAPQznp89cS3j2paVs60G35PbejI9+5EXc+dcheO6
UZzAkamekGAMuQNIa0WJ+w6IteYxzQJHuBJSgdIDyezR8Xjj0zDmcF/c3FFjCToxuuH/XWzabN7J
m48tIedTkT9h3RBcyAwOstTKSXe0Nmukio0OIAiYVOGmVbYUNeMeq7ASORmCp+kZOrRcA0yzoMhR
c43kKT6WFKHY/Nt/qgR4gG3aqd/dpRd7pjbAHyDKz+E89x3R5A73+VvFvnet+y0jN2gEZxboGqef
u5eJP35IgtKbSLC4LGrzBQ0rlHoN2DuXq8xc8FyOWXqpi6o8En5bJSFhiRA613ivsfcF9Nf5hEdC
v0Ga/lLFuhSPWdiTqT9fNExtkxJb1w+hGguSkhhu6f1+FjuYPk/KcQpmk4S0h4FwmE+p+VcemGYT
S0X8CQIeJtJ0i8hBTaAZ9GDEcnuD55lyOuvpIrU/BOcg0SdEIEZJsV/aNwEGHEnUCKfilA5D2UtE
AGYkEZoLGKqMfci7xn4iwoyd77VTCVlg2jgZKwl/tlHjK4dSiPcvyIzmMGkXHztvVw5S+6q3QJGY
HxpXkBMhyZ7LXrx3QQMgTkdUgkwYgSrabf8xpIeRa+3kbLzeulI5nyy8O/bTKxS3wxVgNCioJxLM
LiVubP6rB+n0P4RQZ8f8VDRARQQ3u1a+V9aiPQuAzjwhVtnEPV2Hmzxd8uIv3G4NciAKfmDbznVi
SaP9SXHtiJfrCuzYYoL/bDM7kmYWRtBbN1yofKBMxCRASENz/hfv4PMj9GE8SjiyZ5U169g4uzJo
37rId9K93uqJLnEm5MeI2tFyNgCAFCil1WWGm0hh4etJKTlgTQmndBVScpIdi34sdjKsWLKMW9b5
dwuuxinpQiQ//NrujYbptZvFllCFwibAZy5fWtmkakrYG2rGyZTQDnp0DvLcoiNEQUBW6DdQTXUT
tMYsC95FZ929ZtcnpSH8qI+So7wl7Njxi7kWMR+o3HyZA6NaJOfpeoaSTulC9JLSf9dLnbJ2QbJb
eLco/zzHQo1cr/V/xHvMbZRfJqIK1K2/u+fi7NHMY6i5D2rMk4BuXTLXo/oeWYYq/ALCYM4yey0n
8NZmPjfd06pUmuGCqPBi6vqEJ8hD39QFaORzzqQZOVvxf+qg9CUX2MjnlhOXsCb3qzbdQ/CAvotK
9XLQXL6eiY0thc+JJkgOy3w0Vpnw6QDqk+E4BJGZJ1vJCtnqigWs6KI7otyvHjeqn9XB+X0+OJ5u
ZKm1de1QX6kGAYUiBp3PL1GOphlopJT4Y6ILJgIceSYac/QY2k/s8x6sbTwLdLgndD1y1Ll92a0f
XHBsXkaTm6Tnrz6WlStoeEm+u1MoGUw6mkWHBcnaq1JM5a7YKBPxepb+Y8ROZt8flIWjI2oB4yLb
1uQ0yyQmXAWzQ83yGEkZjWDoYMjn79vu3GpPZjvTsfpiCfJrkWRmgqos/2WHHlBHaHEWe6IwKa4F
R6He+K/3hGPj67ReDDq0uD7GrKTrJIV0ry9sUkY8zlMgoy8O7YoK5qysL4Wdg+apv9QbComDZy3e
3BoONVeYwq0UHTk3oFfVdffQFGPqyBvmser15+lC9Viq5sVj8KL5VOuuvVi/S/9CAE/QNZG4oNPK
ETped8dbiHWyhR9+rQ46rPN/qEhW/f53VPLfcqJGkLgaN4w6KF5Db7pY2+kzZ/8IxTpgeSF9sO+j
PvJhk8hD3vzmCWOFp5iSEOBWdpuN+zhhLug6oQ5soy2HLKeLCUN7oaLenQKTcABmpcijsL7IWTHT
Wx6pqx/TxoHZvjffd/gMslngEoTNK5ZBUhhuA4F2Ij9P/jeJ6KTFz7A4Jz/JjwBIvL5XJzF/nA/d
5AhihgcLU09LN+pDhmDcp6QbPic+ea2YLcuMVavl9LQ8rkohczsIGMGpWkUPP/ucOctbakR7zvw4
xnEv+ZQtcdJh3eVjBEmMXje/Msmi7+9k6Aml0lbcDACDpwLL6rqgm/uk1cctlXE6xtMONk4c+yJN
FOTKF9hnliGLOm1mcEOyhSAnvriJacS42U+zqauIR/mw/ajMfNA+AEOtzQJBe7t4yycLiKRnWGtk
QsUSdsTevFB9s1KQkI078ahdCqyamgXqQSoHRBQGk9E8U/g93nl3YSzpDv4q/RQGDuZg4fKD/LLW
dZ/et2pGfO/w5gnksFVzv1EjQRnEOobxz1HSUf7DmRYbQT8Cw2cSLmKiH0akH89cAWFBAkshiRDp
W8x2P7vQUMFE42yvnIy26FvZNngocZHeBOrW7ceMoayiHASrqgMZW/fCnji1ZSC1jIGETBHJGaPP
i3M6SvselMoDVsYehXj24Y6iHXBNvM2NXrcQV/A4dAu7FKy8ViKV9uEbYFYYz9XcpLLwrjddpVWG
WfK8hPJIY1ZVVPGcsaXu/qyPnk/uy6uTZfEk2ZhuVpsfd/q4SfSWPbvmeUHluVwh67HEvwuOS2Rf
nJB/jkEODJoNB03IXflDkMHq9OS8bmsFtGiP4zIKD+dOppRg5bm4sCJot3Ts47Mlu3nV+jScIDjO
odmh5LzlLa0IGS3uhnlNtG5xKKwo8CLwOIAQi9+wQGLc1OHd46dSYZueprJ8y+uaKbiwMnCkoFh8
t3wqQZ+qCylXQZmORB6Y8BwqZzRxsB6Cp1pSM9xZfjF51A3mNdPgCBgl7cBS7DFKU66AXhwiU2oW
WYKGwZ7CLF5SL5YFe59BCnmP0e8Fb+qWMLQ53inBnpdaVAxYwNH41LLBVM5tjGoO72CIuV7RVvBj
Jp6O/hPE/XlhNjNIctirsxjs+2HTLZaidSahnz3xS7HHlBgHeS+Wa3lQiyw01uqVjxh9eAhGH40y
I21dCGqOGrHTn4G9fPaKNxbB0wgY2WMvZ185D3duq1WMi3keyVYytXhMtJFyy26G+IS7buWPgh67
+km/rXHV/GfJ3zpHCI34Rzmk3mqgDXstSErs2SPkIOGt40GRCj06K7gsFdniSuJeBlKuZsmjCS3l
TnEk5RiK/J3dXOT0Xqvd+3sO3EUav96ruK/a1Y+GvkQQ7pUduH0OBCxMT6sDRyR9I9ek3YyLnu6R
xUV8G11N3x3XQoUtqoBiothuCrwot/izAMFVCGDqAoFAvEVWod52+T0IWtKwNp6kZCSm0bHE7RYI
MtYpeUSeiIfiPlg0Z0y8nQF1H1jXWIH3+gGROt0R3TndGLxQLXzX+1nxew74uGkRojbs9WYyDWZT
99OeyP26zpY9KmUjGEGR2F+0+FVuoDmdnBSGDo0Bfjfjre2qBOXEmM7NFEfUvpr4uKdmCkV1dpSN
AzrkQrmiZs+s3s28e+oBNqsr3FC+E5ns+9az7619+gZXeF0IOpp92Er1XdHk7hsSZw74H26YCvLQ
fGY0E6vBG8u6EgoWUxHD/92wu5ySLSdrckqFYb/8mlsSm26DMX3XOZmSTLlf0UfyV0SoKuu9UuKe
Zwz4B/thynxUsntqqStfHx8yb/OFA7qawKB3a+auqh6TzIlVUMNjKV9kKwtHkrdBYDPY6EvJAZ/S
5j0Uc1FxNZ4bsmawS0rUKFAjhBZVIQGb3kERSq8FTDuNsJ1VnRsGd2lRTpBgobpftElIgxpOQXSl
vz8bsWaa474fp18ZtGDA2ejtk2TmsOqr0UK/hbYA6GuldNoTcpXhPM5vwFEAyen7bftVSNIpZkUh
2Q2MHCgbPRuWmXUwFRW4rx1mfVAHazgC6M7qskwrou6lRfgPB5HCM2nDb1Ab6IpjOKEUbLoTfRSX
RTxa2LU18vhKvwkglWAlGCKJ4ABjs8/DIh7t6pyXZdyiTnMEUcjQkLNqaLbq+/etWFqsbUirsKsw
sCt7PiiPuoMiCxmo9NuIAkRInOOX+HajDukAfR+fA3dMd431Mc+SI7uJzXrIGkCcBqR+pRDlvnFi
haC9S2WBpkYX7mdJeWIXhvuofEPTxHwTE2EgLPRaKE06W9oyCYckvgldSfr/MpaHVXfvN612w4go
oBPy53jLAo69qCJ51V9EoO0R0rEB0i6Q4EByyTFixXwcuNI2iiXHL1krcm1HGsNXXCCD+LzMBWar
wvhb8cl87Dhfyy7CUeO+kljHmK78vsrFxeF2tBV88qu7+ogusMMW6kVwtBD4F+hqSvjByHR20Pmd
AmQd1qF+r2vs9gznSCsoQ8Icgu+V8ySu/1z33/rpsbAo+EfzjYVpy378230BxeWOpPR2b6hO+bqY
+Q7L6i7L4DAbM6oq5ng79efEm6iEDWP93CpcqmQMmG+sdUPNASDDhTn1Ow/8bRZEqYhE++MB9tfq
A0oPvqy8ym6kcAsDoAsfD2NAIplCaQdBrw6WIAOhlKu+joVMIAKKAxVyrg9gK6PsVjZSQeP3jLjN
tNcJ/K2PkRGUALFJZfcTaOgOoPrVdKNVuwZBVUPO/vua81F1TBZkyEoTfpsu/qJWKLk+25yo9f12
ZazEeFz0QjEiQF/YeZaic5CpKdSWLNb7zE8cs4HTomday2RtE2Uv/kDZ1ylUOlaUMV0KHAWOKbqB
SRyI1oVDu0RYLUOnHMj2Se7nDffJYCjWiwmkacOA0BKNNqNwxIlS156B+kFvc1GdvGIm9UfbyQbO
8ek5SypxXcH1PepjayMLDjOQTjzULGJvQ6juBXKWy7kDKfdc46tM9/yAOUWLY3iMtgJWYGnTjxAl
LAryjCKsQWW+ERgBimuZMzHZxbGwIZ+IMPLsyTVwdBbq3oqpeDj6JOco1UT+AZc3QNRtgtCWRJi3
/1AwS5UMXzffbg9xDuZSjXfGVBHzQJJFvahr6cEgtjJrT3NMGa+K3Yt9Z6Gk8kbW8DbRZ4OTIsfS
2armdjqa+PYXh8Q4xzjh7xILUmcPKHB5/F89wRMb+jX2lLZYKzoZeoY024DgCXp2oJjrcYf+noMm
O/MSAdb9B/Cli8MS/yIFGDCdq4E2MrxSEiKLGTbMQNNOUT3vytzHHmsq8YM1JV4cqCnv1nyM7huM
2i2t+doaOC1Rjv7OS52zfV5mJebPpB63RjO0OHpTRCiQR+WQVA8na9TjP3t8wfIs2E6poMbScvET
aDMBxH4SySeXGYjwgBxdCh5ViDn2+Qlvoei7iGcHPjIvGVsJcroZE/RkCOaOQ3BTnVE/MZsykK4Y
aRQOByc9RmZDY+vlE98rxYSi5u3qVcy4U4aeYCJJNXkzc95uegZEP0AQI+Qn5SQvkV6zbyUBpDt2
6SFGwz9v8RGP//fD3k5dJnSdqIoLGm25dLD6u95QpCCDgVghw2iWUktBl47q59eqB9OoA9TYYyaM
qVI4gcMHtrcFDRrV1ATpjEvz3NEHNpFbcaavGZy7S7WlukYQ8eZDSxueh+89i64Iy1qSrGjuFua+
6q9Wj+BpDpttVJoH/FhPOMxhAFHIyquF1pbXjxdRaxp6ZHZhow2Nsx0J2/10x0A6PK45aga95V5K
eEjVnGc3l75wekGf8PPk9O8W5e1vBmc8nE7elWDXFNDno0c3jAUrfWq/wYgMyrtN/UcdnGYR0UNn
IWrjm1PrnIbc/q1t4xdFltv+hx535PrIxCV8s40N2BTBEVlPtzzcMTCQ9t/xhplOB8y9Ed5MVKXr
WutVMax5gFFVpSwS1c+odzn4hzHjjgpvBPGq68q4i8//31D9awaia43sJAf99q3Ztp8s630sMORj
KNJ5ChlirJ5HStHrGZc+9m6RCzoZsuKgef0XA7TH5jfwOxJAwZFi8wSfZiAQfBk+8n28Qbcm8mZN
I5KnKyvBqck0WRtalqI6k85CQ8bB/fg0IBxU4j6ueRk7j1X3gPIwBLeEt8MgitCdoyNCiyH+HP+H
xyIowiJ4k2XiZEOJDF79WVCWm17omFsSlUoeCZBxq9Gr0aYR4whsUzZKQ4oBplMfzzAI0O+7cofO
iYB5BsUjmAdnLA3ULY0AWXYGZ/fJh081OJnZI3EdwOMhfDq5NdVQbhTT7qDIUM7zwOqukyHRyADy
wVduB+dRumGbbU/hdqyGou4Ukds5PnX75PJ9jB9cbSopLAmpke6Rpk5MkeIvxAUDUFzHqt+SXm4n
uGnZkaAHSh+NXo3sq/Z5cfcBR/1QYphhNeFJ+gJpdKGiT80uuVIn46sh0gvcLpCcMZiIo2J9FZBv
aTitgYPn3G4ZnSWGOTmwjjUZVLeLFc0TKDfKkDUeTNOnGTK3eszTC71vVpZJyyWmK/ejZeSw6m66
3xyyBSz9QrN8XuItzqpciNlFYp8dN0zaIxpg2In47VXuKteCuKBVugoECgdq8WnqL5QSesFXV5jQ
nsH4pvRpudWZGf2JKee00mIwp9Tt3vtEaF9Svfdg+w7gpLaEjf5gxpV2tCoWPA7+yWD0//uMJJh2
6yTpqlbfIy16lg11CYMQ+yBe6d2UYqFR9nUkST39mUWJQK7zNKdhumf3QeRSlvs417RmZJDamBUz
3D0arDr1g0KsTltWGCYY+FRBgX3m7ekcE4l82y2IlM9VJJVgvxXv5VpHuMGwwtaBF5dORNU+Vg4L
YgPV7DKL7q1rxeYdI/P2/dvBfM4+0N9ycPmOTvspR3wTEOTJtws4NbVzWnTwScASayee4WuubvOF
DrE0TzXFXEhorCeF7BTvOtXOjJ981tF2M8+bElqVlx4QbeBT2Hc8G2uBL2ysSfxg82yOe3ONBLQs
sI/qCwR95j3LNcOmSx9HKQx/+pgHj1/FQ0Ctw8gq7WCk/G2W85oYMsI0JuhJJQqAdr6og6GRhise
Om4+Nald5RQYDJfoN3BQ9KAJv3K3fpgTPEDX7ykffGL2vPdp0CsLx1hIm7HRsyygDHcZpl6bz0t4
4Kk+n33b8DQQXrBlIMiw8NpcSH7Pl9rbEkdJY6Qb3hu/EnilYhZZAPy9TH/8xKGIC51rv8ARG3jM
Kee6Y3hgVwoO+k6PaZr4R/eK5zW4NIWGgw97FQaUqnNp4wGksDijkbUuDnXwdN7f4kP9wxEgXZvP
zWFYhGhYXeayeV4Ga71uGjp36qWeETnsk8uSbW/cBg4q6NAkRKCH7xBUKhgNe3MPmbmhyyyBE+CF
aGuMwAIPFq/ZuPuCttz53i2KeRccBfJF/+8a7ko5b5VqlSJoeTLDj39dzesrrXYNUaCgsBJ9LvIp
CScjHhGMcL0IOZ3wnMDofUcRVKOA27obmEPOYeMDsNk2sYrKS0YTz3piUd/geQcXAp5wTsvb5sIW
mXveIK6kLEHfKuQxR+Phe/5RkPK+sL+CyiPLtTnvswvTNg52xoSlUflOrx+zdy80yLKQ7DTGMppS
Y/aN9c4HtvvZE/jY/8z6FfgDOE8LvbU/J52fL9GcpGm1h/n4pCphF1V5HPhMlrzj/n8N0+EPTB48
XuFB/gNYbOs2nU0b3UmeJ2M+52r3jX6Epsqs3XtwAkgVFTtL44K6RFyORX4NBXCiHr+/8Q88QnrR
TZxwQBpi7Ii8V8FEpCmvlM3v7UtDimTPXVq0Mch2ibh3x0Gd26OFlfJdvOQYpp/ADv527BqrmEms
zD41f7dJsId4cGCHcQSvF+YKHd5Z2iHLh+ls/5BeYRaV40UBV/pyosAYm83LPo7MbkioNWWGooUX
bBkbA0/cPZStTKJbTHMmMHsIJC+p4NZB+1IsgpMmrtPAO53HcHFsXocayKQj2rpjFW2G7n+Dfuyh
ZqxwNJY7VGbDoCEdjBXvGiY7nD/oYtkqR/wPRR7XsMAnCEYvRNTmcH9ShKME14xFCy3c9x5pYncC
tTFQrhWpteG9RTpVZ6A1/wNp8adHa/Pa/aVV7umYvwtmIwjGJ3QOpMXVBNGR00KxLgSLqaw74YwE
kpmSvIBK07rWIOSF+rN6YgeF43v3SGNImk3OdosDCPuclvQdJCQGWqqV46bDwmL0lRNgL4CRYuyt
WoXR8TgjwO3mBWdW3uz8Fcq0yFOfOUsYK9FiWLfq/Q1T89KfMW4N8HPVPwpf7Ek62e/m/PuppFyg
GB3Gr4JkDgjW+RP85gqdnoZUOH1nfUHa91TpnC6/9ahjcp2E+3RdV6eXA+u7Z18zHdkw+K+cROHH
740sMCiADV/MKFdu0nYQhKeY0akyw9m97mY8fzWPib82sopUTIXDvhpl4y4827H3ZJkePLYxkZeY
nJyIA1NNyi9xAlc4MAGVQodwxpIKbkNAmvt6SIsd162yul+xZ81oIMbjFfjR21SJZB49+4V22SAA
+Gch+Fkl1NH7YjL842WlhoozqBmbrY4UCAz1vXPybVC5RfH8k5jYThrr5gGff4v0az4EYRYqeSKe
IMEwQixxi64V/uXIIqd4hc33fnxU/gU+rc88lYOOf56hATEzBoIpAq1CzxSvAue7IZgFi0SLaJ8v
mzVewVM5QqBN/zf96Tbsly1qjk7okLC23OXpvDa7W5YUdrfSQGmbl4gTtxBGBTqXe/YfcA4v2kfm
uy1cSQhuYKEogcsFuEUaJ/cEhKMUwiQ3S/Gpzh7WPPJzAap6nLGNpC65mKsyp8aEOfI2pptEWhfu
8S1K7Ws8v3PM74HzsCqr+4S3f7QCsFBHFrdouydOc+TlWw1hq9fb0GVqWz5LK1nC/5iAz6bj2BHD
sgGs+e8Fx9ZrlyimukjhK3ifZTjP6i/Exf8xemPF2LIoRwVsbu/WJxLL5H1xodm4iZIMDCm8L3X2
enWE9l0z+Sss1sBO6tHte7FLOvz6X6cGE6REZrNjmeZAx3ifzd9WfyrRmucCgRWvPfiW7hxMas2G
3iJgTKf/tC/cC8al54JsrBYvTmpNN6YnIgYL2HN0jGtblGLu6O9yEBycB/azEf14wCyT1LtEXuCI
QPpPofptUxvlykURDW+Dfp7RD9NKg5wPoZovZRvcy7XRjCBDN/4sRYrJ8BPcvENjJCwkj4zoc/kp
Ut8iXivNPCCFOW69pEPSjc3ZBu3bHOQBNZOAGZ+0Wqz1A3Caab6GfW2EXTfVmJMGIiTQNBDdnBNB
gNrgu1UEP6n7D+ltrOmjBQNG8cD6PCIrHIYWHlHqNf0lJN8yJ6o7xf9YM9o02vgdro4yeoF08lSJ
s/lLv9ZCqroN3AidHevN6TL8BaHFvnn1FXMMZioRoyAyNyLm/AJ4HXUvKliaxsyavEOKmdfDBZNP
VcVLwhAVmSlDvH0kjL2UEMPa/Ci+a1GZ4khpeGH6sAI5CIUYoyAIwfL0f36hRiIPdOIh/fdE5ih9
erAUXse+Em4p1A9S55vuw/TlQWe1Sx+YF7s7PS3NeKLLYVJtq2NAyH52L6OAunHPg8a87jJjL7vB
dGG8H81bgK+iirdXWfw44gwFXLFU2yLoGyud2KMfDXH1yeo95TjGBtEiuiT6X1/xNaI/x0WJSAyx
thlmwTvNgnN9TCANNUUghVq7ePqakPJ/LQQEZUOp0sg43cTHmk/r8ghb6jy34awQxVbe0Z7AAmEg
9AKjNbjrnvR3H4Il358wkIIMRzuvVJJl+EfNscDVoo46/4mX+ssXnmZlrbOrHqtiJ7c/SeXseFlF
nTTg5H2bJoIhaThApLEw3JXVFVhIwjVJ4O1zWToMKBYlVWgwmWoQzXrljK448pEdfy4cJ4v1gsW6
Q3eZuHFRlC3FMGwhVG3OMLK8g5pEaWZfD2iHsTXpvvwHCSgwUThVTxcfh9cnav+Y7qvz8+jZcCj/
H4CP+edlvIx70+p59dTraI78z4wkPSEW2MkPKpBbYAJ7/fqRb/UQy6vPC7Ui4CrRxymrQR2ois/Q
4vfpR32Lj5F5MelMfjq45yJPZRCbpKjzFYUz9AV5E2VQN5Mi/1F+CbjFnqKVrFRKjJO+O2bZn6rO
ch5k5dPRLZciskcxELGgpfUjbO6np89zfa8ADf02Bjboi4eEb4qlEr49zm4qv7qwW8EC9FxNzO7B
uzQsn8RgkdHyDkSyjNGnt+ylVIC2sUKjXM4ZctREo2a1PgZcAzj1bVp6n4E8GME9f0Y/DfuU0OVl
WhBnsbsmPycjXLlZ1ajH308/u9Ffhy7oQRxGKxK+YwdbO1DDhU8D/SivqEzSYo4EZyO975RIQDCB
TccfJVMDrCNeGyJoJk6PUkn4Z0cQvDn/TOn13Bwnb6/zEht2U86lI4UN/yAo+24D6amHUWswIGWU
QPpI01D8guE13wfBtRFedtqrmw9b59qlDbRS14pWoNLJfmC1JG1H6qZMoWZ1PNlO0ce2ZvPNWA5j
lWvpOHZ4HTDGy0kAF/DXJoilA+nfBS6f1dARKvFQ48HUYqGYnks58Z+JzB1G93fBMJGZiQ0q5wIg
yvBH/8Hqv7OlMANasnI4qcR01+Q+/B8ovMGRbZi7JCHrn/JVykYdepK3DXiZQXC5koDimLLFlEHb
J5EqY7UGoGgFVqU4cJWLWMpvPOT7spMVqygCwUjLU5JocLrPQrLIRqynRGxmskE/8oEkn91OT8jW
LwJa8yeSFP+t/g0c+C/ZVRt4kjVlX2X0jpFMPe20cheUjPdZYhbd2jWUO9Yi43o+Pq0hN3tVQZsd
GPHpd5mYagatmLKBdHHZQyBLTXpwU4KQKtCjU/7l5K56EuuWDCAKjXsxw8aK/I5+hM2uzrnsjyyE
6L5ufVkkO0Q5spJ9cojM766uT44FJFWtJ4Eu4433euaokuTCdK1DpR88BJOR8Tb1aG7dsIt3aVbW
YqvP2sKciN1916t6zmebFEw8BZ9LaUzX/fIsFFWV1NeL4M8SDnveHtusWDk6xKzqgIhxGh4sXOfv
FvTsfwj1dsfHxh46gu4B+yFqpZHJwYLohLH0vQdOw3DKqWwVkWm4zTvdDTTRkyZYljBj3uCJ8fGK
nR945w2kjOf7VvUWCcn3hZVD34J6i5Vf+xc8eHCFDX4WOi6FAH7PEkwkzUKH5NXyYl07CuXfW7Zd
rmS0JCQNWr/Mz4/dsErUTxJUawdZoENg14CMXghilFrbc8bSWsyUopOyT8SOyWZ8wqDJGhfEcLnn
2j5yxSYHThqW8tIl0YRnfnYpsgQS/mPeC63leMAyzKvXYE2gx4zc5B5fYGTvSVqfl/DXTYLTb7AR
cjTCyH4OUkbTzkgsRo2qj4wzI8k6QOudmSZ3hO6NosvuwRb6sMJyuNioF5eNJxKeWJxiRuf6T79Y
wnny8NSxaAgk+SnOFWXDK894JEmNsdL3uI57yM2d8wVI8Z3Huy0gpFSr1NypOcRzzMsb7FEIx9w5
A4yQ2B8EenAmdAHHGIFtBMPxcfZ9EBRChmItVbbaGYdBQjGn6DuVkoUzYKH8QLKnia+NlGn5L6P9
DmpparShWAQ8JoMDoYNv+d4MX6S8mOwUfbyTnAx2mS/eeEcB2USP/65A86xPd1LHkHWyXwo0NdTF
Biur9yOMcg4fMQbko3FfO392rI+tTiVH4m7AQnQNF/8uvQRmuwVfTKg5lDut58/rOTYiLNmZK/O2
TJJ2IQKuY9mDE6OB83GWnwp3KP0rRP8kRFkNoHWyqtBzQHMgl/6crX2CTpx78UOkuC45lrIUMyZi
LYucTPz3A1w/R0+w8D5a+qRTTIaPJuIgTrcEp5R/nB0q0AHhB0WvfjlYugJ+AUybEmvYlhNyWas6
OSc4Inabh0o9K2wgH86xEG1CHCDb3NXnhjBzCk+e6tk1mrjHwUC9fT6isJ8JRfXze0xK2P23lZn1
oQiXCJxD8Y/DARHmUrfhnXtL6ujkF629RbzfZTv5WqLTAtKMGjOZ+RWD+552qs7GMzR11SVD6Ije
EVAmMiSYIxNYfcHe7Z+BmSPGkghMyM12JXPjSxZKocfBzs6/kQT7TWo53oAuahzXxBrQPXdJ8KPq
hQj+dM+T8eSD0EpDdla6fisUSUuRGUxjQSUonKMQHoCqkYsfbuBF8RzxAiCnlqKGi5IoMriFQpcF
CThCPAdnjmFA9gV9qd0poqT577m1YkYPPT1YAImUB+v3JSt1bpMC6139UcCpfdpTpso8RhGFev1W
QvzkazVGO57Zx7e6GqtotnORPM4ttHdPVtGEAg7tuW5pwwGdsTs2CmwAYUkyNPrXAQOpEsHoIsY4
Uf2UopvKbAL9fCWQ3TIGzbo/RExjzTKFM5zwzT4ilr3CmN7LdVkdMwGSJs+LoZz5Efo1MiutcS/a
MduFU53W5ZOo3VJCgDbnPq41ZCTw82OfM7znSmg+ApgE1NjfnE1R7bB5wR4CGFV4xbEqvVZLV3iC
J6bsqfG2AqN1inMk367D5mhyKkFlmHJQoPD2aCloYQuMAcrqu8eqgEVB7EdfbH+HZDJSmkoBTNxR
D1k+p292QpknbU+lBBuSv6JtoYBsDc8fJw8fk5NkZToZMz+c8p2jrNQ9xTF6K2Ex7KSXvR45sAK2
Ts79nZe3XgS89pgXdKzYgSRMyYW/GrgQKxNMmG8BfBnPryFrgiyHDAHMU7MAwf1PJGeyo8MRQ0l0
xRycjB4CcBbG3sMjkDJHKYz6CbvDjQBLD0xuD6iFHsgzms55lmX4aIOtK1SLFCAy9AnA2CKBcL6o
th6XSKeCjN/YAWC8WeuqYdmQ+BCE/P/ZvbBoeBuyN/r8KYVAjTCvQVxaEQXCex1G16Myg+NeWj01
Ir2WQbMDOlTfowJWdqXElWQF4/Ccbs/fwz0fNMG9pJLoS6Qcu+crfXghIZ8QQ2jpkg5zx+TOW24y
EYdrhaWqj7U8XOYWP+FP+jCbwuUF1b1qRuR5rdtbSO6BtBMHN8G/FCrElR/fOFQg/Ojz2NYldk1E
g/uHrUsc5rP5vwwdR8Ud6NRiBzNlSUgDWLjyncLx6PKkbNSYECaIs9cn7vxMsiODvwcVijpu5lT/
++7lsnf3cEbYOAqN1HT01rFEzcLrv8kE7F0m2N+sICUITeZBcLIYZVC8s5VyR6rdRZ7zQByhYm0Y
xvg+8doFKXT9niL0EuH/hX+BpNH/Q2qybTz/k13Yl70ZfK3Fz79+bJT3bP23NMA00TPVk7hIOtcz
ipTibrQW43XQ1por4UgSgv8G7dHapboNNI2LazbpGw65X8OuF6A6/jFkyn4dm68g6eXRk27H+Zzc
QFhACYeFx7W6bKJ0H7fvA+vkK4dM3tJAF/VsNhRGtaSNLWV0N37qwx8UnmL2f97cPVsQ7yURKx5L
W4IrmrZuPI0P2CyhqpDtpiF33L2wEP0hFjcP+fwRAoIzKJD1KkzieGjR1FeNQtCFGTT0eS6NVXIP
aW36PTkY+9LThqaOUpCzEKMjkgoGVBFmby5CmGJ6apjitEYJIr1owY5k/euu89f+YQfjp2wPYX1C
UTqkny/Z2Rm+UxKc3rvjVvvGQdOESMe4x1PdtJyr4AjYXwOrS43NK/QnnaHc2jfvF8oyjXdSAmZh
XUDYMOrAY1OnyvbEMsQ7d86lbE1i2KMvBFbzK0/cIR18v66EVM8dCvXxgDk0NQuoAmp8LPDXm+Rh
dWVCB6idYRjSL6ZHaCSZIK8tgK6QaGT7UucEg/gMiqjiGJmISJ3+37ymvV5mO4i6MDwc//jG/Oe/
6Zd9dKf+QvVP/GCsL98xqkhw4yR6Lg4K6Kd2skztmMHgUDXOhHSmHGgpRX52DqiC98+eExl7cnC2
aE55EKKniIw/w0hXCNGz1lnweNJWNtE4JRiHkYlF62/6ptj5RU8FbxsiKQatohQtaqv1ImQ2XXHo
8RgyQIzUXhs1D7nGx6nqyAApagxGREDGkMGU6OSWk43IILoWnSGOyRvD/A8cjaTJytioBqAwvKJr
dKiIxr47SnDEn98ZIDfavYA9zLITLLlhwWDohAmPZCRtV4gCP66cmiGLwjzfsy/vdzHCpz6tzNCd
Hl9cq8e70h+9BV0jUhqOTjqeByekDOabkGDzIBexuGtPXXqdVlFeskbzQ38l/U0hFejzcEwZlxRm
meoUiTvWLqUGTBKZJs/BbO6lzHTbdrP+dvqI3okY+h+MhZT+gL98uhsX81s0W/11fETGVxo3KzQt
3OVIwVZkRyiQInqOicBgpqTd+AbwAvHqDZqYPBud7e19DLUBZa2AJju33kdfsHKnpR8lANvNMgyF
jV2/uyxJkEPsXBgnlp3MPoAyxOwdMFRhIjEGQs5cyYVY6oQAp2Za4y/AT3d9cRR/ef+3500FJgXG
SLCt14fdm/x4TxSzD3gz02UEQ83oCYEN7JuSraUOGVbh9yUqdGLSJ7KVNZj8tBzQlXWCwBXZ/TKf
MR4AHVksuyRp5S0V1foELyVGZoIByzuAi4FlUXOuXRTAeKaBzXKJdovaKWSe5iPX/5ZH90vCs36h
sP/1a4Nd3llqrgNB+AxWpVtcOtIj+P8W9IO3CXo3SOPnA2Zg/CnpVDCCOftYSgGW5htfBxA26dYd
4gpSc7cAtXBVvL0d68PKOSAbspOlR8r4ojBe57+oJ6Hyq+kFsSfM8x26c+c4hqnfcfAokARvMdxb
dLDHH+dYHj1g4nmido8CkUtl25B/GN5M5dYxZr6cdhvTJR01ZJVmvc0GlcmQBp3uD+ecVcc4s+sV
A8eOJu0LufMG1UcXv+ixlrO8kVG4XfINEoPJa/bMvMJ8OpU0rSd4a3rSEb/ncc3ZEJFSKdXtmalh
2raHRxyDxqxU7eZZ9Uhmb3IAhawq/DE1Bz5YhBnvRhaXIT5uYw93sTmKJk78PtcYGTpwsP5YHBNC
c9ADtkNcZWbAIMr24/S0zHcb4ktyJXbwWy+gd/qRuCyo+88Nw1Any8o5qaAE6bScnd+QjDySx1zS
GxTfvsiivSoPXenXJBoq5ZyEasj87lh7uMWy95Z8Vj3cyAYXGx9j7t3+XoSoThurq2sXEXhagp0a
NTHlMa3DG2GHTkedIC5ni4pBtcQ23bLKWVHTYcgi6L+BgS+K2YPXQjI26nRYL+YpJnornjxGeRL7
5YfKE1jwABXgUmZqtkz5fTXWfr0aiSxruE3cHYwOBYkriQq91IJr3ssLnbsriivpeDUCVl0OtSfZ
bMlbCBqabyeDiNAnJ/LLfzFVAlPq3fhIcI9/AlDFCnzp9jnc27lsJt6L6P+1KAVfva+v+M/0QnO1
GmqSd+X8t5ukjqz2iFRS1kT/cz3aVUoVzgT6CuHn0nWCI/CQ6bRD2hEdhkXynNFsPHNaXdjtHAFX
DfiwEwHizV2g7eIxjAVsCU7q7jiP/KSdLDGcdfeErfE7ctStNCbUHBHfPSJABC57NRk+4m5LcVkA
AwsE9EtVDD3oxfzAQ7cVWHamO68k2QGPDugOJQxN1xUbdplY4lrvKe/01TDtC+X8+SRXFXwlaeuf
gSFvI9/wvonSyIf0k9PrJAdPyQvCYX0cwMYXxTI39vSQ4zYLf1JCQIhmp1wY2UPIsmj7IvR2IFkU
/CdefToAztWMIdy5XDt6fj9OYEomZLUL4nfMlUFIbqSwRYqWBula1vLrB3MEFemVybeNTQx6x46f
NCQBeStSdomSCiPYE+QJXaHtgP9kn/vovYDNnFBtsx5mVlnhgLpsaazIvQGXcm2v00VEmW/FAgjx
j2deDuzorR2VywN0aiDDqp9AaPN8BtUbb9sCvhlmfikyBCd76tI5GK+BMQAWtkZBjo6zytP+6JZu
EQArUAoaBsWOOYQCEMJ52RVk+X7e5yoJ1A6y/m4b9llq1Jz5K08IIFXcoOZCF5VetZ+2PQAmMV3v
t9SdF3Lc+3SN+pqrcEMDOTuiltpsCv1BqVy2CsPBGgY9D832cUxsfN6BCX3g3NZJ9q90ZLPe1FAa
cQQ+d7mB12tUag+WsYH1vuEoycxv2FOE/qSTxiEsm22HMgSmKLYUHq7KnvnrESTlK6EcGJNPsxgP
mj6ZDhs3lOphxN+QQXwSQzRLl6CVya7shDE7lDFjMwlE3zAX7OJLQMMn8edNTsct+EiFHAfPopnX
FuHlSBfXoEhBcPBlRH5/rBjm41HZuGpJlgDnI+U2mg0PWF4nIqI6CLmrYonf95caab62VJ+pOmeU
DTJ/zoJ6+fW31np/4bO2dKQTIhmP51pzkCm4s2nZSJdpEn38jUXUEZ3loVztU4e/Sre5Nwa3P81T
UyzIsp3yGLJgzGgf2MXZwVDbr15GsAEAWg2xSHRj4oqE8O4A0MHDonqJa2YXJhQLAQ4gcoaXRlRu
upnL+B9TOH0tfbZttqNWXy+Hp75OeNHGJThXJwqT4Y82qR9SrX6NnExBaoQ9oAcsKhZN4l6Kao+Q
y9IjLGlvwos/mosDIfjQK74MzgZ9uPYg9fRqzWYk6Wtxf2tsdOyPAWh3kxY64bxIq8qoGiyenVWF
DqoS20mDrtzC8IIsvbk9Vk+jchP2DGmrR/UBfX70dM2BOncFNLOeCHXRblDSN1G1QIVEksVC5TpG
/b5DSECZ9DRgp4QC3g67JFQOq2G790R/wWfWclSf7tCKfDwDpn7fWywOEZEXDSi5V5Xz9kB27PV1
PFGHNB5agjRc2JtJTa62L84Xm3c8hNqQQ4vcTYbpb5x6olTxU6WzPNUsgDKXjsJkYvWkz+89IBuR
teGR3gmunO7BrqOheldBpHnnTqEMxhkDo4rxg7QEZu24THlEZc8wB1b25Eo2D3rnl6mxbVmenWQr
V7xuQqUhnjivacxFmKwmVBTcH22SMP5O25PNiCyq8dk/2XK+okxrFgy+gOm+kN3hRMq4lhjcHdNd
mH97EBL8ENGeNwzrkDpj61y2AyRUobBdeV3liNXTet5o0KaKZAzvmvt5UPOwH0KzmHKjqWogTspv
wxHXkz59ptZDup7tX9t8bURXb9WDZ7thyPEjVn9BDpajDpC2N3nBC/VrqzEK8kBFwQQuIzXRsIyc
JbcGQScX2fYVwQa1+inYHYYHnNxn7vw0af0MdBN4dd5Cf2QUjMhewNb+jF8gaJ6dsPpfTKZK9UIJ
Y3/qPn/CQezVFCNsNGlKD1sJvJUVUfV+QB+GE/2TyFzn4YND5mFOn+RXcYN/s3Wfkf+J8EfAun4W
1JZd/exohMNomGqzO+ScBoeHoK82FbqH58K6LKoKXM9sBqoeuUpa0VOG1FUsWg1DqpMUsNWYi2jz
TOQpdnwhawskfF27QSKt4Te/nwcNjyB9g69YdmUV+AnuOcSUIpUC9ZK/mQN2KrjcagTBgVR+wnBb
NOr91hHwBU9DjNdC5qJ0VMWh6CDGuIiNlCLjTefPT4RH/3Pmj4A9O1by1tuKN+ohprRgjMEFK5a4
ae1daE1RDyPdhXxdR2VhQrTA4a7KlmYVVM6xZrFRr6CtvIJ/TAoKPetFRxfVnVcPNeEY6k3+eUmF
F9cWHVYOqsDJ52Qjmgok6dRft859A41OGEfhbEdq6xHIQXnxbOECpH9KAH6N/x2qW2Gm05Jk+K4h
2xiLQpasF/4lwmCfmkYHDlCExiZkebHR/U9zCIYcvEIHDwULt6BNrnqDUo98ZXHkvL5ideQniYrk
P1oUUJAjSUUu/XNH3fDg2Aa6MQ2+IHc7aVUBNNUDeELT8lDSkTCjBmtA87yOIn9TBu2ZTHt0aW3n
o3BqSmT4MRrIojh8Mu1OHJgcAjEyWOr4uqbqQKCpetVcMDa1YF3b8Y8M1g5iLPMPpLFh8CAoqYjG
w+1zV8KgR+iRYPXXtIRDcGraAGJlkWNxk1zASQjZDr5Y2JrbezEoaymMA1TF9E7kdyoyj4UwfW2e
pvfFshG1YFiNeTfUumw0N7bMmlw0oFkG/9PBEqE4nN2E0FSDdTDlbXCjMlKU+NCveEQ27O0S7ZtU
saaXn6Lk/5eSAYnLbwoDgxRA5418Ec5yBUvrckAsKvgwKX71Nn09ICZjrQRRvzAs/MliRV9a6iud
YWRytR76DXuPljp7mRfhV7qVbbCl8kCxd8vkFiBj/iAN1YeySxOdr5ZZKsSy+tBVbSQE3o9+g1Dn
GN2feW85OvBvncRfMeWSMcZicr21I/l+ah5ORzIp0M73RIQAjiag/ieO6441vc3paTeyv7qfuQRl
cZgkmzR1dp8JxXnx7myvINXZvmX1OQfw3IpbAMPlM+OUBaIHMR8/Wo5tZ8Yd0c37Y6rz0y3fVh7y
2mtuYorFP3QOXrMjfd/CMeALnk/YiPtk3Ls+xZSYLgqCB/XyDObi1YaT1IXHcAGU8c8QOegeFlG6
nhMy9KngrDk/1Hv1/ZeOhvZtvuYuSEJWDX0bsQ2VjgA4khlfsnOzKwfEBZ2+cq8uc31usl+y0XmM
f/BKMkHKIYqaCjRENtasmsUJ8z8G1+6616jdLT/EgcMe/rNaTSDfuOBEEjGOPkCIN+hvkY7vsB8K
+OgaCbZjfHMUYcy0lsz+jWoY9at2p3CTXq6elV7QcOCYSzX/SuykTVOYfHpxmmb3tdsw2XgGaLBN
tpe/+EHzv60d8KIDA816kelaoYDgEXYI9E8utUckAGV5nbxGFHaLkYXm5Dk8aI+mgqKtwyFMrqFi
5FUJIPAlZf7Qpp6epLGhzbTvITrfcH8mzXMeNpj8pAzjNIPzZU6/S9uwwlbd59JQxQy+j90OEX7y
PO5A1Y8hyISKqvZs38/aTGoiFgedmYL8WZ6JHT9JvK32iL0lH6suwaMnTLG27QviH67owuHxy0GY
1ZAwJA8Lz1Bb0kMv5JamIgblBPxblSYFymBvZNKeWvUPmFNunlt+6SlfXv5ObNbOMUnol5QKPGR7
9hFl6aE8S9QTQhnRilHUyNnahcrYQR9pdqHgq5ipyegn6qDmKJHktgq3b/MaKleKfubGunYj69au
eV34rqE0JlF9cMlztcE+M2kvRzK5RxEVwuCZKb8I42wCM7dy5oQzWZwp5qZcu1rA8eHLMOAlFQ8j
/LFPyq0TF8p5NNLzDswTpwonfoAXbd1Bb37ki5RVneIo7rmAKYsIsGOPlPyRTqCXJZZwNS/qxeuj
SfqabHg7zTr8P62eJQUJEp7UIrAWNkHIXUc0knPQf7NRYBuWBmwgjLaqq7UF6Hc/t8qmHxGbTto2
HZXdLfsNYd4PGspQYyhawrjNGSliqQrJUDoXUiRX6jM9xTeH/1A4AUkvdKvcn6kGmnYYFlANOf0d
pM5lBdgM02cjk7m7ztWDkIH4B8UZBalLyrJ0JRS+LTimKNBovhYrKyafITyoOkFPOxJqlRgDxhIH
CeEKRTzVR0Mpcdlok9MbXStNdeJKIH3MGhOAzx2coA4NkwTKlX2OVu5vo2XZtBJoGiyq6v8oP2fm
czFzNjZthO40kGHNcB10gCCZ6j8hs+gMBKYoYBDPLmiCD72xLoPLcB5d0mz/lWP1vQO5lSquH1cg
Q+6ckwacUgFkkhQpWImEsG34C8mrtR+yCLExHdkbysfeZNF+zi8R1hn2Rr4pAvqCnRrfHNksxImF
W7doJoRcucgta1P3ck23523QkYDeB0JKUX9DyalRQ02TOkSJumc0skjLYkDFEZ7buk5geL2OKgXl
kaOqUoFHSEm6gM9P+hI0RVt8uY4jzt+6yxpcdsp0kXLIx0J4W1scfp/NgWY4Q5EGBpkohPtUZJVC
n4CiKREpOzL/oPbVGb4OwYn+eHbSXHAsqRLcB/FcvIh2a6v8RJwbXeBwuoskvHxVxNDDe+mR5ayo
lJhjbWKQcUTg+6TR58EcADOU5+O0zXnRYwOHN/ZP1XKOrxZoDVpYt9iGJfZnG4jLbnN7wGxmX5xB
CvBfESfSmRdG0Nu912U7LK372f/NmeiuUukh4G8KzS1+HO38h6NzGUTyira9kW+AlECC2iZ9PosD
Uyfse5HmuhIAtOw43e9Jgrpiaaz0ufHJ6YNZWvO4pDEEowgz2eZxYlHLA99kVA/oUDz50NiBdDeQ
EU+QVfzoAKIuBXXoY7DUt5vXwFb/mdKfpbQe4nWNocER4p5g39W/VP0yK+Ddm8rViO5hVHRdpCe+
ENiAM3CShF1S2w8JIv8ELjid23KN4ashM8nwIr/GhHVVeI9PjWilruqdBsHqlE3104B7AVRJ9yKi
ppkb6G8KWNPgL1+jLYemRE9L04+MJvmorQAZIrj96uR6HMMgxDqAFn+VIq2pJ8kuVeNkBdoAUO+p
5ZY28kBVgDY6nW6TFA4639qhoNaDYhcmsR8N5BFRgTZKtj+dpHtBiBuSW6l3ptnJcUKiHNuCLagl
3kz5TCn8xBQdPIqPyzDvLSvr6Wo+r68z6lB6u41d05A0CxdJ7ZpSAk4AlssExP4zUTQlGJ7QBy3X
dn1r8aGfWXt6Mv9EFNZMSh1WrlGGGxWv5NwlYfD5GIczRLaRogJpZr5FJ4KDUBIRgWWh86haa0sw
iJBwSe6nEaYy1xev4/AW9pKXu7TaXk3ukRZVD/CnVX3W8zSeEi1GTFS5hZPFK0p5yqGFNTMEKCNq
WvMYhmGzt2qMgNAZdnDVNWxnYIvTP1f1REt1lLwaBGa2RvqtHb5NJESrL0n3FtUKcFy9gBfNy3lf
p+1miNZ2rYsZQQqyMz6Eshv8olu3tCetyUoqUBGLA1uOxBGhPmgIszOEjMyJq/t26/geWgo+xOfy
yFMSQdu7WTl/U4L3dxKnkrQTFPDkuE6+0FhrzSjPtE+MXkYGqeVSoOnqQiawsP4OiHZQaVOeRrkw
1LfQzcydamKGQMUNJVZpQFRqoJMCP0J7x7TVO5P4+MvGm2+4Ebqr2T1HpSVrkYZ2S6ZctkJjmN3k
t2fQSeZTKnWoy8Lk9l+JOVKITojpFIVBuIrg2HGCKTy+UiA3/qGP379tXGwIaLQAljA7cIIRC0rf
Gid7Ip6P8jSArWUAOk+3WEasqV9Qhsb5WqeTaI24Uw2sW9O8Pdu4RQsILlM50/odQdLaxWQY7gC+
UbmgUVwZxxDA+eth8UZ0W5GowHWMf0h3GeEI4gmI0tjIPCFqezLvH3zXsfLxc2t6/ja/8ou5U28a
j5vgh9Jw6JIDyBDiBQJpM0dP9Xws25YE7jUWA8B1irq7YyNd2JpRtBiwkU6Jds3/dG+QP7EtDkTy
B8u0iZTMcrEIZnxufXC10UEr+KlB/cA7yhknngUYcTsLdVOWarA1PnjAbCd61n0CDUx69JjrCqM6
xfbNNw3vbO3RkEAvOevMRIBoAfnTML8SFXEb8BQl7Z8TkoUvvmLDpXln6EDBcQCr90eVKc5JatXw
Bhjb/p7z35FSWdFgREOdfsJWQvXuBFa71iTzLO9aCn1OCv9PPKY9AGCut6klkEv2L9dL02GcQqws
shhbMlxvSf5elJ+apJBAfgGuSIZOkXaMJAUe2s1atxyzQ/YD9u3pJ/ZZoNq4/Rq8Lp9D5rJGE3/+
fRvQ+teJVzY3JHRVinWYo0581efugENB5AhOqYOxQHsCpDvUpUDudmoC/AIYzqvEk+hwmSLlml8o
Bbwi2n8cYLYRyB6hukx/gM5h+3jdxIfrbbUSOg0QhQ1K9cQ7UfXTPsN7f334q5/a8tb+spZn5bU1
2VuAin3+WdBBecoG1Ioc/qKbtMeK1Nkikgxfya8UCwt/009Vzc1WeBZvGFwGP8Rdf5a8n5i7JTyY
SrxnkGPw2+EPg8WI92HGL40CrRaXRqrXfWIfzbe4VKhybccWWylw+/nd3MXtpyCNY0LdEP+1G5lo
9YTsp8264t4Wxt3ThA1R1OsSKcDPipEJMq4cFqEVJI1CxV6NpfUsr7RmUne9ZUr/DLKWnDsOznsl
Ml0mzmd75vSsf8+d9hNhSnf1nQZENWZWEHLXZYs0YrRnlRw5A/Sh5RJ/Lq0DxFN5gWtB1EpuhLtH
n2YmjWTunVHVTiVWkvA4Tl+wh4c1pQoBTqDu8l924TwfTWWgbD6NpZsr/H7YNOHDiVpSY7LTZSaB
WXuLEs0DV6xx3IOYdr8Eoz8p/pOwYbDJ90p7c/aZYm+dP3zWJGWMg8OyqHqqOU9f+OeAU1FviTzO
/JUiTg8zPo9/Vo6F05R/pcSMO4mfu/oNW5c/+bdJvb7cFwDO8/KpxDpalTsiC0CEbPmcYt3UYcMQ
xP9R9AW8cjKcf+XfIQQPXxXTsJ5jqEo8TbMxsTshDIY8IPCQItYVqr44DZoZ1sEvbirXfRvLumCy
nCwWd+JE9D4b7zXQRl1K2/OS2GaR8ENLO0mlvOo+EmmNBDS/gF3plqQn69xtkbM5XcWYSvpO1m2W
cbGzuBPX887LzTXnMuwWiXYDGgYIu41xqdSw3iTlsULNCuOuvg/RKv5Fsz1CfSkiAUozLHZHz3lV
r1TzAed/9tMk60bXx4in01hn102trWploHiEOpoLdWggXxOzorGX2u+ZGA4zU99ohMqpCuvoMFaN
lPuI4Tws3S58fAcUsalyf8b74hqVzYFNd9lzHjN+DIkZ62WGw/ujJDxxdav84S5UH0NuI9WPt0/w
2uKuGaBom0w2/DGzZwWkhWu3gMuUaJYW/NcpLGP4CdxSyCR5RJ45nPOxxB9HD5OH9Xj2GSNc+vgU
uzIiNxAvX1gg8bn6+sROayeHqdV+j4BJUmM7V4o9wYKDa+6BavYl40zbiKtL6DhpfWw+BzoCA3Dv
ZAv5jA+2Dka4n2BAlAgdj5QQPbK4l/3rg86xaMXCQ2m4dgsILpaqhD6/GoY85wjEHz+DB1ZRcLwZ
PfHka9jXhh2lyV5ihW5T7NPUAs1xiJRDREM3YkjZpdKEq2jJtbfKnD0posJVTtVIPZIS3aMC8jCu
OAbWZQoND3aXat8+oMMvppYqvUj+tKdCfCj30r9qc789JPRROT8D1/+DNggaIkfLahpiBoSxk2Dd
fhth1THpOXgmFCU54HJpLmw9y8KX5a0ibDqCN5j5RmOk7s4XLsAKMgpqaDZj20nkuEtVrk53bXBf
TNmjGJSZtjtaGcMGej8Hz5LTz4vTU8vVLpwFc1MfUvbT4f/cp9aeoFzqcUCX1T64XJ0gvQz/YJ3j
6ntpAYGaLm65HdoyrwSsG+2zHYTJlWwTUX539DsxM7U12Fwq1jsRgvno3CcekFrdxSHZ/2il6W3W
7PL0N6ilrSo5PfGAzBc/u0b6wwVdVifzNUrpAVU9K+uVR1OPkpX6nTxaima5QC2RmigHrHCA9jmv
/hskBy+5SvPu6XJWu21V8WuK3prqOUi+ECpLrYj6Xlbfx5GogpAqqJDsOp9SAw3S/aOJ8a9QQiH8
Pmw2SGnAGTgh423at+zPLiLxTJ9r0wczEuorSOAQXMC/HN5JC8mhzPm2Q3Xnq+UEG4+Fit0AxZdF
qReLXZYY6Jb4/l5vkWZ2kbJA4EKTR4kd3JTYMNnoNkLVHgIJwWr7YWoJGvRuGTC8UYO3KiHja1gB
BmMhPpNt7ULKEqowfz4YpEp1FGaK7ngD9tXSqcnoVFLf39kcgG7Zub4sulqhRAQyybPNk3YFJQtV
uV6un2/k1wWXgsZjTtAWxu/oYFXGU0dl1nMnOKVG4p/zitquL3y0s1ojV/FfG4x9JFbNRldvCzIc
z6gW+FtChKmWrflnG5bDvBljLy/K8IGm56LQCm5WRaHboOwrqiB0HRqSVwOXXXMMth3yyJnl04jx
8EMy9Lw+dpXO/0c8E1qVVB7VBwqyRObXlqEKwkJfgHafmJHhkJ5rNEuLhKCPSbFgGNHhallPrbMC
y+u3WMrcdrmYsDigjOIl02HYhwzPfuMq/0Rd7fGHBWVYCuWaTkEpOAZgmVdJzdPZjGdm8afoxXbN
0ITpp6p3PwPpAuQkpbRTqxsEG92e3YZFvZ+WGZlp3KG81ie4IBO/EX7DEQ9nHBVZs2SOjj0W4IAA
U2vLssYPguPucnMGJct7BFEU7rTK2l8QvfLnNU3CqK8931LTtsMaFoyC3yx/XJtAQteeU2g0CUNM
G8xkzbVWoJfLdg7Y3Jki80em8IKORsqOXIY4fCwnNPOU99aLBexfRZdg+EkcP4zxJ6nELxx8duux
puxtOsS2EY2RKPVlqZde316CCESrNb80V+rFWyhrgNnkMOu4480RZBQy4Yskh62Xw/nGbx8foK1G
nca9xlWesKeUVqPrRczMnpzC5XjdUwAMvBnpS/9Y9ERzYwprF76DILZoE0GtBFui/Rh/km1oFFrw
pbTcoTfsEBtcDyPTdk6qZUWtCxESuHz/Hpqi9hfypshL6tmoZYgIRWnSgV3edr6C0q701EaQAzP+
V9vvsxMbYPT3WYfyMUsv1WYhjmozUIfyL4ttKolatBBn9AVwHcqgNaQP57PcBOBo7hoCE5EYwe52
aV0T6rK1+VZuinM1SFITcqZ2HZB40LxCxs8p8B0ngiZ95SOvlj/0/MejFXQriBOFng2aCR8mtaHN
F36K7aeM3IwQVWatbuk7+q3uy4q7TDom8WIJpXH+Ggbhi6x2CRTt6ZapagiAjT0UwXbSsPhlMJTc
EETjaCFcIgjCCJm71okuVYuGNJQ8UpI+9XEVCPCfVG6d4R80av4ScGPWV/ImZ4IuTZrqSvzCpkAH
6971ZPnnpXLJAPB9+7Zk/Ladiuz8iz8N1xWPRwqJ3FcnnpYCjWm/Mi2cTDyeJpW3QXAsOTQSJXVs
sLmWl6OlFqlPclicT1kL3k/bBNQEGPRHt8VjLCnVGXENS3C3J/Yy4iSRZnCZgDRz1GiNmACB4rQV
zhy87ovn1LUbF9UnoU7IN/ttRv5A8ayO/+wC+c4kSX2VP0x0b3wRnnhqYukhyJEPqzM9qOoN2ete
P1/hoC4niH4Ufpy89DKSJ1X5DkcF79gCkQ9mTQBhOXFceU68e8VuvP0Zsz8uJgZYmD70UAQoTnGb
M8zoefR8x0v0glfW8YR/RPXJC/5eVPBURAsjdom8BzYXf2jz9c8HsNyaWL1ryQt5Nn9X65UTJ77i
x+57zDtwKgER8hYYzzkba6dc+Retyr4I4q3TBjQOfMQ5VEPaR06+7ixeF73l5EltftD9XOaHSjil
Zt9CUUbd9hXKECI1aWPfDEJ3mBqJeLSMJQRdnLLGLT2ZoflqhTsPXJJt7O2d4W5fpLr9ay6iwN2E
xl6x46KY8vHbsnBqvY7DoK2m6QNwD5m5LWAf/QlWTbZuBfs6Ac4Rhw6Zwsqp6jWm60jNFtGCHO2b
C7/qANGVblp3IZu86u5RrGdbDpQ1iuMJDpZ0MfZQonKVnUNZwTIVHGre2RXk4SHaLuAMJufNGH0W
lTXa/RABz5JfhVs/MUpMyHTu2ZBj9YXj15KfV3ibP+hH6KfGaDqwufYpeexDKno1OES5Tda1xHPJ
kWqv7b3WXq833XX6cZjH1dFzrWdQA9F5L3ikoiQfBcR/MYybeQG5WRiweqtDO22Pnhn/Nmm76pl1
8/N7TdvZ/dqwPBlrmapC67lG+s3OX52K4FI1yg5Lxx3wzC1pQJhwY2VGyzuZGUyduayDErlz9N1V
lej5BAhQezhWmVaHHKalWSmJQQx71rmY5rAz/lzu4yKD6+sxjw9vs1FBeXM4Rqopip9+mLYZrFfI
N9t139FvoiMrAoL5f97xWLcUC0yXE4LPpYjPdyxNgjTyEGYEUsgNt1gMgmfZpbZi1gycDY3d7F+b
byVDEthuy4GoJUtvk9sY2vCTNSaQ3P+N79n5ZI9TtYqpyWHdf/4RfYrouZD7UnpFFSeu6cou2huN
yAIqI2ekIB9/5meM16OaFd60OissAOp0FcHgsNeEeK475WPrt3gvZwOSDeVqd3RF4dEf41u8vYqi
0hCwF2jr4hiZNDG1VGwGeMJmgbWyX5k/Qi5CyuLWUU94FCkhkYXeaA3+ZVrR3JYUr6uk3ax/1QT2
uBbDPQfhWTgcSLsRwml1JGKStbJkjzl3dCrCEm2nobhJvvHkct86zYbwDA//k6c/2NCuwnKLHyGZ
TpiDQlomhqoPlRmSrUVV0Rf2wePKZCguEaUMUQWJvlx8AEZeT9rRh1haQl4FHtEj0HDeQRXHB8hP
plJYL+udGqijzFbnkg+h6hqjQe0TRpsw8B4qvlwCChD005AhEQ7u9wzZEtAn4Nbm5qTqOlIE26Vk
XvtpurUT+GJT2Z2ATWb38HxzFko+AvFXEneevS9AIE8aMtd//5AHqqm7BBOs0quXCVHpf1UTS4iU
LoX3oLjaE/k4eGVBrf5aeFOxKIJyX33ge7mvJLFXHIuQbqtv2xFZLOQlLWmsd4wvARvPBftktUff
WDzXlAN6WFebWbe7ca2kjwh3IXDgefAsxUvJbWVBjyfG0ILDHPYee2PIrpXbzfAwxPtzUHk1Od+d
x4d3LTxkwf0TWT2WErAqI2znc851LPLiZliMhtsAWhdZFEuDNwqOzmQ1MXLDm2telqS2sKVftD+y
hSGlHx1rICNBeHibl/x6EkAlllM4WXIzHx2ldQLEw9TcFJMs94TLH6shyUvh8bXMIWrCftimt1cx
P392BYVaL7pN50iTJsSqXC6fEFN3fx3xecxGKRwi+PzqkFdspSuoLiHr58c9Lc0YoTu8mAhPrTLl
BGgTIrXzR4Kr4Kuh5hxh6y7HA9TT4+eSFJ1tm7vlm5/MgxVEFQBwG9jPrDLVsrSSifFTYitzVj4I
doLekHX6Xi3xTf4yfBQCBPmtNIW7YMoqmZx8RkAub8Xr6n+kgQ6dAuuyXjdQIN2H9Db2fsXwFz/q
8MXt6VTGpKECZoi7ingMAG8UflqBXGWM3i/1dyz6oK5sCVEey4aZgRCS1j0NOhlyH8mN4gJIGDcj
vdo6vX+Zk4Dr5ap1xjrnPEfWHVMJ4BGCT463WnRqJ1OdPwd4rtcMuHKY+6myd8JkZrLtTBxadssy
xqaGSZhGCvlItVDyTt350fzTeFhb3tt22RxVgw8cqIRsIieclhCCFzKr9h9HvN4mCLKbKOfq5Bbq
YI4LZ3hg1480FZ5GOmB3s27POeHb4ftFzzuyLNSalkqukWeLsXE7M3Cxe8UQifABdkKRVcKclegH
Okb2ohlX5JdScj3k2D9fXzEsqxlXcO4e50b2S2SYi/sJ+eVoaJQCCE5nBoo96yamvlbrkF0Rfm38
ny+nb4Mhz/UYkVLM+b0WCBeL9vBTbAiuKX8JnW8qTe2IyKRqmglLK+wTWU4UTRIZv1FX2n48VfHO
YYODBBMWneQHeUJiOzs0A5Of+5K3atpL3Zb7nyIQ6Heynh0y5039ofGbhCT48hlSmonxD8B8zcx7
iJkosi87see24I9ckBiusY6B/CPNLAwTI09rLAWVbsLCWdTbg1ZQ8mpHJb9Q5uTDMj7THe8D5ElO
6wkKDqSiQU/9as9Mm5HjKFyJcYRdRIGv+OS9QIQfcFAi9TGEpRvpUlpAykx9OEOg3B4MA14ykKu2
mhevaFJWHub2F6Meg8K9ru9kMM3bc6VdlfqlZI6TwLjML/jCsqeDQ0E76blXus/MuTBNWBtyNKVR
Bd6YiY8fhnsZrRioBYd6kAPWEPKigbJ0+phpVqZuPBS//WdpcjQbNWnDzrljcUnqeTtS7a88jxMs
xaXoWV1rgrXrwDUOBI4A1TwOhObYiVjSaTbvrrgaJl9OrCVzZYWg8Ux4ZygT7WHvomgKklgpFh+O
4uw+x3kj0GhIK6CjChir9PkzVfPx/Sw15T7YpyjbfDV1gRbQDWNihvV9TwoYhIIa/z/JVq9iBBl4
VSjkRq1sg+2wUDj9tuKo0q3CZoWC2wKEiBgbJhh9OhOkeGgRO9SdoLdofMpdpAtuouhfkvjI0LWq
Oqa+iLiVgxVp5fVgzna2IMbVgtUMoYUYSOo+zut8MBd9CFWTA9Wjkxt02fADH3rrqmze8OxSq0Yz
Ndh0fEWzRuWV+5zYb0Qx4sdlNZqZ6hLVcSZ+bAOqpsRPs5ndqvXyrCZPSp4hthXnxCD45Z9f0o7E
m7Lh0w4Tm3gkQcenDHJTDN3GjubnNqJg2H5Rym38I12oCEvXadO/L89qaTY4ZxIXy3LI3lRVqnkv
ks4LY6dPw/086hw2bRroHTi1zz5K8T0O0yyKvhPqUlttVrASVwAwQCGfwW6kC8Vq06wVpmXGW5pB
WSn/wZdJ6rTHOluRZBer4KKP6e+ltZk6/6hRu0y7ZcvksP81Br944g5UbxAs4UG0Hh40zeR5PBkN
bwot9nxDj5jhWrHi85noi+oDRcREuYO4zCBkKAolt6qCyjpzWoyLeNkjBsJqhHDj/V/MtMrCB1SG
3f6eBATjfMv7gDRAx/uzW2DPN8C8BGrBuwh7WeokIzPVJYV7ofbyfUMIe+HXzOuBWGZwZ1VyUy4F
diazUVg75/MJKWOKe+/O9iMVsxoxe1yn/YX6Mgne0MwUGhhTcZjYb2rk3hn4u0MBjoDSoPWqHdD4
89vafw6M28ajX6CYVgE4N6C+aByUkvXVfHH+dmIQ1TcvGJ8w/OiRDgq1v67WsGbc4Xq/q6ILJpCa
6Rj5uxeDNRwgeJKq0TKTjIXKEZ4LJcV7Vzll6wpt1WwF4gcGwL1DIGgcax/8ISqQ3KQQdHB76QoD
9SWSOviIEARs12P8uK90x3iKqYq8/qN2OWtkAjEge7JbE+EgrX+uQKyaGLOz0oECEX33B6iU7HGt
F163PhcuHA5Q7YZxCXNdKpT2gDsgh/dHx+hQeULeyrPSlewKFjGnA2zXKdSvCMXh6VGjD0y3s+Gi
IVRA9AR5yQp9zKupdXeAc44UvU/EhFoVq4aUshhuAPOwXNUGzQN67UDmf1Pz2+3Y5ivK35J6dVtC
fpEgcQbZODzJnTAQjb/purOGDXIgLqy5pIK+Rmy1gMSm298PGrbTesluo4X0thvt0UeCmMB7uaue
QX+cUVjXBexu4mzYxkOFGcAC9EhakDCZZcJA1haiz29s+oqLhI13IE74Rk3FqEXuECJW1109l5TD
a6GUEKRpl27gZzuY9dw4tz3DN/VYIIuwE/6NOKzQB9nib/sR4Coi0undcrbdYOuiCJrAf3heMmaB
LxL7eh8SdBjaLrvkFGHKrN6vuWLGJBLe4TIyFeAkRE1GtO9XxLAkq/fqOmzwlkewRnqgzZeStmR4
A9Ke27CdYfKquhcW2fcjpMHxQelGynIEXxhij1ugdsxpjlMEbN4j7eWCIzVfjULUXkJoolyUqjkH
cP4UnBHD7qYDsykuV0VYozOxjXoYfITgJ7ZLbBUqnfMliHL4CqupwxmjJcPXzjn3n0Bxl3p7k996
Y+v96arvSC3blfXnOwaND4xqZgLMMwP1VSp8PJzZbnmdgAydatyiEpc1oK8I7+2cNdkbfh+P+C+k
dPexRmtpLNGpCSGZT/Pk18T+/tAir1MThcNhnU+LVatPpviy3bcyLcftN53764MKKwRXAQeLKWvk
CPPmfrH85OzoBseQk/h+Ct9wimlQ9BGnMkF1WyikgivswAZ5WYLo3+0Lh/tAQfVk8732xVUBLNhZ
ScpHLiDjZWeC+eIW6Il11oJdz4KZw8ZYfRvTEHIFdSVsvvjIOiWwuVRK4joTeZFibmIjDUl4hARg
qj4RT50boxFBRkpvIKc4WrxGF63eWKQfAiE0TXZLIGHR8KAU735MlTzZCl746ObES0GC4TxPpPCd
KtPa0u1F+QicsvN2AbVZ0uGT9RgtkaMFIM7DfTMKVdg3d2xS8XzorfpNnewdsdmeEcvxCsNyDG6B
0Ro8BLdwWU/TOe1JS8i7LzXeX8o7zdW7i056kUmp7XsyWypt1q6WHK+bL9Pt7yiEvQaJLCd8eJIC
lTqebJgaMVGClQOJd3EgDj7x0IieC0QnFQAQukhrlpupTm6NWTf12NLiwtvEnzass3r0nauL4d0j
AhOiK8LzDo/BiJRVRgKNO+RDTLY+MvvKC601VIP+Mi4gMYScTyJjdTe/sxDX/DlTUGGpnr3KewYN
X3rvjla1u9e7LfAZOEIhn0tilhca8y8UiG4/9i5PlXBpgayv3rsdfbDaWDbP7eK/wWBcdjMQPNT5
2tjatrI/Sx+baMokmRotYCElipsJYbP4293H4dFlIIL9a2GVoZCTOc/LkBcpX3QqymLnibaGiyiU
f2WlyQW/nBaEAOLSF14PXTs9nOIAIilqaXEz+24bgIinKul2K1NZVv+Z/5ohyc6PxS4EkUchtaEP
wDVNTa1k5Use80vjRtJMsXFVmyhXkLx8SIUr758TjTBk3was9iw/mRo5cZf2Nui1B/zlCQu7oikC
cpP2LH+/McA/4dwVdbt8DJ60ctcC59i+xdxZwv+5gcdJYqqZHcSoPNa5fx/yj0WaDAbmTXG4ozM0
HLRRZHTv00HyomuCYsDR8SEdUnI5m1OzsvToTiyFhdgTKKxDPg+Mpb0NAGHfilpAqCqBPc1ILO39
Y4Iw+Byaxqcx3vgx2hzkBrBzCx3XDSgb1x4cxAdiUTxlicCMbmRAPR0B0j6STNrdV/RIQMZCej2y
eLKhlH75W5mIsKJ482FzUCbBckguMywM2CleefsyK44S3k2gMO983iBoS+8fBZ4PcdPotnKNpNsu
0N7m8u3J8xrO3MERXZmoK907b8MkS8xSSlY5UHUEkJDmDGFwqO+mtAgGVs5+V4D9EzmNLyf5GeEC
2pl5ZsZTPRbmwl+0mHSG6iOzxBwVLp7pNKdkoRRQEmIL3PBpRVw3FF2et7vvV7W0+81G4xjfjCUV
yIUXj9cgMsHbI5M6yj915KsB1BQ/9YirXflouozgdiiK9x1gOg/wvUjiKMAQrGbzf7dxa5tk4cK4
/qc+C80nQhTwn+3A7vNCY3s+lKysK0Famby+/CwKSlj5fItEsa1l7Ypp8OL6fQJ94J/2k8qiPQ3Y
95pfIS6cqciYXhVHSGTv/qjtAxGC0mZuTGAzif1T/chKmbOAY+Ahe1ir+HicRLptPWLrBcNP6tv8
Mm1pq/UcDsrdrB6YMT1y9E9lw70RfI1foBZBcUrKXC5D/IaDthWpfYTrYI8S7xwerp0jmR/H8iVf
v7iC2Cg+rQD7wyD6g7TnqTWn4Qb+pTbfP+Xg8647+OZC70SXvLJEnbayfi9JqPaWVpxpJxCn2otg
7E8mKtKxDH2ty+2pzb5OJANCCJHxJH4bdrYz12t7o5aUIF88RRkON0e7RWaykOIlIv6WspcKDKsM
0WeEecXbRDID2f1eD45prZC+E0aElKgw0IILLkGEqsA2XYHGj/o5P+EodWnXiZfLctVFuBjjqzi5
YNWvm42FpFjC0Pl6eegbnhgE3hd/JQDCcIcBXDjomh5IK01bDGDo5bKvppZ5t7UXG7RR1vWEAVTB
L4Typbu8nyNfrMHIGpq3XbdAXaNzCKp1EDymZQ1a6DxjNGq2Gtp0jjEp2pZ1wJQABxW7KoLqd1C3
LG7sS6GMEdTmGt6K8OCPolLLAYSZEtwJFt0BVm2uEKEvjIKjPj0684lrz/EVJ9N39FD/yux0k8S/
++wik4F8y+udAR2xtRMaoeFRL+fq12Mf7r+Sd5L//QHL4jcaEFyeiEZFDhV8BDswl9zYmHCrgD45
imPVhZpyPF6+UreEFm7Q/f4dbkWXxSqoBXL9KIGAoTR5brNZbWnNeBL/GxaVW4A4eLdPw9SVZ0hu
Why/3pZizNPOAc3KaUGZkpUt0OsIUkpKDMuwSaRWhudgB0EZOfe1WiwSLooW4Roh8LR02BMcW5yK
CxxWwsJszGM8XARotGiMrYeY8jK9iGBcuuI6hG8a1bjydXrXBsQyFhcuzhUS1jA9h52xcNuwuQ6L
qUbi3UR+Ri3Z2QUHym/RNd0g/WsjyHbdZTvJSKQkWhBfwEAri86SyX2FhZ9zUl9sWwGTIEsplK+N
/6Vz+vi/3lQ3P0++NqeMjke9qIBVNWLngdlV6WsBfSksvtEM5YwEwa7LrFVTj9HOUUyXnpnPoIhl
8nJ/6wsQ5Q94TRrVo7kUF5Ket2BfG9WM59VFCXrHh3IRvZYzeZmfx3IvLpx93XNhcx2PUIhq+PRm
UKeMwYfqzP3r0H2wp3Lk2o4QZwRA4d1Pus6mtbuD38yzuyfe5inSasojNPv88kZhvmQgkTEIvgYD
rduhR/LsMeCoCTRfjlc4lqSMcLltXSi/wlrhMmijstEXOVEykEA7E96LPZb3C8ICvlEstnX/cpc7
cI9DDP6+OcQG6KdQOuOyqpInbya75nDMyOC7IZGuR+gJxXSXw7Oz/8jN9v5MHU22uIc6eteh+c5N
qBPZFzGIqBseHCm9me7aeAi6EAb+ZfTQeB3ZFzcH1+9LO/obUtfIUrjR24M5Bcl7eGHknZjBXjJx
ZBTbyWAR9AwULdmgNP1icDRaOQNDSet2760pQiSPMotEjCaVtfjDHjQ8g67pfa/IKPDl7GgAb4my
wlPmeCSTzvN1Awt7G3/GaBXraKm/zLZnvy6DE8GWmHqCDS0GB/Lt00OueYyyq1HTUieVeI0L/evx
BCSzE67jnsKyER5Ml/i6xLqxrkLIs+8MzaRG1NcwIxAQGD3u3hekcG7n5M8PfwPS9sSnk/3E1QYj
q5OF/XngDuTcjr85mlKBrHuO8J6Qg6kMXMMV4kwSR+8YnaNuj4DXlIs8taYickJu9Bzv3EmXv2k5
Nhl6KAAOBI3UqgZpjVA9tN3+2lMGLtSjywo9M6LEDlODZcxogSls2G9Gay+wxNH0OJwVxESINrre
L2MuxWns4sYTJAg5bAbHAUxp1ixZsVUEQAU42q0f1CK1vEIXB4nttHQ32qJIpBudRLPJtWbBoPzx
+SG2GS3AqVKOD1gMWqYV0EjRAN5HynptMdnc5+8hB5Nkk4ZkIidFfR+Om4X1gyngLPxCRrSsvyhC
52BwfoSNe9US5+g07ZhO5OlQW/i0BL+r+9jJJ7D6+ybkfitBbwXWGUdWKyQWYmMs/GSnBVrTtZgK
YtK1bsOz8MgMrZu6CdD5psYDyn2IvFl27REfjA8Vj1I8TadtkBZmGysdsJinFxKxUbIHlAEWZZkw
l/6eOVSsmdl1IbVz2yXYiANXf6PbfyXoZXIUTEdk0T1EqFwFqzdDEToNiHUme7H6CIgMb0aSvDDK
A0IbLeR57ldEIGpbZJ8//shbW8Gvd7oZKfqckyfQLaGCsqBLI3HyipzUpKKAz9VGMrt15iCwDJPp
vZyZ14WVC7JYC/iQqh+vvMwQ5WL4HjDmuwP9aKH01vnapHH+oHUdDJLguhqJnJO71TnEjwqYCQRF
Qu7XfvdKcwpgMUD2SUBo8x5bAr53ztZD3KmSynwC9Q8LxMWrkPVRuhNArE1RjioB28uoZw87UUvW
kO0g+Y7+H2wwpIzD40SS1JzC0PZ17xZ1rT+Ad0eM7K19MG/Ic09S2UzM+F3lGlLruJq+wqpcZoeo
4GbqSoL6EJN7v/TRKV2LELr6EXlie2Je/vUoqBLdZijQlvrU2XMhfyDS0ris4qimkNhu5rv0NG00
UeK0pwPJACYe+T8/OazraFwy5moDdRDJYJsToNvQJDXE9CIdlFbHirBdt1Bm5v26ghaU1+Ly5Rql
rbWnllopQnFhans8RnV+8+4jeB7+BHiSPDN/Bwmq/cn5mbtV+kh8UzIG7SIq2MMQGRCdmUyPsNr6
RxAjMokZgZ86nX0o5m2SOXx3f/Q+flLKVygFqRIREVHCHvvRjoeWn3fjHyWNastccIZugKcVlfGo
I2fpEGZn59HMgmhbGOiuPwV2w6w0BhUSUXv5ISqjgov+VUXpD4jFPbDfL300NJUtKV0FRFhyo1LX
RvwlzQpCz//xAnyIdsQpfHc6CJQh5VFdwb8PIT+ervTAIyqSZ0MwVjOKKrv+ei3AOX6DCP924FxA
3HTIWYV2KMmlRp/HBdPrIJ3ADh7vBdhq2NmRmc+cQyw3+87MzsK6cXIhiBEGVWx70uU0N2N32lP1
4htZ/UrgGK6oZqxC0Y8gavO3kdi/Ev2DEwZWDSPavBLvVv5gbP8VVpelYixTWjFCMeYTR+QN+I07
8W0TNOJcsnXnJmLZ5Lr+NcfXx0Z4V9qBqQyAqSngT8+JztmOSEYSwNP1r8AWvlQHOfpuNr97JH4a
Cba9Aoj7YzzSVASSKaL8DYxgWz7mjbaO7Z7FpGvaf3DX6WElWZiH1Er9zI64PJELD6doC0HI64RL
Kz/NEFXXmtnOtU3I+nXU31yDgm/OC+2x35jViStTMS1Tr0a2uX1/MArUM1apkX2nYarcValrLmBM
+Ggz/vF0K/T8w2nvSpI3Qhi++4XAnkTb2Jo2XZH3X8kF2666vJq+MQ3lLa4VlKXalPWrdylOJysN
HKAmju4K9GsKDCvL6pysJ7AcN1aH3qsEu6+gwkm1gwpJ/q+h/eTcmJ1WBgWY/blaHSVJ/0Ayx0OY
pAXyhRW1hRKF4IShRcXZxLjJ7M4LUX3KdWiH4Q6nB2csiP24c/mdQri8RtCta2nB/fZdymc//1et
CB+USF4UzgVZS6IcU2GHAhmFK+7o5S9sGFwOCLPMrUOeEcD/NR5Jj/+B4Wup/BpoYQ6HHUq22Saj
kWrTlKUxYttycTUeZDhxMOXErie4JJFGxKz3ML8K3uIiuXQq7pLx5atGv6NaRh5ZpwbPBRqIOCIT
2e2SBuUVvROKypGLXgI5NS1CbxaRixWjcrVv0ereqjol3+I5b2DsXIf3f78QVKIFTauRq3UZKo5a
nn0a79L3rd1j/uFyD1thfHtMlqx1CM6Y4BiLrWCBOmkNojwRG0KcIm2ZkkfHCZ+WBuE4GMmhFoek
FqvwJ1N1d3YR/wdEIW2rh1E0IWptka/j9HCraTqp2eM8DecUteluoXMDV5vlPKfsSs96mD93Xfgr
hZ78f8IfVxf6uUm8UoRb4G3R/pZn54eOgMl8kcGuqEFmVe9ph4VDFlYdJ8lqsjZPfVipDhjGEyD1
a4xn/654vWW0lOjTsQyy7kswA0LGyFuwceQSObsO7S6qt6gzxbE22ceJYYgWhQkI4afHFptDDi0J
sjMdtvpZtV53xLDL1SljrEWLlmnkZ7Efqfiysgno0XTrBEP0+KSON4/I6KFcHjF9NTnfSuoZmjwG
Cxn75DpgZrvNpeBLuKcLLaXDTg4bqetnPL+acc3o7KdnU0uEi2Xg8OKdY4LP5PKkral+lKOz/Et2
UZ4QsnmrT074XVH2smN9ICPrY1n8i85izcdrdYwxTFbl+id95LVVL7amR1p2IjiUEEigm+h2lLU4
+aK0AMIzQWl8coGLeBhwbbPzwWA6BnImaQgRfyuYiDn4YkDQueArkdnrl066R5hI6j7K7yRFgX7E
obzQD4Ct5YCZU81InHCOAk+RynZ9pHgauzSyDcWuDH7U7UiVb/SoDT8A5bNXH/Yu5BaVAIrYYxMt
9SSePTRgyH2hW5AEDxGgjPHKdWNqxzjsCucJxrIOKvvkhAoUhyZdQlQ3ygHZr3DWYZpRAXdRzUvU
T6u2nvvtCqiOTAXbfm0owKioj9ByKWTvGcPhM8BdFn/8seaA/ElT7Vf7bsPpCKhhZOxmVViKwwat
UZsFC4Mrh4Ws93+eM3El10bv94o1nv4XxjEALOaUBF6NjDHkFLci6BHKSEjgXzNfrp3W/BT47z3W
5tZcDpOF/Dh6inNYEbBv3j/al118orabAl3hHOad/Mp1xFzCwtuuhcDDoze26JmGcgIL66VTlvfi
RhgFZJz/bmH4eZ6Xi1c0NujFtGK2rzkdLbEOURN8a1nD+BI2qgqRsEK19Q7/S5ALpEm29ERDyZ7J
KhD1dk8UvckyuPTNzjqu3gNnuVFifbbfSowbzpkIvEij15pUKHAXcER7Z066Nenup9MDM856+dat
P+wvObAVi56+xQ7e9jisCixEkqG9XvLJJ3pW5oMQGoXG0IDHGPmzXi0QeRpOFivD6T2s2c+AhY4X
A9muSGYykU2jvE+NsN1q7/sA5ulY0ZXC0+7NJyeWh4i/8rzPjbdOFTPwOjHznaqaCM4qI4zLVaaO
/4utkk/ziazCbun2iwW8LeQrjFbZQ3MkbIQyjuW2o6mA1Qv4uPT37riNzkwGajIkl8gFEmyolKrB
yO7qXwzhoMQq2bKavjPLIgYSgTuq6VMXy/hlS+ZC3A9MiUtW3teTjUXIQ76FQs7OR78mGiGqC5VV
eUyyt/SGDFTG2/4C8ARQ5WtdLThFDs/BgIEeVr4x67baF2fYYac6RwuXufAHNBfVTBDGp2sUVDCg
pavmv82uK9nvUH11LtqvQu4Qa/CpXs7JhUFCUECwmVDaX+wfdfEWa33QVmhldp6r/LDrx3qDKkQv
frMsXrktXh37hvZm6/EsugKPHTeWndMJyfFCWYX0pIub1KPeKYHrkuhwDyOb00J6bnkYsn3+NPGW
VfnaPpGVDSVQNBZobQuRNDOVrK10uTsr3UMICjeDZTNzz4iQspKGZe8rpQgM294+j/wT2q8JGZ6O
Y429TtTBKHsB/LWUyg2QyoiUaMndWezNkVdZIXvii6xhxMRuRd/WLOGxo5fDp5idjHW/NKeYNGBV
zCpXLSdLPcjP8CeSnObj8X/knBYjvaN+X50OwteUEjX05IR8Bnpk/aYajBIdCUmiWeyTTDMygFcJ
7uWYX/7dIYSWEX6FYfQDf1gDIAAcLgOvjZUr5ikLxtXHHJDRIej2mm/kCjXWJa2mDW/a5Kj2uRut
Rlh+At3teI4+ca9wB3hkZMEc5DhLpiWNs6HlJzoKgU1H9DJyzuRXHcClVxsVG7sRoJyoXAj6tvb4
Mh/bgPzc0IIQZU5vzMzPEywQaE144UF5Znlq2E9jqFyd/c8VCOPTY/ROJ2XBeSTiylJudWsIatyx
vFu/MsHVlrkYEnz6nXvENZvkZZ8WIziPYSoU46KcJO/H2zLq+DqtqQx8cG8zT6ib184MwEt/n7Ed
d4h0JNH+qJaIn5OM/cDybX4CDWWSBDEFLD7eHW84p5XQmolTkfiB5j9TaAnIMSyR6pHIylbvkaT8
Ijl9ZzNqGgTU033s4mIN8aHh+5tXmiXv71eRHeGq93A/3L9C9sPxoTQweIbOMcSId1v9uRMsHJOs
rFYvL8p1dFafsJpmjkUIjVNqVoUvh4fC585AHxQUrUta0FNPjpRo+IIdOpj/4CRAXv4qS1SUNPMs
G55ngSHrVXcsaBjRgPEK5aT9MbSz2xth9wGJEkd9JnwQyXQ96T6wNdx5UGreCw5SasgX4E1Qc8Rq
eoSamOMBYQIKbKFvY7J9tM5CRkNplD3frFAIJXisG60SnqaKA4pDA3fmE843OWVeCo3jULjHY53a
CgmbmnuzRiIpT2VyiJL2vFDkUI7HSJ8e/psrw6hGGJKbeQrS2pJA/pxlDApNRswbRby6aO+D6wWE
crQkwYYuqTwlYpwNGLxcOS+jr5heM+0Ow3rwEG7Y4/r4zt/8K9nkzDhxSFGosal9GzqXvnl7oxuD
Y8DHDh7FIfLgOzy8SYTrMzhoZJ+IKnNjw5RF70Kl5cE9Rf9hsRjWl0phhRrBbg23+pRnI7K6hIEJ
67zLdQcz73/lAxgiGeMqiixNdUyEhDyoU0rqbzv5y/z1SAI8MjfExteAr3NSmkpC+X11zlQN9nOy
Suo7fOjChVeSddhSY/GmsPQLKi0HPBqD8dHyi2Z23s2/4hch5nurUfilNhQSMqvE7CvtwgEmyHqc
JBAsUtJfxZ7vqlTgCT6REQeR49Nt/TucHGfBj8kErjg6px7hEozqFsWjwDTz261dnVVwh8hpiYhp
HEcWZuZoKkfxUTIGLf6HCt+xXZc/teyAn74qmKbkLF1ArQZsLo3ZA6sCiTQRtDvUvIVP8VYnI1Qi
b4uOzrM2QTP//bbw8Dl9Hjb1bawTsBo3f3Wcj+W8Rgg/gbZm+T6Y3rUot/Yc3HdlZgoTg7ItmAmW
n/XfyVL6hRYihweMJZ+xJ35Ggq+LD7AMFbRKGa5gBCWAw35v8a+R1XPFTSz+6bdv3G+OsbBkUv9z
DPm6boV0dhE1k6xbf3G01g44yojSR1zg/xSUtxrT4n2AbN2EJwPbRsPMu6LBEb1n+pE3gYqkE3KW
Y4kSwMSGrAitAEhmzakvHUGQNLX1Rm2zDz0aRNuPmODXv3LIkpRhDbVPu7EPIm4BQOnCvgnN1r2n
3ubA4TlAN3TtQB277qAy/rqjdKNoUy+LkwZOxJz9OwsiAiyaMGxclxdRPXWV/k5+bb3OajDvdX9T
dK84Ie3/EArRAJkixYJJPbVRSqTz6DCetQtoJsMYSxgVtGqLsn1FEsZZD80t5OA2c8NCP90uqUKP
/BNf1SBOLG8/GTi+och9kCy5UHzNbUGfteeQVWTcq1aVDq4JPXYW+8ujQDzhVBF2L++zra2j/5Ag
woSks+NKmb1/NqdRKrIWHdeUuui9iXUF0Hz+w8JnxIRxrhQM4ADZk8g314g96qGCChARwEv/PWnK
oop5RrZjikXhW2dYsrt7mlE+IR1Q+1BPLMG16C7O4v+98Z3eJR6H5l/epFjaEekTOUilLLp605V9
Oe2oVirpOAw6FamDYht6DyUhYcTFP9bNOK76TduOEAdoj9IKu+aw3ej/lQkuK2GLkkma3zlJtXOA
Hh6U2yanUBSO/8Pb/oo8fs9187A6Ne6Cp68IOJdws5ZT7x8aF650YNDRW4Fkdz1VrH2Ra+RmK5xG
DaO/1P0G7gmu2PhYvbbmVdtH6UaELRB1FLE/EMQjpYR0rXwAv0IH4+Wlph9qqhdtWTLnGzvJDYxc
aJwCDktTIOr+g9QDbRSbKUg2qcHAapFlV9I5uVskXDk3+egfOBgQlerxJLbMjMKYQ7Xe3n23sshH
+sxqC0rHIdU/7COVleQ0Nf4nlzLRuRITknlD+fhMXP3VugVC9O9n2HvOM5hDqDBnQn/yxrYs1g8t
S2m5ze52UDQSz2tNTfv/+WRwhURrBB87YY21kxTbWGA4GXQA4iXwD6j6Q453vzGIFjxJEoQ1zYu+
8ybo2DGkeaTlmD7Bn8UqamVFijmPq5Zw8w41txj3r6wxp7UrDyS22A1poNsc+thAjVXa5XWCIXYX
w7pDbXt8RERmsMq40KFtR/izMoN2UwTnMOwF45wcbYdsvhwKq11meP10ZhzuUN8j4mtGjamRBpGJ
AunZYxmllmvzCbfytxEQUD0mRUnZq1ahEUU4zb55J5Mxp4PFVVPVfnSRXrQDXwisYb41yWDu16Xa
a01LW7IOU+KWB5DFJ9ZGPW2nTsCDwUsxWpnB7niJNME5S4KixQZEG1JCQKg1C8DnQaXOn9ZNGg0D
YCscDBrJiSuW2LIKWuuCmV7xVyMgJ5tmMTX5COWNBlwTPSvxz1Y7DLAy15PQBI19Lv4Wnt2qppnv
VuOt8OsY4ydEw/+GEOqwwHq57H85w3I4r9p4Y1K2UhBDonrtMiST34XvsRWQCZggQJhHVvayFdoQ
dYHVY+bBepilZ9kmo30gDxpvtIzcr7XCkKxX1sBSdWLPHn6Lz0CUDplWLDtBUbuIE90KLycw6aMT
IV3ZoSxOAI8smYCdHwsE+7XLBEMYW3XEDwZS22/41T4TUkdHQf8p+SrJYR/epCi2RWFkAA3Hqc57
fs7OW/NroJd4zoSqg4UXFxhmeMv8K8sheVpLkgVBctXfQxkyyVYYi0/r8S3FVzF8DHXrqzt47AR1
H4R6SRtXkWxA8lCXjJCj9Ogb03ZQ6T2YdYhUqNq/4OwUkCuKM4yXYrvMvDaqF2a/lIn/ybonfrIf
Oh+WURGMPwGTE2A+VH+Mp0J2cGs3MKIrx5sDGc0Hg50E+yHw3LkiQgYYoYnqloH/IiZOQSrnx74z
M7GnHJh5hRqaiwzKM3z/kqni/wkejuKGzn5rIqosascnKUy7jtrsUT8yMP6fJ4D4Zwvk9fwahhYm
F204oBb46B4TSOlggo1nyBp2WeFkUFm5hhJDeTUS8oqR+XcxijptEWJzh3QvCsnYFeeBu2FtR82C
aDNzMZGgJ7tq/FkQtSzROIv9DqYBf5/tGO2+RyObBW8+sB6QdtnE1wdkQejHYAUIAL4o5GkjaEk9
BT1ysrxnQk8LV7du5e78JagIb7RJhGxDo1RZUorHNFWjIcGS7yAZzCWX9g3b0Nmo2Vb3QyNabms6
AUkGvFgfFd6TRUYWrBYaTtdYeYP/3yothGwSWNZuhYEcNnDtO2Dpvkem4GC6g00Lcuuf8408/0YK
l02aTEC4BAp/8vOvP9dTkVtg85J/Rk6W3rcX9gl1UDxZ+UP1BIEH802bk/o1AaWGmsOWQmm36Rio
MJd5qawvw8FIL1F3nBqCRbF1TtKiG5LU+yIyrHNZChReazGw/xxLCoKpoyvXi8R+VUIqdYm6CVil
BCRUaxRZ3f6ANo3YiddRCI39ubzDFoTQcJZuiEtp3IFkr9lGztRmiR8ZT0wHY4afTC4yuaD8eoLb
zCQo44OVQn+CCQ2pr3/UnwDL4p4FPKTzQkB2G2Ny1wd3a9jUJsEn1FzxHUh8Vv31q0E0VT3d4kn/
ZwmK8rxYR/nsp+QlzyQlkr8dBjbi36FYFVI/QCQdvzXQq6Ji6NYYaqkGpoesC6Tj+uqa3rsTO2R7
gYUHlDnk5fGtBycdLTeguBotqSjzzJSc4FCCuuGCIJFGJ0OOY0uskl5fAa3/5n2x6fvjJG9rlHh5
+cut1qj6aCd49Mp6Xg2dELD+9ebIJWo0jKeUGZ+DFzQv5cXPa/1fvv1k+7vph5E+eZTszkTKB68D
A4aYzIGCQSQzJM3LMHhOvTdlEvB0aA+OJWMpPgDc1Pl4vFOA6Cs1oNT8TF0mmpgiYRN7JLJ7SbuP
A3ShPURb1vXHs8sfymIuZu9uW4Yeb/SnAID1f6T8YPezBfHYuUE8tHQKeFjwaryResVWIHX0oFml
x7G2OUUR+Dpqyz9dH9ERjuWSO4GeC8iDrhKoPWowZNZQQvr/oJoZ0X7jJ72o9cCU1kVR6WvhPe9x
thf17oajx5uBVpeDRefW1SrGOjVH0oCg6/EEebdUxNb13ooaeQkZbKz6mV5uCOcLVodRPiDh77eL
DTgJqHkqgn16CMDyXLNXyR1vXEd6Xp5J+ucDTMhvkpNRIIv57W7cY8ckFzODiftEdlbnnBLqqo0w
7KHOIrmh4ivqJ0PKMhBUbG6BfV8ELk+HN7wyYJ1j69foWR4y8idqIIAH1vDqap4n48qHS/XH8vO9
ubrRY0MdnlwZJFhK+VaqfLLTCZG4EBW6KpZn2cg+xaQSw9ZkwXaHBEeQFgDvyarCX8j5XV5e33dV
L94ICpbfdR2rxyvNMf56QGo12yepIcguhUYPLz58IP8D8EhQiaa9TyFDevuBSeSB7WdzJ+oPdsdc
36z25ZOwd9b076luzPaYZMQj/538Iv2W4zkIojp+4jP6WxYlG0/8oX5ufbcaZeTEeu24gKmdsnHH
hA7OFln4M9Y0sDGoOj5qm/yXcGyfPylThCdznBI2oC540Xu+Lys6xPnCSYolPpyOtx+yGKFFPULE
DqYfkRXKgfgokojIOzABKUOM20YWev8SWWkqq7t5U2g27EiKDnTZi1HLCv+Sefuj7AgBNZcjXrj6
gQtT3kMkTDTxs41XAclclngL/6y79bYXaTdDj4zoFtRoIaraA+Kq0XB8tX3nO2c8W5sJR/nf16iy
nHIngOfRO5lAdbniwVUFSDWEIWyqsxR8BxHZl4lYtdihIxpGXD10NKoDq2n7HNuCOETwgs1qMMAh
+8shm9tQB94jVV1/bcvYNMTLw2PuyYVFaZrp5Ov1U9YrKjK1er6Y6D+YCFk7WwGyOKNp+lE2Q/pJ
6iMq01nRU0lh7kd9R+7Qf0X4f9t9Rky3y9TCTosseSkwPPuiVcqyJmU4pAJWUDT4k0grIbzmTCD3
/aA/9zr0mBPaKDjnzcZh7Bpm1A6wgxQTDqxFKb6CXo81Hkykxep7AsuEcL4SyOd1mF7IxkeNVdkV
4uM7x4VauriH12IzqUa1KEq9k3UHXvFRRgRsiJiBbn+E8HWw2fFfNcx4PiY1hAoC5KeSmbAA56tW
pv3Lnq0r+Im/PdQsFI9cYqiPJW2cxlJkTHnXF/I0TYlPZLGfkflpiOVXEm/bgSR56UUTQ1XVsEqR
5JEJEupsU7/nMI0UMah6B2XkIEo/aj4aWddXKGB90HAAnfj1x1VpV+KukSRnlNMkBtc/NJoBVhpN
y5uiRISZH4LFTK083jxSMqkgSQIxMNG9YLxB0jTkRP0F58oJaoDEF+ZspVnawXjHi9xmLEZ5y2BT
7s1f4gRH9oqzvJ38r7YS3TbsMT3aGQ1vuZkL/eNY1w+RhwZVs2EZv82PPG/c845xcDIjRHiIKQKo
l2bb4hdMfPVK2EqSSFIGui229J6vErbBvWU3iVx9pOY26ZUvQFjpjVhFv3jdRFl8rpbxOHpvlZws
iqWJJxIW6QXN3AnMZMO30MaG3jmLhk/ljsfau1yWGjnK/6m4HLJsFjOa++Hu4N5u3clzi1ZLsXvJ
Elqtw5d8W+kTgPIEdSbSKqzHT/RIhlT+rXk1BTkqEVvPpt7OUaxGyBYwh+St0F5Q0lyfzoTL6Mwc
QgDhItS3dRr6vA+8BsrewYcUwu/hhOUO3xBtu76NRyok1+j5MoquNMF9xy/90zY7oVMZwE4UL1fT
3ON0st4IyWewKJZU00HvsXERKagBlBRvF5WjzSqlp9zaxaz+RFiUGgmPb3U3iG0nKxWgjMpQdjFf
RISxattLhipc6JYQKzmUp2uTBiLAyhzINUTPvjoirv5kpUBCpu/qKPmYZityc3dKiJ/T8vQL/hTZ
Jaf2lSMSSv4zl4S04tIPToHCf9LiVTvCxahEmIsPI6j8KdQesQmmqhZ65rdys+rf7E3kxpD6+gHo
DQe998YLtf9HekEptFHqHRUkEG6KPvhrpEuQx6TPZIXaBYq08OiiMUriv6vsofy8zDY4RKcK2/mw
ZE4Ijp9/sCCP0I4GheFBVFC/eHlmj6+drqPotS1dlbfMmx+bTUS6VRv3uISz6P8S/222FigCg93y
iisVsn1gAWQzopzT2MKcXPgHa7CHbJTNDzch98N9/VoMkZoij9JNfEPhK7NELrbV2kUBVtmrOeHB
9LTpTdfnMiaRmJAAp6YbObDQlHVD7xGvGQ+o4vTPbNABy4kIumQref/ZeAP6+LhPsebZAZ8DP1cr
YtyjKPt+Q97nnwvcMyJ3hCDEXXwcPVgSORMtwpky0csSPhGEFm7hy2LNmdpPfZ0rc1pRXfwUX9xH
QVQQs7JfrTraki1rrkgFKmePGQPuQbPtzUB3WTpU64QXp47NWXr/9E89MklXt8i8h54PjL5+hHeU
MxWnk90OM7DwtgSOepXLJxpnvShGPFSyvNVEx1A32jwji6xpQPFrWd2slIXOX5zqna6MzsEO+bMy
SBbBqghG2S74IvhU8UGbNNVAnuaP1ZVvFbCxDMfBh7xb5Lo8Jggmwtl7QOhpCWhjXoOIfl3YYShh
dV9Fr8+qv57vvPCEv6v+gsgnzRQ7OB9t+vurAYHDh031feClyEtik0FyAADdtQNTf2XCDMmqV7Fb
gmbmwgjbJX5C99pjDw3274Mf/51VDahwFtTJkKYH6w/26ViLlmKUqt1xzkX65hVyIeGEjWbwkoZ1
nMbTWZnt+2oWCN8oOYM//+ZSVEjDr796gwkph9Fzpvz0ExhiZH/VMvOvvGU2DezsobdMpH1VZq5j
9wWKn4vd+bEoiSU9otvzEglpk9om/W8F6aaXqD+P6+2Kap255T0tCHP8Am63/q93cYJgMgUIdYea
GRa01DJyXYId6pCNLkNstHOYuFhClTbDmS8spyIgObfvOvczfBhlMffv3FK3P0Vp/1WUCswJ30cP
xsFAXY8JuBo8dU1wz3FKqQOXb/PQYOxUC5KYcNWMpCk3Tg0ZfwWSgnacXfLtTAuBeOhjI1vZ9awQ
wXdaUIB6bHDG/H7ogBGcUKNRxDtG44qMmcYgf9ABLH+p0/M6noCArhVgqDWLLtj7ThlC72dtQYbP
tuDiqmTw1F8W4xJo/ZV1vtcJwx7GdlqQ9+Gm6a6XD5jYFcT3lhWWq/j3VOSJxEx8FyA7L20v1Js6
llDL9sAFKLBBd7eSOAF80pENI6KL0Q10joESTXbqFqhjkoDktHSmwYUgc8NulGVhz1XQCNLCxfiz
ChETn+TBrvTE15gL28ZQMpeG1s+fPqnMggYz1yQpgwG4mFfkPfhzxhiNQlqJ4iD24mxAb0ylWK8g
UEu9IX+4khQw4VBaa2SFDxDmTtPNhXNrOcWNlsRUGyB3UMdN2oyv6sDcvEbfpAZry6MwV++z+BP5
XZ5RJBnMvRBwt2MmthBcVqx6EfIyEh1IgnklCwD/GxHg+A4K3fW53RbHf/Fn9FFbT8C77hyM9+vb
BQea+lHTdo/LrQ0EeW0MY557jHfHJY0VWj0RONHN5LwNxDTs+SOCkBKsWUy2ADDZJJvUnqSo2/Sp
3S+eaKAeH35wTniRfeQS9OQqEdJ8KIvF+rMD2iHCBzkhlKs9gun/Say9Zg/zWC2DfZt6BxMLWDhV
fvh3oJ5OM8LMCedEMmAlUsh5qqFnUF17iKxQk5phtbl3ig4JgOIJ7wBthsEensimQhqgHMlsPDCT
YHIS0wKJlkMS967XdABOgEQasstZ8v7dN2xOJjRpxVNYxIhW71YDcPMQ+vmyvExwPU10OU8ysgr9
h9q6e1j2Z6vF+XnJEmoLDTphyXo1mDAw3ERDNc+sqcwmNFopkSdQSuktzNw+4a14Vyt8jRr1yZNe
mP0aEoZQl2OwhA5DPl44zwICqfMG7tDzNkFwHG98CyQ9McKs3FVQWUXsDfl+gjrR7KD69m75R+x+
QALLpaevaVxXQR1JneSfXsxD7414pOEXQ27js9uRFpuE1Lz56KXLnPQKpAdR1MK18uKTx59MCHf6
6PBqa0Kc6YSrGx3TTH6Nbp9jnOtQ58VlRGOd/lEsh6/7J/Kp70gMFzkrIaEjoBeiD13qhaRylsMT
C3iVkrwQFY3Wq3aaNSDZtVZ2wuPLLmz7F59BIFyaAIJsz4s01vBIITRsDeNeFWW1v7BR2FyqckA/
LKGSVYezJH0YAcR38JxU14URf/8SSVIBVlnJTlpU05EX86b+m9m6tufhmoIcYyKBC4sAYrZbevmZ
bVoYIzowjzKofMFkJONI1zbJhV3KSamK20z2qeAMSP6dULLgeLSr4O0IPkA0JVNoXFTIzcVjfXTP
25YUNbESt+X0hEK7d37hff2DVMQHbwgf65rCqtJtD5JwAwFDzBMWAOhcdXvny3g0O4umaR80J6MC
xrVl4BxYNrAsb98QYr5W1nUeqTY+g0LBMoIMYtKE14BQ2CfAup3rpaCKFYiIVukaiP7ZgUMu0pVC
aHCgcajxP5KUv8GVxWxRZz7vHgDBlcKGG8C4bJT9dBiD3ERaOqYDDpL9OmJGs2Kg2pBSxynd/qyb
iQjGm6ixM5YJ7M9yobwnXQXxZyU7OuS9l7QCe4FTq27Tc1k7goL0njQGeiq+8mI3KCJ7O6WIZ0Pf
fa36sW9Qb9GGW4eiBHnSJqXdcfpzzeZ2tbajGythLoqtivKE/tpaOsT5Ad+Z+gnfpZQS1FHzaUAE
g3WWf/9Y2TyvTzqLZdp6leITKrXg45Z9Bb25iAg+9yhpyYmX3z08YC8TtCsnL2poH6mwGhhnoIYt
/dq/aOx2hsPrxhx723QJD69CXF82hCaeKMT/SjaI6dzLe2wK2nih/N1niXuR4kq1XBulv2mBnd43
oAechJ1QiJKwLNU4zXOtDLlseyN1swowwr0cBd/jA47kPhqvXaI5SjZb7Rnc2zevr/5sFniG7uoQ
pCr4kchUUyi/We+zrFD1QSb50x/29ZWjcpYy0cJGDkrGEPubabMBz0BmWmsA0K6J2Gi/hQmKlTTp
WIAX9v2E8tfl7wGCH6p67LQMsSO7z2d3xEHNcx3Eyilt8PgdwHb907DFwVChO+cme/eNkgACDIQp
u7tZwsRgxAKiP35C3MpTMo99O3IKyDBh/IXMIETukiDhnNYIKg10xaZEHCJXweXkh9UoxCea1cBA
QZgukG80n1zFGrRA32xYgjjBqSvEquRJZxeJ88Lh1eDqe2cANpdbsGL5AFwozT8M/Q9GGQwqputY
CnkpBVvnRBrUtDSzdzkaFP2Ia3Jp4K0hEO4nG4Yfib6285Bt6bmDKkTfO0yz0BVZxcNFuvmvuprc
R1ckmAPZA6afuDvfqOtXvOOKuk85jk6rcBeH1yOuNFp3d/LCiUouDW5kwKuNP6ALBlHq1Tf73cUs
BR+BzzXUcBirjNNF+F3Uk/PrJIGW8GA6g1owQyhh3O66e4QjIcTA5jH4vCG3Sz/+C+XfNhIXnW4+
ce+6dbf8+x7by/MCcj8H2I1FCDFw+ld4zcoPfoH33SU2LlZhtHEHHXLFkqAcx47FPaiZBQ+F6DuC
4UO7u9iM0tdjEC+JRaiBMYweiaB3h3J/Mt/2EO+3foiIcXiWfJEaP8RvoVbCLRmDKWxGffW2HTJj
1ysuNsq8Wwh7oE9eNDur29ZIAkGLHnB5eUK8ASYQLzGVIrSv+2oBmaWB/4kS/FO4Ah4J6UQqnxJF
xatPTJQxM8brVODWBw0ag6AUiyDCbXSyV8FXGkE1XsrEDVHLpnR6klAJQjbd+X1vLr6OzoHYbZN9
6jYqWJHVj3Nfhue14ykFrIGaEbZY7wDUM+6p6oW4ljXZeq5j9626XGnFdatgnSDBMdRuTU5s5ocR
vtJql6A5dYZhfjZV2UOOM4pe61dJtG1ogEmQCoZWz/yEoF4mSoj/XDnYUMxlWa36x6wFeP8ewqIl
zE8sJSnqvYOJOBBB2QV1o0J+5imXjAD7eS0QZWgcMyOQYboz8gx2VjVeGtdRJw3KmKMw+GXD2XW9
TKeaiPbwDX8WP4mebpPL7RXvMjbNxWTYb8S/xYh2ZIUIeAq118XkstfrPKhKybZ3cGqCKWamxxn5
fM/Jnr/A0iigjc0vXEnfAZSUohT9YUIJgLD31iMlbAWiAo+jRQbVzrMkWMgXjefvV6gd+wds2Deh
sXF5ohcx+x+lrNkjPh3D8skE+aeDh/fOWU6nna0vqcirOdWaXZUcZDEgO8lowzr0WNA/qmV4SnRO
iRJR6f0OBoBKNwpMwjpYreSVP1KtpDeKjCZSctHH2vD2+p0bDetYA8Zof/5XiEedfuM5iBj01hOs
tKd1KPKT1b/XKgwQmduH8ydO07Qdbbiwi+I1JAZ8lBJWt71nR4OZEN0JwUFJxed+h5OI4yuq8IO1
V9BNUF8VvSOc7EXRrFHOZVYEhiUX4nChWLfuKFTdH3TmUZCZJWNTJ+qyLAy+RK66kLYwMZPV9GW9
3l8V2Hny/lj+iwp9lvmE5nmZBUNKUDiXixNtxCjnXydTssk512w33ianW7xD4Fow1R1aODdGaKsL
WT/d0EksJ/Ibv3JgPQbPB4BxpOkwxdiZnJbhNlVNwNvT9YumjyZ6Stsn3Gt4KWcLF+mfuvu7KmJ8
/2x0IUJ3Hyox70Qr/wgcbEZv87A0ubXweDE6OLb6zvZerkQCIeNz93rQt8LH9sooXRtIMTZ5NGWX
0KGmEilhAblRIKKEb2gR1Ha/gBAS2phFwHAFYD8UoxjEw69948osnC5nMOUw4IXJ3aZXVvIcpjt6
w7gelfHvmoWhnPfe3mOJrDeO7nM/Bk8lAqQ9kypsO3FwA6tvd+ooNxKJ7jw8jxNPDvFv6BBIptNh
YEmrHHXODEYqi/E4MXnQ8+uM5/r3Wl01meRTijgW20a2nRAu/2OFJDbyfD7DmmZa8qB7RZvj0mwn
8Cu1WC3JK85ck7OF+XD0kgU3edBDx4ScCVkE0qpkiv1ZLV4xrppp90t8p31XLgJs3vgbQkkd5k46
VKXu+nev6STwjkRF0lIu19OQAOf4VBAoFq9GcsGH+BlmoIYJ+N/KExO6/zwd/Jq4qb5N0xXBnFQY
bTqkfxDk8YQlSMGCynHI6j6mASFkPxxm6yym5qxgUKxrTj8oeXz1T5+gIAMNkE+adB0ChYPbUiWD
1GhO+wGV0iuSiuVhAN9/VTQWuVAQOj1Kbg3s++Eo5bAxWeUBPnYKrlkxAjiTGMvSEPaOzOz8T7Pc
OmXGJY5MVrKEmFyWbFGnKIE23rAGedpgIZBc4Th6BAXCMLf9ntYVP7ZPgHZnb9Jql4lSK2TE76z1
xX73ji1D4/SoGa9QAffZz7MkEyIJh5w5MUOLpBGDn1AV13tAqmIZ2VxKQ7YtCunioYuWiZrmsq1/
FsG+xG9xWtzQbt6h8Z9lmBaawNEvAQWPm1kXiZEgEZhb1uZLkF7OSsfEKMwSpPqhGnOpozEvFe9k
LPxI085bWMGlbIUae+tyYoO+fTG+UrcBwDV9tsiWfP2+E2SVwfg9kPxEupK0pgaWKV11rC8rtley
OX9dForK4rA+7kHBX+jyuVFlBNPvv3bmfzZzJbFQ/cuxnQJaZkZ1Ypj7fum7jSWZ1hLFUy3enFPQ
zOx0xS9EaSofwDhWSgL7xt1GenN2BMPUjAUyzn0+AFeU+mpcfnWnQLuMzm1Ctl8TviuQiG7QYLle
3CbJnREj/miCQw4pzzNfbvJSwhw9GEGQuzbscfn18QRRGwy6q8RnYg5eRGPnSaS4hXiB10gpTmzg
uycrj/O4+pM4X5kMu8jQD4E9d+Fy1wFQZ6qPWGyK3WGYHr5wPJY9wuu5h8REsd1ivXcfXxS9wFMZ
X/2u+doNYusb8siIh6p0Ks3qSKUQOO+LTkEW0lrBeQ/LKG3VyHHEtG7KtqQkpLObImWIzE0LddVZ
PJ0Ro1g82q2Q5AVsBfMJx9wL7iF9Tmrx2NWtUeuIUIInxKrQqmsZmxd6zDSHVSqMLBSZL5l2z0sZ
tZU+tEMnbAfQFIs6zGE3PZD2cftBrELaUNjD42lEpe3uuUpLF4PGVu6SZ7piG9uU0lpjFl1EIJIz
uLx3pOaDE+77QDq/iciry4I2DgjoYnigAO9pVVE9MDEQGMtk/MaIiKZkhbMDQXoeI/ytXl0149b/
DSvvFsy9kXlat9oTka7eu3fE6kqlk3jKXRxoIs17UWrZH96/+u8/ITSya5XYGGzAqZ1Tvcoo3uNw
/MF6ai4RSqQt7jePm2sxp5Znw9K7r42i21AmN02lakR0FW9kM6FU7yJdDG5qpR1Dv6413GoABJEK
9if9zrkbqTK/Nz29ookF/VD4oEu2vn7pn8B5exy/BaKApfdjS+YWRzg7yLd3/Rj92c/UtHuXR3gq
neKgB0jyH82tiFptcvqQ8Q5d1Iue31asEIgbzG8DPUvnc69OAwd9yoGRyDEtJn+cLgd2/X3312SH
Anaozax03e3q88OgLlnWb9EXcGwvL1XHr/bXLRA8tWj2v5FeMwi66GcMTxyC5iZIeKdFLftIw3b5
x3ABVFn2ZWDZq4LtFiGjCPCrpqr4y9WlsQKUq6Z+qasEG2kfhbo/qp0eydHtqh2cjJcEz4FkB3Um
VCenevr3kp93NkRSTjeELa9CqLuUOzcrizReZDa7PxIVq1IV4JjOj953qKMT5Y8ABwXTWTvmQ8HP
muXa05cgkRTxsxfSQlFSzq2IR/JBdlYuuYvSD71nqpJ0STNUPNJ5AybDkvH83Z+emigoUSL1+i5m
hb9YnIjLojjtlxbE3vdy5Dm6XvExIzZ4xsLMgq3DTSxdVidVgxOXgSGDCCw7gsHV/AHpab6FycNa
Kvp9J0a8T3cRCiD76qS7+DZmPUtYeKA39xRUvRE2JMj8WxpYwDNTPkAxR3w2WgVbapdqO/HCGynq
tPhFEqAWr1nZ5l4q3k3JaQk+7qeSpoBL26M2jmhhqnNoHEYgQ10RS2mARZo80TpYHll0RNEwoRIE
oRYoDP2bFQ44s0oVURPEucB5RlbKpREsaVRMXgGss/l0fjtNza7LxfxWc9bUrgTzTEtLUzlS9iI5
riGEW9CuEn+XBar3XXKkVlHkqJSXMMeYHMEUCmCuxJaL2iegHXhpv9VGS5tj3XtLj2Qi3MJPbHbU
+orCz4FL1+qouw9MUBp/RkS8wbAUqsujiCwagKmOpJuWjeZswysH5Exse2JpARiCVDQO0D7+UgGz
t0HuxgQ5u2BX8SG8povUS/2ISO8YB56Ep1IUWBobCrhHjnZ/S7bMlnMwcSEkierXmhsv7KAKL8s0
4ewVqKdsmvjKLye/GHWczXq5nuWVTyl7J995Tq8RpvL/DhyjpQVC/w+vMFj99DpOTiqDVbbnzChl
lJqCDV/gyj18+/rKEH9AwMY88NFzdIPDlMuo7vHskBks66Qfnir2Evmwrz+uvp64wmawN8fdOlY2
Rf02rzIAMf27RY+pOaXx1i++zqUX4qwXelawKlDwDn5KXT2OLnvvKgM1FV3scMd4sZPQeA4wpw6D
suSQ6ESExXgks+meWURfFWQ2Rm7Wdm/YyCSewoC77PL1nCG/N16D2Q3TrKdl8n8Rrnw5VQfiLBzC
8JmF1CAO3sBB9E+7rRBJCtXJd18UZytysqWTmWEFg2sNzYHp8srGNrkxpmf0QD0pI/2K5ATp8egq
susqgq2hIMj/crWJwX+EgIVKTxgzMvjUBbdjPS0dJ7BQc2abZ57djyKHdMaECg6WZsd7SBqFAKI7
kCNYSn6kxEkfNValvU2jtpB1ZbVoN4rnBKn83g9sN8mWeqqlfQKQUJcpzQ9Eu24FwTbUlUNL4wSV
nI27JQZVuIrQXSy2rgMlSzjqB4Y+Gr7jGBiRhnctSb4/P7QSaw0PkWGSwiTEm0tJKZ2BMrwV2Iw+
KBawhpf5i3EDascEEWRUyhm/fQSkIeseDMQ3/vMTckl0sKB/0grXkcY8aHxWdrNZsSf1msM3bll6
mjCb727tLRkF6iVPYEuHgRixOHvr6tnl0SPsxRV/4VMfCUaX9fEHWxSwD8Ozp65+7EKF/Su/Zu+7
QEeCNHWeVj7o6Ao/r6rOrLJhowXctIVlnvgrw8WEcupNvtsoOZtFGHBpLz9BbIrxvE2D2ZEVWprm
0uCGi0qku2cg3PMem6V16g7lD2wCtYI7QsrxLOAzN1BSfeABJxuIG7jEcyBMgMKHAGnyGeBtXiu7
Wsbfrsfj7V3tyvvVIgGFal4DfnS1M2dxPzLUmlKqq2alKmpJoapbFgX8CTvYP8YKiZjdZCEHsWWv
kWYX2mRhiEQwNifNq1MnPmWk9AfbbhSBZTI/Naoon64YBa8YqP+IRxsoTnGq1Vks4IdVcUHzwQeG
+rUdC1oa3Ijx158tVATYDaUZ9vz0eAvFgpQO3AGJQXwsT9kpxOty6m/FmmN6Oaej0WdCfYzoX6C7
YRXr1MNNVbxiaDy+O6YpJeQlh+t8TfyipxRNhfmL3GcmP59S3gaYmtD9b0IiMyou40zpi/LLAgTa
XHtEbLfVayn/nds1Vx0cCchgrDP8jt+QAR33DREfX9rSTRyQUcqKt5x0kn8e7Xmg5jlnndZOU+Ui
xgIlyzhAL2iJPGxZdERl3pdjUsh4P6vhIcBkLTOt9udku9yWXfN65mY51Y86etN4JSG47tQNu9sD
n11QIALCZlUbYWXBk5w3G1cFEl87xB0hkWKrBsgpg6O9S7NobY50q9kBn6EUUubB2FYpDFwAqaIj
+R/cEaqAkq+xUCIM4GmmbYkEfWNtcKAMxDKKlUfu7NAEMtGBO2j7Mekv6ivOVqAEtsVdLIYyAj+c
MOXWEYmVuopQk9yT0IDT55ewSP9FWiJjRZ4fQ1b/VJv1GGt6+4vNB1zEAbZut04XrmbdOdAOPt3+
cjQ1ZMa7Wn37ZMwxq5Kf/H1Pp3uA8WJ8b/AKOADwzxtCs1pZWxlln3HjZgA+bTfY6dsVw5TujWGR
+Ijnc45s9br6EXTnwD1K7lLXDbYE/HFeqDpTfSAYFhSvEzMD/Q0NHAaWCNdgzTLmkUn2ceeWw5Vw
sGbQNhQ3qHem4NOHRMADtiIerCPSJG/zcUQCXNXi1yikIsvp2HgfJ7MonnmW2Wg3FDuVppMZrBLq
lzoaAsmfAY4eLM6y3J6vor75/6jPz9OUkqpr+xycz0+OgfkDkpv2LbPyVG1/76mkHkZ4bkiLc2kx
AaIjvwHJZxU0mXWO6ep3ZKVwkSJpsQyZqbA+YAn1f2rVwxRVNJ/ZLOhp+IDB/sKclfQQAqxiY1TM
ju12BpJ1hP7D+vwY5PuTQr8sDywLnEvDRj514IXsmHAQ+bUv6qlaESHBYEZS6ZwFLbCIjh22p3dP
1Y8uKWUuZG2/ISEWgJmp940Yb4Uw7DKS7wn96M199h/CyA3lpLmQfSP4AGBhYn434jm+1RFWdLyn
IRq/UAFmMz4FxLPz0D0nRp6puUAjmWlVphxP3gK35KUIp8xSRuUTh2u2Y/0b7t+WTD+x9e5/2VUg
Cv3tEcjZoMUldiyyUzevDIPziHKxn240bLacmtHT2Rhqjr8Y+U/AqZJjOmgosEciK6pSiHJJbYHw
Wr2UzVE5UkHNB3YrlH+rzRvre4mN0IPWi9z6nz6rFrWaZhob3aNb5WulMfumMAi2p66b/8EdZefa
XYVSAWf6h4erlPgV6p/kt+FzAyY9rLBKO2DMiMybcSFPBAe3qQKjzmU3mHqx6C1KWrDm0SnXygWo
r53YXDqYP0ZNyq6d1ts3Sg7oQi3pfvsb7BW09RxASW79ISBUr0kUN7Vc9BFA2uA2olijky6+HGVz
7Ji7RgO7WM4psTKlAPnou8yjbTDN9KMw7bLFVBsWYqhSARGuqmaZP/x2aznJd2WdOSzKCQqZif+/
qpnWuA2eZ6GO83/frGPiYX8fywWU7QH7lyR/aaudKboJIzbIT4qu4gWsNCdTQ/wKbxxIl83dJw89
sa8FKuulV5/l7zmSzvIMT+nWHjo/70RMf2OULp/2aPlTNb0gFHxvjKuMU+45gI7drzMo7zhvYVnl
HDaZMPpCdDNIjKGRrEcwpOAEe4zMASfB6fdLsWYhF1b/OHRjGStI4HRJJhMhJ3qxkN9u0EHuHT1o
8hYtz+/MDYNY9HE+4ilrJHU306rCZ7oph1S8KfbOvmQ9/MKrn8m48mm9f5PSbJMXMC82y1e0bzbf
UvTeVfXEN5bmhMpA7iGI6uINmYHyynjEKpruKwI24O0h9Zc6T1pdqK1VGEbuChKuT1hC1QUYzPH2
k7hBrtC2+R5KhOAdnEcPtZf/0dLEfm13e4svTSjvxngz6C3j2azmgWeFH53Kz1Dek0XSYs0TC+BE
pTqRNOySb1D0gm5wsIj6bpwWjofpfiWT8h2i82o8TB+rZZlpW0T/b3k6d+4Q3NxvlStsMf1Q5yjG
QVHIbysgfawGMJETZD1/U8bUnaZVHn0iWJTl4NmjCIfZErKMQN+Ek4tVMWRTVmStbvnk12XtcIqM
4MH3vEyK7/d3HGz2U4Vuh4xsESh+EwnjjaaXxs7Yu1N2llp/ftyD924mCb7QiIsGC5vPQO1JV7+N
s+xGux3aB3QWv20a+34NN9GoWnJ/uxSn5ofhanGYMd5nyHdM8lGkycyueckUM6gJIsN7toqncgkp
U4ClKIv5NkTc8u5bFm7LkMHql2JjgKnj/G83DWvTqt7+oTji3WH3Yl1rC760iz78W3/VqXUSslS1
awuO7ykSKM8A++YztRM3Zv/DlekktaqCb1V7HSy1X8hyMYKmcdDcswfVcxDu7pUYuFzLcMhCPyjq
+lk3MvJpd5PuAdQVZbX2xUSHjtKPHP+4n7bC2WR4vMgAWKpVc7ycSDp6eXv3uktji7lkuHUv4YP4
38Hwk5QqgSlITOSIWfkQHTekhOk9TLIIQYW3LWpTAPmCGfC3hpSkD9lNGM1sa5tJsAGe341c2Xim
BvMtNlEfK8EJEG/ik1+8vyAgqC5m+PIZ77pVEGePlsRv+8Bx2oTYhOr65AG1J8PrUk+EATP7WdVt
MrivGh4ZVy0C1GkX3UEF0or/OxE2QU3i9bXiaeaXPtxthmku3aO17ymarI58i3ss7mlNi/p5p7gn
9jKMR6Lb3JmU38Hc/Rl4eLYTM9GxbeLG4rP1E2WZFqYMDs0a4HX47nu8Izbp1bxZpDWjzVOIdcTl
fSeAwoOjJlXlRBfhLUuSrAQ/uEFTjwmPmNeipwZhIv7IC39TbbqkQZ9DmGTE1zIjZnwQ6yLaaOv3
Y3GOnK4bR6yE35pbkWlb2ccD+Wv/bV6G9r/22JJFxUQQcuafnZO2wWJqnACS6JUjZAKSSO2PHpp4
nMABaXzKwUmn2r+WxkFOqkJTZwfMQGFse4DsYO8H+MpfotZB5w9F0ntwWFwhfFLYTN1TO7jZx306
+d/PQEBe4TyrYTC6g6g30dt9+/usbaTRsd9hkkFIOz7Lre0hQNh4PyWIUAqUELamVztlMJKeDKjU
fmwyLmM9FvlHiWmKTcjwncw+3LTWwORzHdHRT5AH2sDj1S4CeBUfE7i5actRl3oUs+6M9+uco4t4
fRU8evXox/pmq5yb3CnDsrwl+7t2sT5WQUgOPGg2GrkGqGZcgg4DdKAey0C8fPR90oaHMn8xJANh
4VuMm64+HJWX1yg/N96BwBOJ1Tcb99Ag9FBeubrZy5O3JRMUzN9njV669h1rA/Q5eVg0v94oaBQW
RGnCZBt0BbwpVnFiGMci2hZ6XfXq6+A1jwGDdKyBx4pZtU0ObDAJCy+CgGoKO8W2DfZg7fDJQBsG
Taz/+yKkO2ig5WKBS3Sa80ofBJ8A0FM60SUroJkWZGrc59RIiF8Qk/TpL7ectkz42/Odlic9EZ2Y
DwvvK++/Ps0ZuwKZrzxs+CgBItbBpEbnhlju4wvfvYdCszn+oQaI5bjUtLFxQwrekm6/Lp24I7y6
F5+SPj5P9rjA/u8MjQlYLSLG5AW9hR7d6ohMvRi/9hzFiEua86oCYOo5SjBJkxW5txa9S4GfqLn/
a45SMKUD6xj0BfomL4VqQBgLaIs7h4vBV1WJLTW3HMd4e8BXCg8wQmJegDfX6BmtdeAlrSOgWbZR
80aKJpXt8GGyKRxkCaXtHVRfziXiZKESParGXRpQ4EJFcNu+4/SwO6ORDQVPpXLUsq4AY36ffdk9
6Cfh8CyFlIWO6htkqkp8bL++pTH6NQ+DxvGacctMj/2OyTj2MPXUKRNSfUB/NcnuJFGY9IzTqUKr
W/nBmBHJq60DsRCv3r02RX3xy6U9IBJUZrkUG23I9Ua6ZSgRD1oeLUe5Ekh1m/gHV+EUtOBe3EEQ
Mlj5VOWKYqJPiS1UHSIgNOWwzQ17Il+KnGUBV8h58sbRTghXKoT880G+tHm6sfrm9tZcYf/bQMl8
2H/0i420R6JrXnoInBNhVdqI0mWfbRw5r54EtTHTa2KMlQxvQ4O0UA72/qKuSQRj0HNsbIB+0nXu
5jszHbl/0H7wjMQN8fb/UEYK0JkTQmh320jZyAbnKBCe28frYK2cuHzebmvDOfKEGN9HtrJpaDwZ
AxdDwuDKiKIxVWPYD994xT4Nc4kiVLbvMVsuAcrqIZs6PUid8jwTrYcfo1sZl86DUOMyyyCzAg0R
11oc2Xko/h0Ga/homBftjasoxi453IEe4E7pdihSjB049ngvoHl8zHrSluIKiT13hm485EVhvtqJ
vo1mL1MrgQN7Lu92AhE586EJdFomHKMvQSXJETM6b1VRL6hhi1IoKYSm9WBedKeYxtIb4iDxHbBE
EEXbaVFqW8MRdv8SiJplFt04ViJjZnFrOhxPYkKaAdoYEv9RM2oWu9Evv9pH80RabftHPSt+GbNB
B1Gy8R/YCSeGkkW5ijPvPxMm7CjHcZ5uwceaeinmypuDhW5FOcszucZ4fgwrf63vya3U4jU24aDl
4Psk7MZZrKbip4Z9P0IfAlRjEsMYgte310XguDYf9CtW4biWifL9mPX9AXLALy5ScFWd2MlMkyaD
/oUfz1c6u0PiUwuXsOTTr8ku7GVgMHh36cJlkMI9+wqRjQw4Ls+1f3JOo0MF0s0NKiw4aFsofg8A
gVO+OtJ+jkE5IiB5d3J+vtVFjEhT52Jf+vDfhWBgDy9sn87AmYbBZTuFlxRKOBEhaBgwdjCEu00E
3rq85J8wCVue0QFAwXzm8NuuJ0GlXlX8VGzBTbO+a0XGAiduOQfwB15jp8CJVHuORp+/BjfxuJpi
JU3xYID/oKIebkpuQ5QUbirPdiOK0KeB0LPsY2pPp0CGYuN0C98yW5GNlPT+6Y0MlUl64mELl88F
R9j27U1dyJq5E5BTAcrc0rYrEQcu2yVVL7vK2PYThPI/A/evhjDYbs3WRtXgmduJlLk7jpqzL3Dr
HZMzaomUWA3GINTDVGUMcExv7ZDXXuScggtO9n//tECQh1HrKUfaUJqWUf/dwd/qBX5SGt2d6tKG
rFcCllEUy+1go133YmVAT91CDUJz7W1/R9OknMbIkIU22veUzwD0xK/2ulzdxE3/zIi6Xx3B6+28
w8GyXi4ChCaRuviTbgsVKEBrvmwCiQSLrdWIUj+/yQiOXY5p3sYHOfqpq/BUUG2DxhIKaSbf93pe
v0GQWEIRUQ0b6Zh7Jk6m8vgrX/i14K4iWny5UHhIa008TlNlpOtVUTHt+pjSTdIRtTJWzzgBglIo
Lkvc2viIo/pqRzrt2csyWaNzrrFh/SETVso3JcqFDq3WaO3rqFk+m27QdgHDvkw0ZbK8GXmUa7xY
6z4QXNacCLIxgPX6aVL0lKAqGqoRAkV0hvw8AdfwvAR7KJ3ZiRnRrKZGKnMbYbRnI1UaQG5E/tvI
eptMjBD8s2F7oSETXLheqGOsfgHp5mFJbgj3PsXaah+E3micInB4Sk8bXBJLYgf30WYOC9I+BkTt
HGr8IWkAZu8CrR7ZJ8AAwQgjEqsATC2C70dUpuf+lfjEAHeG0rpnEHLi0jxJ8RaOwnXVMxitX/Er
lwrOze9DBAPwWYZjAhrBMeJOKUYI2SMOEGc8hbJGJh+mp1iQ9ooL7tNtNVtXRNd2C4u9dY4OxSzP
fyBZUO5phM6ttU2EgeO37OVyscRYHlsC8Xs0KxDvfMsiarTXIeeDG6cxpgyrlYF00DLI6K5DAnr+
KA/5HasSapakjGIucYdmrqi3xl/gL4yTi5kzg8iXi3D2G3juQzXj5XNpo+yZPF+HEoYgAucr4HWa
xhVOwBIGc52EZ/Y1/Sd+MYeZVeK4DhVioWmIzp1vkrJ3228nY/NxE46t6Xs6ozlp4p/4HbkAomRq
STHGDdxXGZX8WUurGTpg3Cl/U3wLTQIN0iTtlUpWepfSsdXD8Ghj5Xl2zYm97FkzKdmqUadmT/Ra
cH87UvsED/iWlVtsVsOtNWngQOIAc07UwM0iysm5G51LWgSTSqnqjfBzPKgoVhM6rNrE8NPF4Pv0
ykKSzxyS4PbWYHXfh9nwGPQ9lK9i5wMcksdf5pI4ytxogDZabB9YEAQUQW7sieAR/O8CXMo0Ck22
3e3gGRHRMrjKckNCQbZ0TUkMxARNbxMFa4RK7NV3JoQpfAzIlwOqyQVllb/2A08mHpouIg+Fq0Nv
5uHrAklSKcBKw/UYpGPNnPp/6uGr+71Dj3MbyNEse9T7Z5CMDF2Id0XlKs0Xw+5c945TWTi7r+9k
x9+bHXHrK7yJfun/qIdoZAOk3CdP1J63isxnT+1vc7RvWIkT7AS+kPyovxcdJhauKmNbGQcvKH2Z
o3/YGRqlTU50RkIgaw4czFfNyhoTtTzq3hTJRYSM2DLSQEfSF+hWcKpwh1ELRYgwH6+J08sTdstE
FUN0WVk0ALMDc9jAswkRiymWIcIPunWPdm7E/5VM+nbTugue++hrA+2zzdZqHEClf0ZKzU/Ik9rD
velEnwyYzrlDdLjmxYs6gkzr9w5pfOjF6fMtct9bJLtRjB+iWk0Dsw8eE/xEzb5yXenTB6XH+DFH
EYEwNDhV4jSNYMmLddZrtj0A12TtUtuDtzQ1S3ElqNTPGZSIhqWaa6mXaUD8MMsfwgzt9BFQ6Kp9
EdSKVXjNZupIKyiAWF7n8RP0K61WJdM9hlN9RcX1XrmRgdmRnBGtBetnXSNttk/r0S6/wEs7Q/HD
3BUhpanU/nDcY//33mgjhg4ahumISlY+HeoFh5mgf6yh7+VxeIV2mITtOrjR1v74Ye6xWrDHZIdI
SpHaI3XEiHVCgngSOokRqxI23OIZsjDwYQTUDElr+qIJ/byl2DlAnXicf2v8Z4iC8S2bGG/ydIBu
9LgiqH54loaijxhdzBg3SeegOY5Ba8rfx40vnstXfNpx0gNZjIfXj/jzI4KUsvPfiRLtQ6FA4QTy
ubMBJGRjpf+zHnnmjHb8smcBpm/IWAtfQhRARCzGULC5Oz2pdjQ/QT4JWpCQTvnXIyWgOH7TlI0C
mOXnciDPuS8sGn4fjF6D2EPj8hPL9p6/gDfvPux7Sua4u6tby7H0fv6+yFQRA1Ah3MIeIABOtGWx
2ItRXUQjLtq7ZdnvCCpHMutg4RfWSIIUiYZSzTbz4TslSEbzzAqO2mM0m5Q/eMQTvVfpcTKobjb8
re1SrLqMzlQIO2UJOPvWAXWrHvW3rvBBqzhUmttOfQr008Oy1S0S3b9VSsZg9V7teR2JCakz1Xeg
JEWdZT8hnRUG49eYLhU/Rs/GWVlNLXlxI2E92DAj+KGqNkE1p+5Ec4JwFNGElsfKrtxcASs6G0So
M+RPt6+yFMdmNVBO2LIlH6KkZEq9mikntX/IcrHxMobupolib/U79d4ivOMZ3d9BGuTM0ydrTPir
OHYam37m5PeMesfY8m1XZdpSK5UF9Ji/R7KkOBX+Axq5wEdI2TrTZ/1cdLG42lRNw6kjUvY4b2C8
rob/6zkEk6zkjPzqE9A/y+zcV77b4FyLUcPE4fQjQym3MDaHL1VzZo5utB8olx+ywt/FlLvAHdYr
Y7yXZUdGPa4fA+MbDvtSOPGKLLUneNBXvOKrj9JEY/HjBh6AtaU7CEyNr/xMsuOkrpsuJa009wxW
igYqtQkEQKiYZjAko+bqncOuNpdlvBaJZiIhbmUNq0wIyQokPWJMGFdp9Jo70e8XxX+nicgXm/M6
skKFH78ljxTSZz/bofHpt6ztYyVDfSIczK/VAzNvuPXnrD79DdjqJ8qwp5/Iqym7YOn+SVqQkeNO
lU7v9P4ydb/YQdK0iBJU/cvUtZCwXZsVVP/+mooj10oxSugeQA4g72EyV/Z4Cw88Z0oOheB2uMI4
qIlRjmPjymxm0lsC4S6l7JJGNpXY7B5nmOa/IJmgPStGIwzv54TN1Gs2JvF1AqeQ941ieEoOtu/u
gCK3Nb71p/5qd0SkjkOIIwqW/VHfokmV4LRSagASYsPHm/0OmeSHO8zXsTLw1ayYYKIMt4vYQJ+w
vS/urHbvHBo4hKeraVGVK0Fq244E51XEAt+nDVdDnOtkcG4BrrPuPGmnqK5Sgfv2FSijIKBcpIHf
KFUsfDFSWwVmWGJ7SS/doyBTp6I3z9B4F6ANyj4ShT4FiU+1c05ZNyenkek1yvDjTXVn4cSSFzU0
xbzolV4iYBwE32eqLafUaCHrUAXTRW3CWM75QC/ianvH8sM7yI6h+raG06zZeDFtKUcGyU3P46Od
JxONIjcSosXLesoiTpxkp9ErNuoa9bfxF1vP4pZJEctv/asAPxEkQ4klu8i0HBD2oRQ/PUOGwEWQ
xp6gQ3+Z5efmzbnPNWlbGTct4SCe+ti5lPT+a6OJDlxE2IWnz84F1u6H3rHRNmeDMROHxJXSA52s
Pq5CgqleCX1YOeWQr+juLO6oNKK/uMowXmj7kDDaWYAfaJevRObSKpwsBlHryXkhxHOpmYoWBObS
MCeLmCLHHE1YYjq/KYGRfUMHqwqr+YzQYOzVWtrp+VRHT06b5+8lbaQFjIOCA+u31ljeI8n4gWs4
4xcszT2rKwheF92ZV6v4u4nvBO2kplPvgJ99qKSWtZZ3aq1Gg78gZHC/CwYDGDdazEt/yqMYX9WT
wznSMiLC7eqY+8L0TR4v7J1d71xg+1yNgwhyYdUV7UEgIYHC1laAKpfE6uzOLM9p8UoEMby0sTZI
FC4ugegk8gFSUKJJXFYSA9CpKDgpS/6KQmSPTLnwN+dVnYaaG/l2/OKRrAyHibHNcceB9yRJ8Ode
Wvy/t+/hVcmK3YBS9UrgcGF8UXXwrVQ0vOpOBL84daqAyK38AcZsl/x6u4tRqWwcnz5sM5H9tQNr
Tckg7gm+MkH7aG9XoMXnHfrCxYUyneTD0zHs8TMeviI8OyiQhH2UbJxcaflkITxVoeUcqciSaDqK
LDTL9ZjxBCjOdSVPvhIRPKAnqhFsQwWVft0xpGuRtI2nmE6TP3Qhk8pMovw3z0kqamXZlNQs1hys
Tt6Mgbar7cnYKOF4Haa+WpYJo870dw5sjlJ8540WzvvV6My7cGsrAlwZ+MuXTO1jXN2FJgoszimS
2Q8qZazIKOdvntbUWdxsNJzvJLhAU2PnvzmV844p93oYcijLw/pvkD82esSuPG6Nrc1qKk7L8y6h
asFfY8TnZIB1QY+TvIZS2mMld8N196UAUwtDzvEHgTdpe7DbiK+uM2ovlktsjsX5dgkYhAyQXuNL
ZaAdRB8opNuhZylHaHwJOY/NIIy3kf6OdJaEDbzd11rtEfP6cn1pTOy57IrXfdwMrFaXcuF8nVOs
25P+2GJl9UrlpstycXCzETKAG9q1eBlt3NmFiDK54U6Tc09i2Fg3pAJ2xHtPhcckmqGTnfO8A86e
kaICd7z5O23+NYPJXevb2FF6chheKXupnilQbnnVxUk/daUMkTO4vqheuABRfiFyANM8euVUlG1j
w7xYH17THY1ouZiQdfSJbjvKJAtH079st9DDCt/ePx9rbHbhLUwcxEZschq8ZAn3rQNQg0cZwKvj
nwjCNqmhl2eUItoIXgjAejO0R+uqEBbjZhAWFHobiQSiTmV13NFh1If4qt9mVV3b82bQpnqA8QFZ
SRO1E+bw3qKes+o7UlF6saLtRSb4jFvNFj6pvMvX89aiibmvL8r9iE/QSBAindIEIKQB/EgLGeFX
2UKyMtNVgR/b5x58qQZi1Jc/cZYB2lSygwPnSMsKMTJ91flUHM/cD8IPTgoHYqzCScZi2PIa6Cic
1H3zNOxNLAfkHdHoe60iK4H/IhMFvQioezjWFJoRFEfVJ90L5m9+KjUCOaekDvpL6VXvRNSNAESv
cxgitOj6iCxyTD6G/6zBgwiV+nZLtqi0kzsOrXq/9MiL9fF0WOIo6bCj1JBae+/l9n5kGZboNSeg
M+n2Wbn0JMA2s1zOKufPIYaUHvmpk2Ec7EHsJBcEqm0BvUyPdPnSf5UlYtftibbqUUJ827YMCgil
v7lqv36LCeR7u9DHgxgm+kcouWHrY9bArV3+TAg0QRFFCZw/eP7YoYc3xL4d1O3e1U21RBEvUSfX
mzkRSI/t5mMEFRcwhUTmuv9TXMkEL5j/r+OvG+yT94BRJcvEe5yr8KlLSuk9eGo+6uEbMhQyTpme
5xJc6Yy4tpkvJ9DJ22I+zop5cYQwFo/YhyyqJ0Yb+tXKzzCrgw/TJa6nH+1ccA4X0ojyJ++jbj/+
hA87Enc2NT6NQFoD5awVcgxGjrPkoSo+bOnI0ytoFmhh9i7obmkRw2oCre1PZjvymHd0GE1UMw2O
ag+Y3bgzfN4NlutBvni5rRg5jobtECfNThnHLfLOep8wHDrlQ4adSaRKrP43Cidm9gsCy3jvQ1KM
Jzw5R0ClP0NCUZ6uAKizTbH0u22yp7dGOnm09chhUw+Fv/2R1kiE2dQpp3fGGkSKwO+n1YPU0nPp
4KTe8C2hVzwchGmSz/HWr8ZMl61iqqyn2q3GNZdvh61qoVKRnzSPBW2cvxcDXDUNPwbz9ImyftQJ
2JWOrKjGadyvnFm0PPK4vp3caT/y5CPqCrSM3fViB9fG6l4RofVh9Eo2pOBEUkv9D93l5ZHlpIBw
qrN1QRL2d6jdPqVjNmgmjMhOPzaXntm4+NbPz3edltlhTGK7QHs6/W5ulTY74Lblih35+EpNQS1C
GD6+AHRenJwYQmuu32yMFzWn4v+3cWyXzOEiz34aksthWTVa0sGTGRLCN1lkqnWnynjPn/uVzlFV
YyVe8mAyAtP9GOsEOvhT09FzN0ER7QMKAkA6QCwsKH3elRPERUokmS36WMlbpVpP7Eh3wqJxDtI7
4JQYAqaD6LtK7mJ5Nbo812znhCPPf0bcCp8ulwVGFv+JSA98kv8K3CQSotkOZv/FaYQeS/Xm33XX
WZ6uhvXUzO/tvTyIu90MrxRnURILteovT75mz32WjMFFmQALOQU8yDLYzjgjkX/VdM1TiU4iYoOQ
cbz8ebYByxIS9jOLx2PUmeh43jszgk7ZNbm1Qh4UJxdM+dTXX+pNLNp88hFoDMxw5rcuWe7g+jBl
BtASSE7yUbPK7hYlluK9WvAIOkgTVQFGTWauEYUEVRyGHyqKROPuytL59B2IXX4Ojge47jDxIgKK
19xfqwrLKzBUcUzIEzTJtXKM6YaSwBN19Ojng+ePN6G4Z7gKOhui7bDPeWqqLYeaVr5fwdbmZR7G
r66jznV3+yPoEFcE6PA3o1iV81clHKqRu39BnulUP2fDsgUUytH/vNFH4ahAFDyMWnc8tjuYZGTu
5y5Xpr7Lb1S5q7rulyhOpJO3xt34EnsBJDfbaidnPC6FVRRBt2T/iUo1yUrthMnsh0FPrj3Vc15G
RGbg4RUDe0DT0kmSNrjU8UYardXSxduu4Bd3Zck20nZr3YTj/8wHiIhWcLuqdbyooGW3gxYbjOho
lO1JbdXDr8incccWP/wGFEuDEaUjesYRDPUKTW+8/YwEtXPmP31ATYLIl32gsRh3wOT2sHzKY02a
gd8oeoUjcqJTeWnE2C5u6XlBOF9XwUvd5RZ2xvhWwTfnkSnaIb9Si6xB8+IshPXVSXKvhoEyHrPO
azFzynhPQ3/b+xFukG5EQJVr4HzhX5S2pPC1rCeq4JJd8Nvwe5n+LrffJUf5ScrWJMZ+nlrjlze7
V8Hpz1+p5CqS1dgxOv6BNxEL885E5qbW5IdAtoPuutRYx1OCGpk/a7KCnSD/2BNujjwl1se7n805
8kxddGWgubvbTCCBeR6+MPuyJXjOW2AhN8DVFuapV9BErs2Bbq+JpKjrp5Uc3Am3Of+zOQ+dF5C6
w64Y+l4DHHRv6pEHxqTmL+SqTC1NOjXE2ZWTjBvgWBHAuUOb8ph24Di24lzKoNcnnx557D4dLeaR
owgJVWr01pqrlTT2ioYT94rRp9MCgS3fAIw7FL8zFDNvAo62lOzLA6Xv8XRe5XL7zMP3bXRr9XGj
sBTU8MH/jKLKCbUEAx1TVwe3Xw6He+hb2YIvCZBch/A3Gw8XOtIa21KZqeLua4pNhO8M1sgSyF5s
E8W0rzVu31u84h7m+Gf76ikwKSl2VATGCho5iLI7SPhKCaygb+A2vHK8Wqx3spV0h/9xMTtRMjW3
bEoAc0k/sUJc4klh+FLUzuEwahiUSbHJOLvFyNjLh1c+249+G6iMIjB7nb1Ha95X9DtyXrL/R+Vo
/8O96wuTcS+NB9Wjnk5zk9+7yBSEpWN/AEq2s1QmoNKHPktWLPygH14C9zCN2ge0iDCvAO26qNdV
jedn2WgeFhogCpDLdQU8Rx7lQBU+aPuH/Infyy78guZy6NAQ6wdibZ9qAfHWbgWTrjFFE0Pongls
8qKMk28/vRs+qKLkFrHHtlPw0DW9XR9KAPQKcyLR4geX0u4/5u39DcfwnJJrlErO5KzH2s0oVPvG
j7K1q+FpBEIkw8TbHHS1H1xm6B/vozCJ/oMWIrYT7vae7N0MlePDNN42Kjt8VQbREgFJuq1FEv8a
9wGKY4iBpgZeOKZUFr0UpxARvyaD4g/KIjaMZVHZ42YwHYBAfbvW55fjy4lmJwaXbP/YVOoxS6sx
T5xjOdrzt2bpPWzcmpuzT32DK7NfPcY3bkM0VMrYtTVR+eRAUWJUJCc51TAURFGT75S2ZOQ2gP3K
mwP6P1vBjzqHtsDk1IGa5sABLqqkyfFbngGDzh8pKie0v9Pe54vuH5sLWBWgWNfU9TWbyoOhg7R4
pY7sbqfxE+PueY65HAyLNZ42pIHDdW87KDBeMvY1KWyqKt/k1G+6Xemby+JaQSzPqYZMXdJv9jkW
vP+/ZL+9T90z2aVQWAeKl9McRbC83XYm6Kq8XJnSIzsEqnYahXrbPIi0XHpthph+XccRP/YtGvNX
FWKpkK6PlKA/ib45jUFx5QdnmFDeOZl5OFTvEeO9i279QlGNqtrQVQhdDdhIORaxbLOHMkQefqIh
xaYajCYjIk7KqL7pT40Syb8NsM2H3I1qZZ//IzWT5dZcX9xA9339P6LjRGj/a7IKzGqfgRv8O+K9
Fo7HHfdnoI6o0Rn9ri/CkzojeTvEAGwNTXBpgFprVcR+qzY2p7ES2hdrffXNRSEUWaU2ZmIRUics
lMMDpooDWH/jWDMiCnrTD7VK/AERUvBqHGtfcBxU3eJpXu22vCoQiQB9jhzrDJ43wVeiIi8WT2uv
LZomxCHfwaTQUa4BJus1fJmAUaRj9Cs3ulYQ9BAQcLTsTEHsI7s9EBFc3e3i87xbtdSYU/h9uOrJ
2TgDjULYFF4gBS46GuZP96BRmiqf5jI1cj+NToag5QpKb2eDlYB0oV6rUfTgoX5n9aH1M07nsClc
L1pMvcjR2Wu1LrZ0L7jDTNWbaJLIBZeZLxkO/sgJInOAOAfMtgC86BJWzh448zCkBHpohSC2RgzW
vrUhZiKhe5dFHWQcPbxOGV928iE/B8rrzv7W/YBBfZ+Hcb8YQFux8cXItv//i7j0qsFlPJfLln7m
eQZe/7EyKqAIUAXFFXsHo0qjrMtVbUL6+bCv6kuEh15XKHLdN0hgzX/511xm3uwc7xBtFMZwOsaU
n81ayFYY+7rqUjYKATb9FeyngB1EEwdCfrr99H95iCjfle/9PF1n+KCoYYILSfgv39FOQo5PPW5Z
vgjZLfVg1zyFhbcmKBhj4/CfEU9CBK6ay/8WHbK0ngFPA05B7fgwBG4IVvGDWTS3yJu7QpUQjwM3
nHywTEaiD57NGNM+5KOH3yD+OoYTqO+O5dxHT8t5AwuJpGNnSkRpDBEVVSQF+nHxyORThNTte362
OoXd/yO2Pn93+0NaHnuQ5iH7WAi0bTC1gglpDpmq/bdIMcqnFlyrifrGLFycSGze2t6F3CQ43m5A
1Qr0udtv1pZDFafmysyRwWPEqg0UAjm/78Cct6z6KBH6fYbdseWpzrbe0+jPMZyqwxIJ2zPdNpzN
HtPgZkiqbEfQolXfPe4NXFSsVUe4VfKoJOZ4B9Lc2q/E3V2RvMbYJ6vvZGYnEitI9UXh5dF+s7If
XTG93rJSGnS+zIMJuTGeyx2OgN5WMxWz3lUyMFLjNtYxQmx9ArfEL9WIX387vvqCyGepeRx+TweL
dpyzbe/W8xuygIbPdY7M7EmnJgVCQF/GA1PXO8GZrbY7BrL62pcwkHTsESdmc1/PjF3FLr4+RjQv
uAeZvF/w8emcXbmaHGc/q9yKq6cE9tg0dDt6Ghvi9O07vyG/orWmb4bnbY3aoqVL8b57IIPAmeFg
KRz1PwjzcFsFVKNA8sPv2yJhoD73nJDI8gCv8wQ9j55/4THPiOJfB62AkDDIEjWL+gs8/nAnb6zR
YyoUelqdGEvE5HAndJtBDRGZ3TRt7NyFtWLsfF0QVHv1QSKyjeTdd6bTE4ww75Ho04hJv/uYQg9A
RZyzSRgfeNYNQB6fwucIK2uTMHHr/h9hiMxoEO4f4KAEOjsUwIPa8D0rPATnuBdj1PxQTp0i1ehk
NX8VeEHyE/j4wTO30Hdwh5lbjUMiT2dRPs5tT2UU3C/ejKUU6YGMBa/4zdgmgx5I02PUCpe5m1A6
y5pUGKjGVixOmgVzS4qjVt22ZscfRAtO9JlGWH8gxFu5XNXHgDUVtxQ7+lmdk/34j3jljDWFEsI9
w5P+CbV8hqJbTbmpkSIJ1t+kQtwmvrC00EhpG7LZj4GqYv0mY5gycHM6DiNk/7ocxMt/myYtPQ8W
DyCHBiGcAYJccuaZmH+z16hv33aqc9o1q0hs9yQFU9jmT0BGrJ961c5i1bJAAddwFLCenq0ILxOw
Fof4PBjOfJhPsT93Sk47vKIzZR+VykWzemtQpGXj1Y9dRkNw6i5tDHo18PdsbRYmfUXrvX7dwQEy
r1ZYRyt44U+aL3v7N2acCFZqKlqAqygJ6xe5HmKxJ+in3xfCpC5zBw7u8yCnXJAmEIX0vnCDuZdM
xbbUr9B8D1uHLoTFtQD5dOA13gqo9MMjr/bpu6K9vqDbSllAhYYtzM2RSmSs5+/DbdMcZ7t8ROt9
9Fvzsvjp/Le3VMAyYIQ4RWZRnsmhVRFW8cdlpvd9dTqmZ0vlK/SukwjM4js8xSg1qpI3BZkBYwAA
N5NrSQQcyumecMJSDorY/cRnJ1XkQQ6SrGEzALQDPS61bKcpmFR8s+c7AZ/EODTTPKyd1TgxFrBx
Oj/IEdfzNIKzoAIpmb8QGeEjRqNKadmY9DMWpecOdsg1GjLqOwWJN0jWoTYw3ZOvwXBq0Od6cBIY
wEPpMDV7733S0SGYt/hN2CBm7RMKqapj16rdEz/Oz3W3rJODHJmAx3jkavjOUy0V9V1IdyLiMKY3
CuNz7OZ4SkB26uDTZOiCwlqNfzznAnqiRLouuda/TMw/E0eL2e+lnO5Meuz8ECg4dTj72oWwqeUH
PPH1Uh37+quxePEZNptoSt+nbW/kYqJWTrN83gmCI86jlpgebHaGXSlYhUjDVTe5GOTQcKpgvgT8
ByRaUDPSPX506nrkz/WFUkJZfSvbGy23UNVHCCivGJR7F6JGGVxoMnBuN6gqVo3VOHtI06x439ES
F57dQ2HBp1LafSmKYYRbt4FzX3DLLncreU6W+5k+bAsg0EAyvu6QQEGog1+hOVqwOQJLM99cK8V2
ezk7GPMEl2VJPCJow3glsm8iRKRlrNCAYVivXCMbhHUHOMB/hgcRtsXtdlkz05nuwuY7bk0eEsmv
mkzMDN96ByGisElpDqZZRIQM+i28V0gplD/jb7fdAeW7BGGV2/bYrlzPUT9D44UW9RBUxgG9JnlT
NBH10ruu+vOUtx1frQloNYBdfFlYFx/45txGOLHiWa8GBGYW+fovKXBBqrV/1QuQpRC8tFq6XzYl
SDjmg2NnCiBG99XM8ld18WqrfVdbx8sBJgZsSKnEDj0pD3N44981vtuZSIOSOTBr4w1H/OvNWnc+
QPDHayNpCo0F06RIMGTWrMhi+uvJnuP9x0kJkXTXfZ0tcItDjXG9MiAzVamjJauYifXswj/ouCi/
RnHO6BiCC/zuqcgTZd1j2khFcvI/K2wN5winh5fXJcfgyy4UW3927T1LXA7hvM4RY0uf34PlRHm+
LY5rwdQMTXnG+hKXI9aZCoXbbiA1dqA7FmlTLLVktrWxfLm275IrHL3YAHsBTuH/zDAU8z/swLa/
awVrv3OQt//IScIxkc0QjGFI9WJdC/F7eEJxlb9JImzFHW4InvlqrmAAcAh0MRJHuBPvUwhBkgDi
1G8atrNr1WVSEzcymZja8oJHvZ6u0pTpGhvF6B4prHwgVwab33J/so6Rsn1uqjc5mS1nFa3ap/Bc
YXEJE3CX+rkVlGfzZSTnSPEmVm6+Zb9FBskPvXmaikGbIAy6ISA2qQxa+wccj47iY62tpafJN/Cs
4aVS1/IZZ8+BGz1M27r85SwAYZ3MmutdT3eQ4EJNd0u7lfj2fDZPH/QkKwTvB5QT8wVRxuyf5Veg
CegrOwCzXMHkXBckTYvta2w4Z+foLs5TI2u0/CPUogVYv081lzC139KFq2uZRRw9/71WrMB8v4Lj
PfVAuiMVaxqJwLf1X8GWsMcEcWsgpvIyjdJl94H7a88ZzyrC51Akwlz3alap61FZkWhSd1J9/OCN
3QG7bMzionMATkLAGwq0GeWht28ks6LuBcDjzsw+zdJuK/UjcOtPBWGtyle1gaRaXlh80KtfeCn/
WR1+HWgtIURNAtgl2SBfPt1h9QhB6mPa+VJr0YHTGVWXDFW0VYkh9mvvMOPbpbj0oE0HDj1LjscG
8FOrt3ZXfZSeouT6wimtgj2YAEbA8aQZ8IZLJkHSL3d2KPia3MA/Ao3I16uplhNS5UOgtb3SuWFC
0xTG5jwnO9fTt/UbyEFFztFbBgcmlquEgbxHl9gxSngRle55NLv939+fSEbDvnuOvf95SPvGJunR
gLA94r2xtndXPJC1QDjNkj6EuuOfVMixiZCb1cwLbG4xifY5H++dnjnZRLFQwI0VoV8FAgC9kr+d
RLDvz5hXnkDOSByN145TT9q6qDvUKxRQT6s+zuHDDPMF6hleBn97/yUi/4OAeFGLbyW22Mzep51W
fh45yXntC0t1FueR0lcg+cRCrw64ZFhr0Yb7fkiDxor5xTdPKXQbg7pC1VogftrDJjsD/Qm7Tx4O
IVq3Yiq0SjgZhBQrrgwIUw/WtQoW+Wj5EZGhZ9LPtItj2z6zvIqLmF2Lwp6SOPsS0u0qnIeetHC/
gDwWQXzoxR8Q0P1aLOa4PZs2XjYVPnVvKqZ/GS61T5NRVBsEFsvUXdtizI9nethl5iNDT0P2USmg
cjPBN+wl8QYi6RSOT7Pbfri2VjOtYDZNh0mvgKSTSGXXkFjGrT666RGB5BoxADWQYekwgtL6J11t
zD/cFay3qVfYL4CWW6LD8sFG8tCDyjZriHptGt7a+xxlHfTgGa9Rv+9MN9mUvU9J2QC+nqfe+jwN
WNEuhZ5+qE1Q4Au02Nc04/ei7st0OraE6j1vXyFvQQHkfLQQ8Izq3mOEuTv4cKmzxilEAFqFe2W2
YtiJceGDYQ2rH7+c3Q7yizSi5l3F0COkaAIFOEvFDnhuTsvcXl/0gd18JAZOxR9XiXNC69prE8AD
I2G0MGPS1v1pUL3WcVHSxA5jQNO7jJj6PKOAs3N/o/KR2MtJj54Xz7F2PRFypJfHeqJ93S5V51UO
h/xp4G2v5CnxzBwakLvuTq3JOSPNNR/qLWqUct/8DYwiSsNUnk9Lyu54/HDFGV+5avYFAoSJ9jML
weXB7qA5bXpxXMqDQX1Zw0ZpoFzabIcoSnDr6lPy4YgAuoc/2C6P2GODruia+tPX07ssBNmhM5ZJ
Fu1y/+mEisYoNj0HFPoEhhnJHnmbZxrXI1jQ42Y6XYbdGjnpgX/5UV2ee2kWync8W2ORDaDTf93+
Qf0gF/jkb4Hip1+NHB7iRF/GZJiwxZ8C6d/CdY+ntMHCpSdOihcT4DuftYPcikGm9Lfs4ECJc/nn
KowTQLBetY3kBsMmPWoO9YWQFM6Cy16TggMwnLEj/8sbvHdyADQXEwa4GjKmifruI2uyhRn78qaL
KSEWT1n7f8gDmpp56PFUeIQCs9jfl7lm36WYrDpIUlfpGVsnCcyPRemKwLJJBKQ1WAU0+1EUl0e+
Nmy3ojmeIz09u8JEPBNn8QnUxAnoqzGs0GHsGBh0XKhNTnlSo/Svvk1Rr5aPFnckBaByb6hQjuI3
A8VxzMotvr+DTo5gwpg1HcP7MywORSSlDi0DpurPpDAdFqGzq8BI0uHY469yxquZUS5kP+3w+rO0
Q4vSP5I9GowDAAQ4+Ps0cnt0VYC0LTdFwSVIOxg/8GMZmboMFemmtNHbpJe8ytXFpdY4/Gagh+t3
yL3zkvpy/X8PajfO53CwG5dURRhC6Jtv0rZlXec/hqiXVAKQ8jtXzgiGU6+T6R+IPG21tDKMEhgP
fi0emhAIgTvyLpF8Es2igI7n1rGOkUWNAn5v2VR6J9qvJ8fRKT2EssZzHsEi1nCWr0YDn61mTKsb
iWaQGgXrtuiYVSaGV+y8ZbeLlIgdSkRfIlQdPwqvw8Bt26hI9RhFV9ExROeKiyETQp6EqGwshapi
gm9VnD+4nxSyskfY3IgjpK/LQ1GlF6X0O5S16fABqLKBayBpCRWEzdbdcGKag/MMENVgmFcQ0Qsy
B17a+0ew9MoDaVEvWnalobJMoKiOMoKqMYFAwicOdq6vGeSimQDfJ6Rnk1tIZQ2Xl2BVAFn20rcH
/PaVsh3rDg/vUpaAA4ILcEs8GzPcJ7RkUfIJaDLWKiLg8PLxJNzuB77H/XYGzpmC8CLIZ45eJkqb
XQUvpoinRBw0z4AkqC0lymQ76aSsev2hgKLpn/k1y+K7F1e4LTufQmHKpYotxPVeT7x4TVLE3F9t
dUDchiE0bHW9XiyNi7GjQz9pl65agr7vG7bMF/WEvxmq+xqa2l3tBGlEebwsx2O33a4ib4c+qZAt
f4qmY6MPjKFhjVWN/9QQSApDPl2WsRqdJ/E0jWZp7Q4TckjoJAePwm/taJLVi1IQYqikdysfS6zH
6ySgPRS7CVS5fE8El+FTYmJnOLTJq9K6JoCFGPCrrojNTph+xyZMC3MYL6zuclv5KcR1QhmqAeDL
nZF34C4KUYi74bHKGKgkrYY/gTaRJe0OBv/EVbgsjbDzx4GgDTTnBo1baAcEqTzhNj//wwc2/AQs
uy6L/XdkwXsYBvg+x1pFkUd4YOmMCOyUfebhdrBmjRdIpTrN7DJjbqDqTdDacemMdDsNePmDAjI2
AOdl+zhNrljmmqFjsBV2/GQVHbv7IgQQoITRlbAIaPEFyW/pYPy6MQ1RWOs9K83c1fqN7Za1AXik
Hsq2Qkt8XjWa6UgbuCt7QVak9dE0Zku03tNLeuLIM4aeXcXdXYFtksyikyEaKLwUlY6rt8aQJ9d+
8QKPY5grKtw/mNUXSV9v/V7zUX46SGATE6JT7xCcDeIRpyiwTTR5UsI+Di+j0OjSDj+SsMZTDgBG
K8gdDZJSmC/P6h0rymbnALpmYxMGsJjliAuzVvreO5pwpPr+jltFb8+rN3c3UuDNV7oPMPTdZECw
uoKkiGMqJpH8fARahGNTcOSM4r6Zwx9J1bpnfrBysKIUilfWYxl0sv9QkxynYunmE/UrpcJhvCvB
4m2oi4YYXF2YPPRgPhYkk6mYMgAlJKv7XAun/D6PlEyPI6/nS9SbOxsjYnnr3Rfs/U0jFWlXRZMF
t7aqWcE5EAjwKGLstxoDAKHICmEWzYyuio0TZECrJfveymAzLGWHUDSLGH4niIxfZxxlEzBQb6wO
rHkPAlGH5VRnQB+7GG4OB0OXHKeW7J1oS5NT6vk3YJhaQwBObmzgszUjW/nKBSv0r+CA5XWC+lGD
7PsYYM2HsfTjNI7lQqfqnNEPmjOR4OAQwupwWMrTiEyTQSxDmTGoP2ldVvPoRiwO22IbnTRdKC+n
qWF8ftsMA7e31Fij+6Em0LkpruSLYgQ3gMiwrLynmazoymPny34bSy40S0q7cSLE9+1cPcn7bXxa
FbO3pPt9CZWiFIz8UvSP6NObt4QbF8TQORReBH3HJfl8BsTIaR5Jb9+79rlvMnBkdrPqir2SUPfE
Ulh8nkWtnhpdVA1L28E/hdq+ybXoKUZb5rPZQY3LCxgZddN1geteXx/+n7wEHvDSSEOrlSU7NUjw
M4D366ZJGgCaBDcvO+bb5NLNlxL6puDOx8JYdg+E9jlhnaVoNFIXcAT5tfjjb85I4TlJt4yV0qNb
IJFOZM9+wEGkeUM+hCp+8R1kvjVh5QsSNsp50EwMc+J9ye+/qI5RCM4lQTWr28mV9WqroNz/0/H8
0kWChZYyB2fGS1gvfKFsW307JCACKmgVSwlpdw6c6a+88fA61LTV0yy9R//aRhheqZy+qTB2Ha0x
HASWsBTBdfM1BrQlDZ3lfMVQIOhOTa2OH7JaQ3UVF3llXHplAn5fMh43fXTWlMUXWct+VV14EleK
k/XXlzSa0GZiJCpVlG0nQc0ByTjNrHVNsFF7Q9W+zP2QeV1/ppN3uKzPZVO9CoSbWhhH2/5l7b+I
ygGl7n3guw7yIQqKkTchtWjmF1OOyhBWOQ7/P8VupewPRnIZVDFbImGNWdp3WzzDPo20HcTSIpZq
iQtblS/o8xUFUFtLiI0F5MG6Xs/+ZgzQoDICJb9RbhybtF96cT9z6dqxp1PYG58j5m/CNhYzfIfo
6LnN0dnPf9StLaJYGmp12idyiy3PQp1EGhU25TbazMPQdaqCQ3OPgG6h00GkstHVtE3ny9qfQS22
Qom7fUJzrOIuIiqEAXfGmGEDPoR8NZgPbbYkuf5X3nh+ghlRt0bfWBNmmZYdB0FSr4p7muHeAL7r
jNroCCZLpKbPgV+WthXVPTnbCDkzmmyDu7xCWEsyt9IiAvvdTDJ9KKBuZ2cWMIoJ5Mn35raDoT0R
VoIBTycMOg02CXINCOq01yGR2MiPdIjYLkMNBXr/Kjur90LkqlM0qlkm1siBX0U1GWyCV/Ru2ZgG
uI+EPzh6jHC/tu4dkUj3FqsWMl6DZ2dWYLuiWeiVj+PZUy7D7U879Q53TvZkz/73CWzYMWXZ3UY+
vBu/gdQfoEkZ56e+OlOg2WYq8Hp9LKFFKYb4k1PAlomsDtcOyQg2Q/AzomPIqKr/tHcuSFavCKt0
dPT9zu6Qf7mrH8YUrqHM0OKBNmsU2ojXsd3hs/l2p/1WvwQveDaFtVMxRjojGHfIT3XHyJMyRqjY
I2OosRATqyRp3OCwANokew7qBHsreri+FAGfyEihYBoVkXXNORXAO4ck/cmuHOp4wsJzqrc7WrDl
MFWXflBnSuICMGSPWLk/7L8c0117Fa+5u7Qwln99VB9HzZGAIScdXdHmr0ttsb1nG4Wv7rwpm+ki
r1UjWUZ2VWi3vzZwGe3P00Rbftaaej9EotPJs78cse3O5wAPrmPtWiv/Mb5jhL47KJmQPoHzKXkK
c0oYHq8UEaXNYGR7cAdgHjTDkFVGrmN4asIoPISeQ/Xg5NysWqfOs9rh7P4dp4GATzJL3s0afgm6
+IOqK7Q5Wkkj1kvTXTmjwzmrdgEBvjfdP8EIgMTuD/bOxzkidEZctyU9nfLAFMirv6XPUGGzRMD4
dbmNa/yVxEPlSlZAZ19lSCVyYmQkTHH9HENmDfxpsuFKCl4bfwL1cnbC7KYo+4oxMe3hm/BmODmV
rAWmlKa8rhgfOGY60d37gBoleIURfTKQg4A+5ODULLH9qJXZPsDXysSvxIPwp7MRSbz1x1m2hW39
S9ikhxy4rcBwU7DwRh+LRWdMS/pLvhz9PxueHl2jnWKqTK/gMEkXCEep8ADwPON7xWhYFZFP+RcM
5l7Cxk7SnIv+/4HCan+Pqb+80KjdgBeC7mcAMTwQ8GISZzdf9yOLDxLyihUZ44IL78TGGrUN3kxp
DOj8btjW62fliFDyFJxatAgWtn0mxRz8jjTuNz1yzHCfftszzcroTaDdE5wZFwiFdH8mXVxhwB0A
fAFunqKP8opsMMVtl6IpSkja8/nc56QPIXDfKrV9mw8/fVyVubfic4pyT4woXdXHXi59Ybfo3nyw
3ZhVlAc/cwslQjL8rAwL36DEHg0Ew/WKs2cWz1dVXpEDRJLdLAfzg63kWR3eV8LDZ5NlJy6uJIQj
UtVVzxDYsmJ8cfVLAuLX6vIVnHClBNZSSXMZe7QV2lGoBQLEkPYyJMwHo7d7Zv1azl1RQ4QcDR7Z
ZGB6TISKwz4vwsaGmcuxPKhZRBVzLoVnqWs8ndXLJ4fRl5qPasDdIqJ2QuDRVTikD4lnIlW5c3nT
yo1gsTZ8NAjQXLAvG/Uxz9te+AVXqb613XyQ6NnVeqrrLLV3GjFDU30FHACclGGad1k+iffjq8Vj
1fRJNEXQZESOcUprYsEZ5KXR9W7E7XDICkr0J+FdAt5PquzBhyeS9kfDJM7kh8k4tD6ojf/Yrd2P
byqkGWxQPZHjkbuaIYWxMfbnjGRHf83KzdsoQcfEUSIk5D97DTfVlRwVWA5SuiVs91TDam2t70cJ
ubzyLNx3iifPvxniFtgjyq0moMfjhJMPSnoshdImoJkhsgyAOK/qopD62NQ+yjadmcwFrbWHHsSx
qKQY86nfnAu6VEPz3b5FJrtgqs6oVu5urZxVJPxWsr9Ij/SPW4cxY3CqViaAg/CRd6bNn0bSfmxB
kKQfgSaSgP1N1qimS4TZQaSF94w1lh/KaY6osgTdpBqPhqvOjQ6IxckQAdWZeflxXKMwig34QU/E
ENwqXOmsckngh2VsJyG/Bld39IRND39cRy6P+OHOybLziPQ116hwPzEfniUQXiBYgZIEmKXMxamh
RD/a47Z1bqznm4ursiJe6IS9HCD3XD6fFOSqocZt4EM0sVGfazRnAMKPBmHyiaeBztuIp4dJQiOS
EMadrDgbAw40A4qDXzOMG9njzm1Y1C7v9UNf+g8jUvENYRth8Ar0yjPUByb87XXTXrrJjhcxhp8p
B72uoXOh66Pb506pilVfHMS/+7jR0mUtMHv08KO0qtLx1X3mo+MDD8jwv5xjY10on3dwTgVRTo5x
gppbGefk7yXBlOBpBTbPBVlGDx0VGi4ZLhSRnCeGgLgZIcy/iOW6g7gl7Kf/KT3MuGQ06cPsx+Tr
xD3Y8HnGW7PuK+bLROGFm+SqvhWg5VYptm6X8O10rkINxehi8CvosqzYQ9Quuw3w7Q6VGt1dkMsg
oe+Eaa3hw94jKQtEeMXoTiUBbqL2kUSEI10pXLMZ+HqhpggCQqSN6wrVIZHBH7+rfpiAruHXj+1h
CAdvrag5/ChxtXBanTTGoEKtPsVp0f26Hif/Q7eMVA1kg2PuYhbZcsEtqYX939x0NfvjcMnFoS/0
ADK8hXXfi6Q2EAye/nKJkjcvX0PNN1wC9B3+vv9zFJI8HakYo5Q/F6XVjRyHyD3C5MMpT8t+I4Ir
7ZCnlKAlWSIwptFZufaA01tD5o6GpRS/Cn9tvz6wvkjKdgh1qZI/k66cUnK0QxhurygHA5Vc7MrD
RoqKTsLaccEWucYVGk1ugnOM2Tmy01vDd8wTzGGIUnPxd5OO8zwsQFmn9UNOa1wb6Ay9/lJYciu/
E3rxY9hpPbNIL996JQBJ5X+VrtnSKCc8inU1ynAct23EhRfrqwedG8CoqdSZefoRRV7F4qoxbjrj
gDz/3D8FvT6ILATM2Orc8ivJrQS+HX2ONOFPsLWav2FAwp8VP9m3pIQq3aOx9DhKbA5cljqObVUn
mGo5+iiDU+Cg8hjtTQZUeW+p86Pqlpq08f8xZ9QuL8b7gun4Tnf60p7edz0CqpCtFRhCBTrq7dFi
YRd6DQkSoUoVDKJ2P59ubekw2HDt3An7JcnS0K2LbcBGSs39ikCReEYxx14BwLPwiZr6mSo6XyDy
6IQAvMgmnchjg7oEGoIK3hF6yl2kAm2FFeDkrTsTc3UIRjzXuHz3uu68948pcZi5wytqHTg9afI8
wLqrlTVKVLTDscjCvV5EbMPrCU8cRrzLYWWRmjAoxDmOFDXEsns5QnOH5KP04YSxfRfkwi/pl0dp
LHyIIQXo72wS63WgnhPfP9NGYB1MR5wcIdqqNJUuWmrJf7FMQyfe4U4WP5Rq+KDNpxbX7i/y4Deq
VZMZHyexHN0WaVGHsHU7sH5IaN8lE0QIDHOT+7Nd979P81rVBkVWLQwXQe0odkuk33C8pOcoN1vt
dr2hzGD8uxxhnCmRHXM/bRdQdGOv1a4mD/cEml8vxz3QFxE275LxoK5qz3xE2OV2sRi4WedZM45K
X6E/AJA0b0H2B28lduGu0aBT46P0mRYe/ZKKkxSVYHzsUsl5HZsO3hyI1LDAaS/akLcUcY/dOkja
s04S3+fPq4LDzp1tPapyYP6pY4/sLPtgwl34zHcRx0d1D5D4vyEPsJXCFGa3+bm1e3a2EDAx1I/q
ikv0Lbs8/FPWOtaOqkpKpkHpYp7uCL/c5WIfjbas2/DqjxJZgfRtgMtiPnHClAzZglTmvca8849J
eBV6R8RrlHff7ZP528NZk0cFjzsVhgkXGcDJZUeDX25TUdWJx9Lh3zJHfL9AqZ/A79hNk0MnEazA
Q92B+lax/KWV4/IRGEaJOGdRejtL6eQxNJtHpHbOQ8TPe1MxF1+1zWPiXARQ76d5LDxZ3I1a3MwK
DaXLDjUiRBWljx8xhWuz2OZq24315bjqttwVK3uzm1GomqvBLtQ3IAryB/QaJmZWX7mmES2IfkVn
OwFenL7mEnXC4dpAtuh7qhABgUa1ZJpCxRYNvqp7CrUuXaFcWDJkNiqzNlvVEaL1CVH1IwTN34R0
xy6zd59aKlzDBebkzTvp9/uoSC2BAT5WW1bjFlHY/sCbkP5odxOg/ExkXvuiv5XJ8JvxcK972yZS
OMpTGwqOQlC9JLeJ/5bz44//jcPB6ifOUZMxidtYvncxNqIGTR6daJWY4e/NZlipeVYGX2Zd5l8K
yO3SdaN9m6ISlJ13e5DYaMgbXe3v92qbe8feRG3bQNwuVp74fWcJ2eYCx/XZIEIgdoT7nv9MdHjO
E1DKIByI5Y95f8/XmUzyQJtNwP3OEBp+l/f5ZlRH3zJvZa5J63odDbeLobPCe8TdndLTPvBBkvRS
RC1HHsnzzjzazyJx7uaF2l8khQ1TWXm2DLjFReEuAOOWdXiN/RuvhxkEYLWiQgC5rMc6PfC628E7
1xgpx0ymBlA+61fa0kK0KNTQSXCBX71n8YaqJx9iPkmyGEtsCWa0Clqx4quELo7qH3lW/n83G9qo
jgQadyyK0g1r7CSaa2v/CD8BySe3CsVaCgdGjtyZLSMBv6OE11mApZe2qy2NU56CwCDgc9Y6tyq3
/ZlGoedwL+tA8CmPgHBr1Yvvkawo3m6DXcD07P7aOKDVs2042ILJy5Vni7jiDgG1Il0FbzVTPWvQ
gGu3+Qj2Bn9MkIeJhNRn9dRbeez3YG/ri063UPfXVohb7bJekrUXaDqfKWGT1jimVM7iLTlIE0Zr
KcvzyM3AFQ0ETbY4iHHxGy/FQ7SjRxKrMKBMCrt8CVzFNInt8j3qRTmZbbqJcrAbJxgSjQZYXxdX
rx+pP+Nq4opVidpyoa9UxVMtotXVDck2jqtwAa4RkThbSmH6c++fpU5vGGXdD3oC3CobcxwbBEo8
afm8k6+YTAmh7JrbjrbwPgmBtEB3X6QQQOI41Jh8/ebQBnzIugYJgu8ppjNgh/SUQLq/xPbWC2LT
YyYdZi05ByhyAsDwc6tq70PULELig6xMk1B8aUqZLLrLU08zmBfR6nvGlmvnSaAzVDHt8cg0r3ze
tMSqA6LMUq1Km5dgeUkciGkJgJeH7Xym5CoP5RiQWxpViPL1JPlmEExHcoow/JChCCUya/LVEGfm
s3EISNhM8eibF6Mh4fuvqsksPxBh+tU1kPvhg0xIdg9QmRdaOcAN6XrJ7nbIT6/8SS1w/xIlz5Ev
dqNXKSGQqEaL+7Hagw3Pjcrb6Pw5liyfpF4u8TMqBbgdrxPSF6cf0jSLn67rps0DdZVoR68frKJ3
8TJwhBSlH3g/WT5HGubbL0WLG8NvXoY3M/LHOGp9zkNVMtbDuRAxLtJ0GU1OWt9QHInL+YNY/nQv
Z0v0pYvr7isjyl9JvM36Ac+0BC7Xn7Yk2dORpeL7e0+HyCiQ5McCz16Ip8eRKsoKhaoIyNxrbBi1
FkB6hsANQ7lopVlBJ7NS7v0zWeRsKiYwnck0c6vlT3BnIU/Gnoz98NY6nwsBXemZIA/0RSV8AGjn
ikYgAO/NGVwsla8usUlBFXBMjtoqNOb601rSvR1/1tc1jGqpl7oA0Q5vkpC7+PCJY6Se5Rvx0bNz
6ay8L45NcIYeKBadHxCzWipc3Epk+F51oHVfNhrwHDiGvng/0KBGV8u1WioJG4rZZG1sFQ5FbXn8
CjsY3qTnqxJ8vFmcKorjATXdsZ0xneVK879lwHwRlHBc7YY3h+RV4s2CsvJiqaIjQlo0bPRU0pMR
TMWdCousDckkoaRlTD9KD7ypG0flxRxSuGzV12Okhfm63byFTvDM4RBIuiQ6wKORx2oH9V5AuaJx
sb0R7AF9cUlYQvdFuEydzHDaSlgpjwOV9KidoZ1795mQJjEzlcX8ZPqXq9dF1zNKLRa2bPvJWRnT
tVt0ZWhR9fVL41mEUqCQ762W1knofwnSq/VP+V6MYeGTnNKbXqfJWgfzLBZ357UUUp6+QPVFmTX7
Ezw4oTfcEwUlZ/Hzf8qxzoiPNSNBR17U9oHMooW15EKzhhwvJEhJjwiTz1DAgLSkR3wvwUSgKBd5
ZyrZDyL2Cp2KPWWryP7wbOcQazZzRGeZvQ4Ls1rJ/dw/4jfs9Is5aRIoMGBKVTuSrwFlYn61fQNv
PN0XPbxJLkBHZpLHBqPfwi/tl6ZasL7zHmK9aCmxMbDwS8migRBz2zJXGkayoXFlBz/9wRiZXSET
CA1g/6jXhoglwU60PEDVofGI/4+1FiQqsgFRQBusaYjkiDRVOiHeDZG4AbMy9s5pyklYAE8yFUov
Vroxxz0swodzhNKrC8831X9q1Za1/8qpX9luNrSvOezK82/7wIF7GGnbTEj/lxbIgIaZGMhEYZhc
dHoRTnnlLD6JAB7vXkWgsJcX7HVo8nIy08pRT/ZV+wg569VxptBL90SWeND5dNfZU1+26u/jn1j1
Hg55KKEHq4n9E7NIyS157fFjUQCGkm8eXqEiWI0Ou0kpDf+948TnAvZVa/xh56BK5Ww34BkXy8k/
k91UMxsMAFM9r0zU22sFeCL2y/IkRxYTYZ3Copdf4aO1v6p1Cf+kvrHS1NbLF7Q6jLTFCGlL40jT
6TdGieq8uBQeBszIuL9vBdHRvjHEFVkJT3HbSwHy1SI0wOfaN71jF629HzngMJ24ljtNjdd+YtWE
tG3SbjKzh8VArX8iHP1pLjK36/jQFeYU6TEvFGPARN4YszNuAcdl3QcwnrgucZ3bSuFQbpg2xAhl
MKxF56JJqI344p6k37oIv4kvhLcabGG4bmIilxasUUI1+q8Vktgi+6c6tE4PTO/LuNcDG0cxiY/w
/2XHw42N2NbM8DhF+j+z7FMMTYUqL6qRJBf1z23lDETnuh/QJVWaJw5Av9N/iBSdtKs/DGzXIU1M
cuVVow6qTcTWJWJl3msoRwNYensXJ6Bq+CDrwU9l0q0VLb/5MjXa7w0TZJIl4+mPsJoUEQ0vDZxb
qE76Zwg+TuPeCNLo9sBG1eIf33d8oHNUSBCXK67v+ukDjAxXaxgx9jVxY4ecZprYLwjPLCXvmKGf
ybKdcfy/LxaiYlQF09uUvR2ZLmldIOYYw70zsVUZLoDewZnLFZa/fQ/X3h3JAo5Jd2gP9pt7VIrZ
n3f/9lGVtH00QEszkVT9ENgGQkNBh+0EUGxK/fyPTKsGXSFdSBRrZX2Ej3Hz5b+8TeZ+37IjjaZX
/izRzb681E3vSD0DxnHdh0o/QCviiGVgPj5J9YraZ5umj560HFH7VmwbP65Y69ZRL6WQJtcTct1X
Phrv8eWNkiRIehGg9wuU/ZI7MbNu4VnQfpT7QQw1ue+43jg95MYZY8JEShNBNK+V0PUGLluoP4DT
vXWuqWFZs02VUuJBNyKKDRHA4mOvQHh3tVHdPJa+ir/4loM9DI5GXZ28fVPrnREtyDol0AhR0xIm
UYlwo3rxfvTNXxJJ5n+f0NiSS5JHebhOVT5GED5ntwNiItU/1F8LFGhqoMpYEwVFhnr5zGVuqOWs
KysKgb/QVbSt3Wx4oCOr6SWZUh/0AVmLNbvlMiV0mQANQdADcgOM1FnRonN2SgQGBNUIXKAfSFWr
BdmnoSg/seDCeLflT1lxSv6MtO7/70pfAIqFKlQZCVLlPpMd4p+kLAa1MHWqAbrOebq4Q/wpPZMp
YeOVDNct/bcGwgNBCIrfR3toQocJJZ03Z/ZnyqDeAUAsZ2AoBOp1Bamtr45XCaHGLhUdRSxjTvy5
XS4EmfDyZR7+gEHFAbWivA75ftBOoa8DMfaIJ4ArE9UpqnFnrVXlgwSnCJMCaNLoOIZLHx4Soztf
LzcKdqnEZFxteqW1N3nkTfu/ayrozqCzo2rVlpaOAg7v7zDGu0wqiWB23yaxA3xZiDhMqU2ZaqSX
MdmTEbqqM4tssXT5F+ibz2zFyPyHBv/JDkOFYp1r8niJd6feFSas3GVMy/IKI2FI6Sun/m5yNkBL
W0HHBBMG0wBfwa8pTCe5ItOPZ9+O+vkA9V9CiLPWrlnk6nL2dwSyYD3pM9/j7nf3BzxMR5hAnL+X
Y9RIKiZKnHvOP3ZpkOlhC9xmFwXkkDaa6YPIShq0dbtvU2QTiPkCIv7fjWOGWZA6CTyuOhLtlrEf
CWCRI35V2KemmRi2AwyFs3ztFTVz7k66Hb0Hl9SCzZj2t/08zK9RTJTQHYbgXjO6fLWknq/IOil+
7F62nMvoB2W7l0udN/1T2U2LrERoNgCZ1/tA3KwR/3ZR5/2cwiqGanGetZTvcvsfhMs9YbAlWpim
Dh1sDW4Mj7X0Nj2IgcPAbbIt72RlSQaMpt86NYXgJZrMRuK3zRXlC5fGOF+wMPrlVfB9nEfRKi/m
QIpROcd3nLFGyCFinuCszADDAIGQPt8D5t7hVcmkIRLRyM8XlSoZrNMic6GLkgiKBX55SHKznhm3
YbJY+024dOgx0Sm+LkVyXdRXIb7+wDnoHWRKhZD4NGul4vzlPYBJNR1KABvmyxuS9RGc+8/XAOKj
OatpIByAf64iWBhTCFjVb6UAPIJDjM+v758QH/qv48Tn4w7Ouy38PZAX0cwuSOB3lVp2te+w63ME
k4WgDhXZVuJGB92jXzVPz089yPRpakrRSQ/+2YTXYY3lSD3IhkGN/a0MgMD3wfyiplr24aL74VoK
UVu0we/sPDue6wnBr2LKaZBLVvMICFauwpgQSXKwewvqn3Kiv9/J2aP3rc57GWNyyCtiuNZZ3LcL
xfz2CEVJi0QRXkuV5cJrqZ7asbaTQKhSKEaDC1vqWlo8FVXD0ZJRnWiXLAEycySFW37lKmKHnfpn
87DY3vDejexQ9/bsW1f5MKeDZJHMNb9hg2KKX/4bp/Z2PIQR3on0ivZCxMC60Zf3N4ixIU46sPmF
qtVYymzSZ/2MM0DNzh41p04JoPhRY364kZV83N8lHBoT3s5O/0OTcGQQ9YdMAKi0cQh3fbp1HCi8
xkLDmekG2ep+4Ss618EkfmMi9+5wr3kcDhgUPuXdlTzPYXQvp+/m0injRgC5AzjqTbtk8AX8Ubv2
EWNN0NznyjrVWCJRSvgtOoPFzncgYbAu+MDa3PPrg8zu48KgnwT4Pm4K966fZ9hbtZQ/YN1rX1Ul
IgCGx7YHRQLO1zTsEz+t4/2BDsAcb4/0cserNkHkdSTXHDUlAaAsE75yAPONh3VwFlDoneZCM5pl
5n0Ruzm2hcQP0TSUEQ2eM2ZWyf7S/H/ctSIns0bfiRhKam4dxo7Nt6fKQ+VE9hdi9uOyCmjL90Dx
VCZV5b/ikObvOIUk4gS7M34lkszshWccY0EAo2xNaKg6K1cJcQMgWti/wBHKFQ2QctOydVBuVRv3
n0RiCgzqBavFF80UHZR19Yls1Af48mKF4LUKR192yBmE65UpYRklh21fkBIHFSK4rm6o8zcEHoLW
tDGlbNlMmaT9RjjrKEuqWin8EkI+oBPo01MMVkI5pobpmQaEmM3U+5iCc/6RRscilli9vENQ5Scj
DR5RbbsHtokN4xLoJ8jc+f2RfSsoexvwrWZnOFB/lFxxgazGm5s5OFaIW/yZhAqA4Cq0sq4m0jMc
CJXZ0al1+kzmWyWlSiVxdHdb9eqHFRaswZS24zkt9hHAIn1+G9ujwUDVD02PDBVToU8hrhJDEktr
I9eO2lgZQ5RMfQH6ZvpdjylmBnqJfIVeO9/HiS+Ch5c7X8bWHpENq0ezT7MDVSq+lnIF4ga4U87b
jyeigFqrvFAKzkgTABdvPT3GftbLjJsxZZFVNZJBZkHmTsr0H98HiZigKUydrKfnBACtVVrV7qeN
1snzoxaIKYgZUHQ+6srdMU9YDHP+v5S7RKdcQO5gB4AGM0WDKNZmusj7G+YNaB/fvyWMbLJk5BmE
/RLM4UNv7wfjix3W30/ZtpEuLNTRJ1rexzswNcrQrxqDF1l4xaQV7+kdJ8vdVuJRWat/fpGJaXqj
eJZjAj1nsovwFxJodfZR3//IS6Hys/Wot1iqSunsbO2Kn7BbEnH1XLd1EaVl9umisnCMmYVO8O+j
pdtSmjvxwdjgchAE2d0Qyhqh0AkW/dKzc7LomsitkjsSrsr/SlCGjlsZIyf49R1GuJodWFLZYige
iDKOG7V1vETCuKygf2m+wf5zyhp8NnCm0XKJaXdPI4lOOra5yOX2d6ED37GrkhCqXAHP2j5yH2bt
xPvZJmYY+a4djgYE6GHiQGGmqBDvxOfA2itwxUb5OBIfdHoK1BEN8a0GXn2uqdFOzA3Camrhiu69
53OIxE4jFvxFFfwxe+gQQqZt+tvfNKMrUf4VghQEkzPGNpyIO9glAjoR7/nLg/QCDl2qf54mYZoK
bR8xgAzNY1SE8n4T8VBQK+QhBl79rgp2FSJmTJwjtmjoHuDn/5eGjKxK1vos2zYWzze2MgbxCWS4
QFQXmdV8kLAyOpa2a9RokijF/HN/8hgzLK7cxJaWfTD8Spk35m/Ca2rUPg5KsIaspUw6dEMIsk6Q
LNnIvy96xK/wC/wWueSoev6fA9CaYsJlVAZQ8tywWLneFvFxRh1RacI91YwSbGT2WxwgX9bRToZ+
Fj7lDu/g4np++xHliWvsWLU/NSSWs8sr2vaElZa133CZDKBd+6ZAkhlwFvUJ1Hojo7Rh3dx+EdCa
TUJrDsJ2qVvVOw6Q7T3pGa29uuJcX/98sMFNt79rFfk8imYoy/yjBpaGJHqQUa8nSeYkY65a8KP5
z5fqwnmULmmzN5xQYWBW7tuOjCsvUoeEfilYH8DUhfCk1Ppi5JCFfDzLZvxSXJs9CpWAWYpUWQv+
CtBbO38Mf10Zm1odinofCoB2ERGH0wgOFL74JNjHi82PVY53eYzCXx6PnjNYH1nFu5142raztGBL
kLZ7ZTZ7i1kP/aNfGkKuZfSjt+FmHRYo1f2xioORHpo23OVGYmKEJKpPWS5koGnuCORcP6H9mtoC
tcB9GZKkAMTGA5BCTFs4alilbX5/64lG2dii3FRBrBz7Ku5l8i+FYnKbWtFSt7QnuBF6/9dsiqsk
TsZjaBnI1hKGZ1GNTgmF7THxIHU8ccAI9U5Yhia/chkCgRfQeeq2lZtu5CI9vDcbd5s32QjxeU55
ML5opIvI0JyrnH/lq5ZSs/71S63ZQg1L+U83NsiBl0w+0B7hnedmznk8wQNJdB7WRE/dbVQ6+jUr
mfD93sQz7Qo+UUzsG6qru0WO5FedzYP44JvdhNfKFXEu4aM9QJx523h+yF46i2L069PcPmukabqW
norseFe4SiL42k4hHzVU3t98pNbxuDBWzSXuaM47TQ/4uaspSV3gZuFUOBcX43aDbF1BVbjuGLKY
IctZmeChYtB1Mq38b7HgEybNyo8+xypgDs2UpqvqzRp6ddLUuuuDRNKFy4z7CnDD0OWiKLiy2rUW
Of71OzAhlwumz/oZUFvCJmyN2iScD2LPrDUBWI3Vla/kShRTvHk4lMxmOgbAWhHN3TrrGVHVlT/b
FWCgMq9QyN0CVsWSrDtIuM2eIsl4mV7DG0OtvKvsgcmXJNFoswLUapQFf9at9TNLTLlliGD1/G1V
zbuGiwuvN4XjA80h+xUdbNfLbWURCSQ9SrKExQf9biH1FHCnaIArqoeZhVJvpolmCN/X8tE2KEPl
O/lf5b559l3mNakp6mdR8B5zUu4Hu4X1XYrznmYJewoSr2aVmgcsngGEmJkr8xG0X5//1Q1k5TcQ
Dpox+4KhqxDLvZELaIoMoIfejkJxRcsepFP4k/ItYPQMPQmT0eYccjzE5EtOwe+OT/cyzYDwHS98
iIoVntNZyxm60l9Z+ccOL7s3rZyBRJK8ZqlBsliOSaLiaf9rlQV0EqrEQpy29RdRGrnl0UDkf3oE
VEcnrQzV5GCf4Zz/Obr2hnQS5SvU+AWYuPt0PwOO5J5Hohg/485iq7GegXvsmypnpc3qNbVyzfE2
ybmWpaxeihPUvnTC7S/QIS3bcbWmAvG62VrQoehyMC9zWD8ep4wIGuTrKs3vSdvjheDMTTBOepBn
HRk2ni+q0x6/wMdp8HKlGmOQZkjDhnte4CqOyuwqUtTVDEAQCPCtuLg0jj8S0ZdABBSpuw8UYMhB
zEUkindZPSjgRrjGvAzOHg0fWODzfex6b2XnTJRaspo5Y/iZo8y/sT3pPTrGUgOudAYArU7PKmyA
Y2VcNdOLXDsU8i2gFYFiWrRlxYSXj422JGIgdQoI/v5AkoFugtHaKRZJXsTYbKrOTiYYn1QAZiKA
OsJPe/+0VpyrTICHD4ugFByoWFs7SOPTxYTP3EIpeAC6wX+ozNCthDoW0HhIkRY+p81T7to2y2co
gTJBQssiUR4JIrgS4ym911K4L8J0kOK8UQCE1NqU66xSmaJTzOMcF+tFB8Q0//wrNlA20Wemd5ti
u3HwyiOsKXcj29hRNLZYSsSnThmk7lf7N1Meh90aorsFHeenMz/p+gaku/kXC2bmfkEK6N9u/FiH
bKwe3l3gouGuBhirYjeuhGh5VuEeEx781phuZ3nxnQV52UT5WodUXfv31UHsNnwFQm2fVfdoABH8
leB0O2MgR8NptFOdBqLyRlmMKHh6ZCmkkk8sJhjYEBpKBDVUfQMYJAgrdjdljDp/OSJrAUZgEgys
WSTL3spvqJN/+Hhx8sF5H99aK4LDhybKQWPKlDk0t72Q9e0RNvdv4yHp+Ft1MB2SFBJfg5S5XxYm
F6pIu+X6JQzxb3/jwMlCFnZwIHmV7M+O5s8PglW/uRRkPNW3SutNDFX3AcCnXVLZN/eUKJTRA+M1
eAwdAuEBs7tX8rYBTpRzteDVUKwsMqHZkyDmGkxa0Sz2tCUB7Eo9XPcEgtwoUmLNP3qeCgkh7aVV
t1B6z++H67lQom+Yaw2PPndw/ugTYZEfMGjI/ePCX1yYsewlj2KIdclBhqudh7Y7auO26eTDEQgT
Hc22hLqIIK4e1cERyOIdcVGMWNyCf88LGEsFOhlun4w0RpxoVq1U8xpJvOs1DoTRcLBW+UsD9hUx
h9gyBXJleRJ7c7wTCyrmeJZNd/ZuFPtNbTBA5835IVWotwlUKm/OVyhd3OzndSutyfGCXCf29C7I
XxsV5MiWgS6v0tBZbyKKa9re9FmFQEodTDxwgDlSXdtgYU/sGR7Y5CmXt7JZ6OyQH7Ne6K2cNEw3
FYmnvkhFBFXKyGtQvU1Z5gkVUD84LiUyDlIgFni02GO6oVHqVMcE3MSEKdL4h0HHt9ZYWEOtY8V4
9Zbz9ByRiRflYf62Lc4AMn7KpazKQLrNq41fw8OOH0CpJ6m8owCImPRQitee4mdf3Uw72U2BHkQT
QcshGm5+O7gO05Z8u+lCpIftjPjJOArRr89O4D6hDEnjAnSXUNlqEXej7z33Ld2sahKUuQmy8tPD
ioL/FoHTBFVdXNKN9LkUt277Nb7lu6ysF0QbE8UMPVyxu5YYIuIsc2zzjHIpvHA9P+vciyAjnXlq
mJPblxwIYco2OtJIj/0TPzPovo3vDbjPHjfiJw70AItHwxqeDtOwFVtKGjVW1tpWWmoPtGZqcEtm
YisCNiniBDKpvWWr4KRP96Uq2twcczsx0ml40mNBinvtucPgEfU50TaNKfzrezWr9YysbHXVdKxz
CGoFXxsAHzoRi+6R2+F4u5Z6u4xym1ODQorp7w+LURYjFN1/Af8AasdSEKigckad46NSW5LPiWmk
F53zjd3fZu93z+Lru9gUzoa7S3YetXBGga/+l4XV4UHWiRN8ixnlEmoYUF9qoRh8f8uKbf92V2rP
RYRce/lcxpT9LVl+2bpFw4iC1IxVsaHVFpnpdp37pSvb7u8x/3+VMBZkVL9+LSC0ApdpkY2BUJXB
L5SrQst2btLF+vA90itTKaT8Xva2O/yAssIHdcXcOqgH6I4iGF50fGdR+dm8hfQd4NE6ShnZ5zsm
V0kXL/NSwu9nW/118t7wPA6UDazLtw8H+6U0jkvLmy3jetP1WP9h1ReLjpCldbbrLlU1+ZekZPlO
hquQUUHYaIkUswKGLE0gZ6j0J/w2YWjSTWi4btXCfcFCsJAnsFapfznvJA1G0ngyYT28pMV2rIoH
TmWiajac17CDASngi3GkjSb6dDpRt58Yjsy8j8PGWbAMCbr5v/zesykVUwjkg+KsiElu9wiQ9y9C
LMKj+RFwwp5sdiRE5dTOmwS/cB9lY6k+UF7h8ZBPy0yzQnIbECITasGuru+h3HJZcqliomnAJK+h
SXaG00Ljj50hqlH64hZCPQvMa8hd6TBhNte+Cn68rnv/TNuF8KWzHXDo959kLK72JDcOnZd/uFzz
l7K1xEwDK6w+xiFjvxL066e9+FaKwgMuTOSYjbj+jCnW9y+4MrpPajo+XHp86+KARVzYC06b+WOY
Qs82r6HnyFJnX0lbhyXoMK3O6jXUi9waE1VjcBfGEymAmF69CBfgj+Bb6gWMwkxksQVruD0UACuD
b9qE2ElYo8+FYEsggpeHbrFeVL/Sm0YF2MQjWg2uhwo0yHAOXIuqG+Rcu5t65d1h2qu2TVHQ4+sW
tvLrXUWmCeDIeEBmr3rQT65OGVb0wyWN66Osr/GHVaMlC8EEchHwKniXUTkglkb24x//lfPD/4+H
jObpLt6iEMu0GuHJsHLKUpeFAXYOeq7H6L23pb+ztaRLI++mR0HgO2tbAOjhyTMuordmDgZrsnRx
7BkAlw0p0GlQdjNvEBBPvlHwYQ/wVW2TkHU7R5F3uYmjTpg9xtN4iZV077y772OuqbX777AAyWNg
OAOGFYntwjJ4sDAk/5hBoxuzcmEFImPsB9NjDFMyxFIM47cT2C5RwWEgNBx9DUmhQWtQ6D3OXjT/
q0k2hOF+WA150YkEtdCj4vEvqjcoGkMP+L2dPwq0kjUquaZQau6wE/bAWZbcOceAaM/Guxn266wW
+tJtf0f9jgenfYRMdX/AU1NHXIHr1pbAkKbUt0BdfdmvFpS6nzhKbz9ZcnjblXKc/y3hbZI+/UVf
a7ZSrVleY0WstRAquWMWQ4JnRus90Yf3zJLrdtqLZqpDd/cmHwUppOFfzb0II+ruMjad/4DI//IL
ev66rTOed+Rw8ZtxL6Xaapp/9FcZ8UO8mvML7/oRbhcA9zf7qzkIo6ztFB1lOf+t2fo9/ve2wop1
6vkIpnjt84n6yDGOkWW17DufemfOr48u5nFT4XKpEkIqor9/mJ9L0OIIAiaVUBqHcK17cQfPLkGm
cryTAys/fG4cqJsBJQow8va8OAai7FF40Nl4yaDHkjVa5UTUD1z47DxH9zw6B61mU7FoP8yaKNo2
Vz/1yciwn9DUHOybmSprbA4WT9b4Y08LisJKJ20KcDxquHoSuNonRJvIRUn5ws1VEEXT2x/piwG1
V2Bm5fmsthBQfXdRMuGgLnk/LRotcCh9u/qdfcJxmPLlREB3JSwRhWSqOBwoyNvs97ABBxemYu5b
zhDDpY/abyxf0/UEgTlLXnYzsi7ibawKgKj77r72/16rWBJ76Yqzag6XndLqoKLvKVRfsrZUeSUs
P6Gf1Ti8+xkau5ilj6+sMcExpsg/KDHWwz9BZhqa7Qvluh+fe0fOjtPsrz7TAx3H3/wXQ+JrDScB
br/1U9G9VD8rhT0lnQHkx0UhAVUn+GsmmhDweLvQWJDvs8gBRBzD8gYwsEdzto6g3NglBWftHSEl
8mWWPImyFyDhewO5OVugu1nNKl+1l0x4ZhUv7hFY1gk7u7Itb1zSkKftqQaigmc8tTJrSY9J+Bmp
bsJO4fIsEts+1L0oKnO1JU0v0ofGnxJ1qaxn7jiALvajcOlhR15HMlO4kCOfQwAupeuWDPlfC3cz
12YF/YXR0xxTxePNla2SR0NUthXSPGStFmOfYlHWM/A0zRmBGymJSZwPrvMuC6tXSKwjRGpukvn4
//YAUDxxSG2SuxZcoDpZ1kLUTTLz9KH9ue42Mdk71jjo4kJnamB8/ofnrMzjnLxjiV8CARmrpkZL
HVhHy0p5f92NqPDOIQE5pO+rCXRu/scmxdVr3uWvtI/lnKQy8q72SnnE0TE+rassRdoL5OARJBj3
9FIbJs6hXa6d2v3rNwgwRlK/Uzli+OzItq6Y7RoWP3akeMxsHmpMSL5wCjhhKip+U/rZu6/zP2xm
foLgSZfxI4GnWHnJkpn5lLcFVotzPtxSDzAVeR9El1Gr8DJgw8YKQwaQsfoZ8pfW9oXclljmeXqD
MAEPXV5F95IPmOtX52nEHVPWmwkncqyOC2VJ6AdXn0pApInD5lmnCGOL3MjFbfJsoq+WhEFgNZHo
XMHY43jgVsTjWB7UiRCOixX+nOz+ut7aXtmBryo4YkB8djKtWr41ulq0hOoXDvn1sM9nxlK4tYH+
JviDHLmhJAoIyr6nNRH9qjV60DyGcHpZoFN82x+c/+H8u2U46aLVInEOdWZ84fk//C8woY1PjhFf
SXQIqJTSa1/n0lEvKN5eip/IOnCIihMMTbkbNCREoPkrQSApfeSoAiWlvTwnlmkAKSgD3oQo1Uyu
1CODROBJ+Bj+7FQuRnz/cr6matrbLkZBQ/o3w1LtsdCybpGGbVYTJpRPkPZ9ZKM38Fm/2qswFZ8M
eSEOAgMXQrhq9Yu94KhKHOBhBVQwRvNLalYPSgxRkIJyi3vUpHgIelSqcYYyj4JrdrHdR3ZnUrFA
W8G5IkSYGmZFNClDUpOncyg76CD+9dXFI3hUJXl35awILd/CAewlwtdsOn+NVFrhgeTeU/PrmEOV
7tsm9zhUROPhQXaK6QDgD7MXX7EPAc9E2LpkyfM/V87QrorVzhS1ZUwYiBPwAD8WBEWAOEuXjjkA
XRuCpvUpMsRsp5z4yUM/6OWdvJ+bY4apggXu/Wgp+H1ryu7krsZYExWffurzNWfSrCvVnH6Uwock
2p6bA0oPoe5cQQumtlJ/EomY0jq31pv1yxye24UrIJlT1Y+G2yVslKzdm/SRXh9ffqze/WF+M/hf
XBneS7JSwQEm7InbeZLa00J4qqQixU2RGjccLudYxolv4P0JfTWURDlPT+d2qTFM0n/MnzRZTlIT
PpmFBtB/87be/0OT/1oCZmBYqMLZ9eLe3/nEBc2RkA7Cmmfm7752zUYPbkUqupgKfoFGfNz93TmB
RrY38YIVduFgsiVRWcLlUQkQf1E9ziZU557pltKPHyEZ3RkaGzz1igxPONRYAsniqoVBue5MssvJ
P0joYUwnbx9b37xme+XuyfiDs2oftwlWS2fHkGfiDqyN9JQuU06dPo99VNq2glazdrckdAOWlUBr
E3KWp9QpDhjIn88sKGwwYps0cY9XRBjjXJX88Y20M+GTQsD4q7AW4rmx9R2E5ORkBaUOoKgJgCxf
ScUTa9FbsotL91Rh6w1KB7f6g9SGuVN10R2de4TxKvbrzEQYD/hXn1bFsh92vXt710DAciB9MlY/
seVpHFALgL3A20BT1fHLSUpczneaSjGvsm9yqKkHSIbp8+E6mY3bFfVRefmdcSveH21otiQCiw3T
1kX143wz1DwyQcFhBU0wOKYCv1JN0pp+yC+6MwFw+ybG4z+T1iMWhoEeMQck8q/J8xi+SPdjVN5K
x8q62i2IUW5rNofSa2mj/aBIej/mOaYRXB3Vb3IlFm49fA3F9SZ0JPa6MahHZka2VXJGgDyZeY5E
d4vdFdH6t+mvYPeTnIgnfFRoM/85OZtmfz012/7v+GMBApdfDxlt/0DDYVbhTiTxC/a0R8lKvhic
D7cnipdZue/QDKLi+w5COcdhCT9bLfc4le72s7uPAAPj/7lUHqZ05OMVoX67FUOLSIMOC5HPTD43
prcgpwJZLK5KYGGGvFCKufLqL/QyK9QzITxEQ77newByElRrnq/ntWdZME5VyG4WvKHKKSwxYNt4
EFWVjAN5WzQlnvyEMSD3jXNJGSWLeyUnDyYpfAiSBLSdkl1V2XJwXOpdmp2UvH0ZxttvyUZQRuJ+
VBMMrdBj2W5Z8n9mZe/0vf/sY9xDvOJ7LNcaxrKruprllqlTiRGXHNVcxA7beTNRv5W/Pa4Smi1Z
4uSRO0jYtueXyJS4VbI0QE0+bCL2My0B4FeQ2GH7AprSyOnD2oyKS2I1aNG6AjR1iK6jLp2gVI2n
A4W1lXb8HgZXUKZ3ZHN6Xeg8RcJEijV3c4BT9ToKgkeye2q0pTx84zyzya4xT+RjNHD80ncZWJhY
oFDKqAif76u5kf7iA3PxjNnzL2H/oclTfZf38OlN1Xp0U98SxA8cvpZDOEaEbLCKn4/q+uvyBcIs
rwy4KimKKVr5EjMyeGBm5EXUB+vSpeM/EnNol12FCRBKSGZEC10maYf+A4KDmZv7gmk3mI/a/ICO
DtS59TUkf+BVN/lpJzJ00VL7/au9rBkUzRI+jkrfhempBCzxRuz2sJy5s4k5qqK57PW0C9142rwq
dJY4JpgVjcMoPzfueIJiWhRlsJcKRkpGpeN0zMSae9yexkGFHmkQV7klDYW+6sJH7hvM6K+nHNwc
HdxSWvGkfr55Xv2zjri+1fyZTtV7P0mXsqcLJ/2BwbmIGLu5d0ISaK2OIqrACDSESQC1+RVXzUQu
BXEZkpjcEk3yd/JgrONQ1JZjUn8yFIr70YL/kKfoEyLxwIVI2csmyoNyWQD/0HvK8901MmVehNVB
dzYGnXM/UwqgV+ASybpQYtqCMRJn2kH+PduaVG/yO9R0m+NiE5khCTtexDTxVJDMjEGY9BRgAswT
al6Cc+i0Hd8hZotUady4tMROmRl0oJh/eFh+zAohd2HTdV1G4yEGy6fPVxqQjms+FFspqN1CfT1A
2VGZqMsPJOsgcQnWC27pb8t9aleuETOF+PWAThRWK5pLd/PbdMJyxAuJMychOAuzx29psI/pZDIa
Ui36j/x52FcMQufwOy3Wp3guwzPOL46JdIhYTHI1I5kDHXkSmAtXNJMVTrBG6iC8NTmDCKesNolL
ibqd+NHrD0iYKqZKK95Rvc4iAwNgirBRJAkTKsVVGJNRtxKbY1idNIPwV8Z6zMmfMHLrvAjsbOVu
S92jjfqZC0MinEkJDJ6aFd/JqK+6Aa/qAKhY+5UIGhAL5b2EzioAWW1fCrvpgj/cBmAkjzOWwR+l
FryiTuNgdlK9mSrYX15cHZ45WpjXidiiPIOwEY4AN3/eLbvXEpEMoXMBEb64UxSrU6gGMhxDF5nY
2HgWRn+KL1pJ2HsgQnleL1BokZCUm+08eAJiGD6UCaW1sXx5R1wGziOaBNm8tOy5OKSSlQlRy4/U
nhGz6xP593TDu8kp+OWPVlbqDNxEv+KXYxbFWsj+x7NrC+HZwqbCu70aodjTaRNITXGr7i7AeB9y
GD7WsdVWORQLz2R/K4b24wsXnVWd92nti0aJlGM1L2YW40ufiSqsq39u0ampHMXx+JLqZo5J4oq/
Etm8lY/ERtHThHPlUnsA3CZGFr/Jsh/MOyH8Yt9X30Nw0RGASoNHZ+m5N7zNYUqGzKjuIRsKmmJ4
qMWOiH7vdvtVtF1kwn1KTvk+7UeBXrZra3sPQ2ZeBUD9WTqw2eVp+yFmtW5UfzEBpWeqXcVgtOYq
1ukH6aq37FcNyRqWjo0/f2wxdoJydoIuZNbVKp3K8WNUDne4nH5B++UyrnXCYktWXTA7/6cPoElT
WQ1ejwSG2ahpqJ0sseRvfxJ6+Xm+kpDxoKsXW/jqQT6Nb6roBCLNBhiHtg8FBbWbATAZqjC8Umvj
WmeDRhv1EClfVLBGCKdQxzGzGXsuqeNkXyltA42iwo1cbfq9d4Pf/QmGy+TU5eJqRaZ1ToyJndA9
BMXjI9iGfVrNpWmq88VC4uPtjxnByFvgy0hq71ngEdmEdc8PezKcUm+uuSxLGR9RH+T+Ku8z1DC3
zQh5Bs8GApmbJLZc0vdcQax2a54hvkeC5EDaHrUtuYY63s/1yoPA+F+q9puVzvK72mvC+0gVgsAO
Io1xcfc6ACTLK+dyJJ0JZTjeks4NBwFwZmOf5gfvnMPproAm9O3xGZv835saUpHpSzD2V/Yj2sAi
4TzM4jDVOr3fpg3sJPZsYzNnhL4J1a+5XnfPOBN1TAA1ze6CIiVaLF18A1i2C5rrNW/YG3qUBiMm
CD1DjPW0NEzMCLMrPDV+9FxoQhLoFExZw8aNsxvQE0jXsXEDZbRPwBcT4CwVMfowtQL7rIIeFa5D
cnXPq16PWutkQuCs0RT5S5pCqEXGCBjg5U7IpKffhyW6cpkfA/B9P8yOkreQDpeLHD7NGD+Q0RA6
JQWuJH+DgyZxIk1fE9UMEg739yXAIp0FF2c0GaVwtw/23E4jxlfyDAp/fZILAgpVtWS+ceTUR8pZ
6lncYTJ13FAeFflHe6V+X9FahDLi90yvZxanhrqgpAWD1IuRs9gQmnhJOaOhrnFvD1J+yoFIbjue
naLn9+MP9EP5H9CygkUwRW2fHgYX252wlj8Gok41jpwwfg90ORkpXIqgm20YQPBh3EunrX7eu8Nf
kdyoDEmqaEiIZvsNmlM5E5yAzZTNCwLUDvN9jzpc9gUEhw9IIn9Uy/exbG6QFnHiRGDii3uufXhI
ryvV7l4tbl72r5GLwgRHztphlxMdf3hEbLlEANXUWAAd3F7TbUJpFlM40tolo5IjTbsrSiFArOzN
O6loqWdF2kyOFsho2kp+V3+zHNxMhD993ZvOzQ5AN3FTHQu7eIyA1QIHbqJUzMPKr1Ksao7nl2Zb
BNK8O1D8wz89Lxnipi9wG/8XR3VJeqWDFsvw62s5f++2HULuCHXRdv6FDtyMgk7YOb9YmkcAXI7E
EVc+D/+MK2WMePaMz4aQACgwaRgD1aYaP1difovMaN/yaQ3yY7PaVbv2GPFo/4deGof20y2nzy0y
0clbbwURkc6muZy1mD/VE/Uh23ypc46+Zb0+F6jLsiuCniBktS0tEGM3fWQsq1JgJJhKlCoNXdGd
Ij8PZ3f0SC4eS6sIwmZqWcRBJxL8UtHQxcKeZmfWDIvO3bvV96AFKVJtlcA5YyHTekK7BXQrF8u1
toNH2dS9Lu4VAHcfx5irxaZBTjvSoHJNcJTyoZKjelx5SGsLRPIdK41kIVjAT7uwwbAFc9WMr4u/
+VIh+NaSQIlMLVeHpbYGtRyVeExX7ROizzPDpNm5fHZkc8xgLdwLd0FrmBN/fSLAPXabtlO69F7+
ARJ7WbbFnE1z76gbH6WIRgMFSWlN/S+8zAT5ea5yaHTlx0XKpNJKy/um7mUvDoqQZdQUvtZu98j0
Nb13PecwwWX9vH7Y9+wXnEyeMbzgYkFken1ExF/NoEvfsq0p7QdDvKjvre+DhX4OPNTGupHaV7Yx
pQoXnql4p4sA0qspM9Mj0yenB96w674IZo8Eyyng6BlLAuGzZse42We4Tf6Xb25vy9GNwH+MsnsW
NUKxGVd8Yul20UN7TM9L9xcHGui34+iEsy+RaV4etRxHdhwNLLAdXb6/kSOqkHcVHNgWBbVQOeDp
7kL2ojYkm8HfomLFr/LXKwtL+ON0xj0k1PZTrQYF/TGk/c1zaF4StokfJ+hu0wpduqIlNc/rLQ9M
JOdQtUYzj57GmP+PjGLdkqfO1yQr9+U+cOjOnYJmv0i89lJf2ELzeZ3RTndFEZM7NegM7W89f669
QZqFdaifiDngg2TopUE0j6NcHhbQKk7F4eFzDEnhTXhgZH2etjhqRofjYarUl7O9pmB++DJM/mPU
ezKrjfILmH5w/jC1gzp6XXgUd5WAAdEDvGs5oryUvp+8m26bOyLy/JhhetmWhxkVZRIoTfTB294D
y/cXmi7b0D9gmWnvbDbIqkh1lbC9oG3ZveyOgHZuQ/SVTaEbuLl0GS1itzsvlLp9MvbCp1RsO2my
RvjznEB51Lc7VLiUzRLGbkO0Co+tEGl3U7S0/UU+fr9c5Wrpk1jEeFm73uWasOnP3n8dWja1Y7uH
fN6QR8s1Srl1mC4b/Iu8XW8ssIvyUZIpkg95OWrZwJVFeobEqf2RY/9nDtgXm76rXTAD2s5rnic9
1lim7zxwi2NUQfBqubO+21iv95PDvKuycBlONCjGw9zZ/aFnm9NZAhWFT+q2HmThdvvkjZN2xy6H
7OS4yZ32UmHNgd1fOmEeZ0l6ouD9r7uimIqeXykIvRrffdGHfuQ32RiMYNbjf04rcDSH6xZA1bq1
kP4rWI/jTBJ0WYPo7L+rYQfvtuG7PQ7VXx3wiYviJveY31R7CbzjvZupyN8Sys01iZZ0fcOyfH3P
qJytAXefDB2Mv2Z0u2uW0tiq73HHJshQuiSD0ZmIlh0JJSdqHhG+2Lr1198brSfsQaBLvmK8F1Bz
bBdnDBKa2X4m8+JirFCcNBGUArgUU8JPmB04BtDyacYl2v4GOODk+MrwrnqTehZjERD4YwLE19Af
C4ZC7jCmRDArxbtbKfZRsBUwOV3hpvoRIExbyO/BeeJu8knX8D1BO/nIz5hTfSbfsCv6NeNxSRCp
VfyP3iRU9sSaDTSnC+RR0YYGOzYo1HwutQLyHyN+wN9w6oVDRaZQL3oO5/M1ZFKV1gglAx7RNL4n
s5w4RDxtY3gdKrUdFAf5pOKhD1GF37xLJNinSiFqZYffwOLNNiTNUqIrxv0LP61k8CJsKZnA9CRD
CsJVGR2mvyppNh1XMVtooI+s0+nML/lhTteZXl2sQqqEpkj4nm/QiZWLJ9CHGFwgdGmOKm695MiL
Qx3xSkp3Q4TwaA2DlYAIwLy7zhrI+MuGicX4IPiWYeVuaTZYknfJAWoezuQjTY074+34LbWemysQ
6kLZvtDBmmhTm1U5k0UMJMld88TVmMzZ93ltDLrabQuO+Z9TlGrJbs68PnJFXF2CUYw597jE8xwD
qLIdT7PVZRX4ygioyvGwcAj+fg/2eAw49yvk7SLBwkdrX64zlck9RIkTCPCG/h5MIrqZfSnmw2SL
eNYuuan56jXapzAjflN/mx/Id4FuTKLl0zg9jNMxQiPXYyRr3PWYOU5Au3hFp1qZ449P2eeASe7K
DFXG0qJEyTIppp1IsXc+Isx/wpoX3ZfTMX2r8XsSCbyP9KSh9CYKKkw67LLKq8oWjTFV9iLOi1IK
O37qxXoANLGk2nchtfrGcRifltoavnJCe6KCxZpixVrKhF9MBkOxnDZuatdoJJW27vxIyE9aJWja
4+G4AFDMXxoVaf2qbmqd86XnMQNsdMuBJRarTRjdBiOqJHizH/M+eVjG/PO3OMrOSEKfYisbgVmR
gfwVrZtVY0oKVmvlbUX0bJQ064orBrLUwV9uJhDW5Z/xhu2sDpBFrRSrRcH/Hs0+R0AxkxbgIC42
FjVdKA+ON8Z7dInoducvuUMycF2fboCU6d/FXLCwIF5/EpsaOx5Lp28yQf4IdHmlkEL3zF5k3PRC
Gj29YBv6SK8Y0toXdjNdlcqtvtMeZVNmquTAK7reGuzkWDXVADa9lFg1kUZmyZoh+1YUqreSCxvN
zipb/zbCao2brk0V2fKS39/R3IHphq2GX0mnZ+5FpywXIHZHTAFMBHSHuvPvHWZc3vxSFdB5Ra6M
m8pp268pX6feHJvvBiTQfXQBVw6LueYAzmcMMHRvlDthyVJNflp8v5RtkUqegRGX1hl4ZdXpnXHa
n5bZv559ngetpkKwEOM9SAQOsGO0iONaYDoAuIAAmIwd7OYRGIfMJQIUaSkbEQv4JiGR09dbhSJH
YkW7BP5KRtp/QCL60t81mA8b0cnOesmQGXEyL1ROtA7aAM+J6GAase3p5op3bYebhDdopjL6snNz
+moD40qdMcHJprinuVdRt2/RmiTkcwAh+Sj2kGmSnoGVVjwpRQq7KCgkdhAZjGvW1hY1K+bj0Utz
mnj0Ehf335Qp0v+Pjvk5G71TtPliT2u+J4sfhNwRipc3e4XOsoG+px03d+mUkAkweiG1+7IfCEOH
LLU2+wRPRPzMxrp/acgdB/qFO+Lt3u5Y5fX+dRmjNwv1DdLDU5QVXvhApNGJiB2GDqkUhpDjA7ey
cvb5kvQpHbooohSQbuf1+B8onUK+JVjZUriI5uHTv0QoghbAE026LZHnomHF9r+/EpDOimDXL/HJ
BbHzfpsZN4B6ipL8g7a1eAEqJPOiptx5EuDKqX7l9lxCmrO0hNRWHdzUfG9pS2WJZaEpTyc5x06u
EdbZNqEh7AysupTUYvl6A5XD0yGAzOvgvp5dfn1D8lERyfLyrhmCQWW9QPdl8m0oE3fed9fDlJ1l
P1hVbMzKuQpQLiArxP2MTqThqRujrqCzga+T1VuY79pzE0n0q6rvbpGXtsZGyKenXnolZ9kp1E/Q
pevxXdIpKAsYLBbndmxmi8ydw7fSvNDtmW2p7QBYbFW0FmlFzJd4UhdbCrzPbxnDoFNIrDXSZqTR
JP78vZ1xhZ3/YZBh7thppfcsELjVgKg5n+QHSLXBD7GB5+TY1Gx0/LDNp+HI+XEKmiPi7JLagHwu
/StS3/1VKHE9ZtqRb825JNwcSWzAeMJV9k73pgRwuLTbXtCRlrZCW+4LxhgNpnjGFNTpHcUjudjx
+NeOuaYgTqNt4Wqd5Qijgal1NKIzE4P0RSR3aT8WhZP6R5EBUUBhBU7kAxyW4Exo713NqMnoaNrp
sum3knY7VZIHuikQjiW1SRFS9CGl5IO7MIjoedOf5bjTT6RwNQj3QPCJ7UhsApeh1VFAsIZDhKSM
h+mwCaNp3JcV51B1KqEG9yPEm4nmtt2GgOPG9eZVfDd31rKRwl3i33rvCN/7zBqsHFzRJTte/nEf
FMmpknffSRcyHt2n99NwPtbeLNiapmjc77l4AVl5oyoVsABNg5W5fwU0Qd4/evGRVYlhgbD9mUo8
qcqi0+KC+14lD11KphU7fK5BwpnguNkakV5ma/SfrW5F5lV1InBk0H0jBVwcditFmbGiJO/98Aiw
ILwgU+OzuHnCUNx+Tc8Nk75cDRQ2BWcWiOU0QwVqGfA40EEWiHEtvsrOHMCCI9gJTcv9AjJNJhsn
I8OdeURaigy7+zgw7m7f6LcjzGTyzTnulBM1ZjOBNpCpvVjXiIbNx0G8lHrx7koFvwwJ6x9tnPBV
QVL3DIWffbqwrSu0qY6tSSGAsblcionLIJy8YC+My41AVVPWdRmizyk9K3K2oNpDbtAG+VI/jNm7
6AThxEj7cExLE+1t71MhIGJM2sORw8JWXD0qbSSizvFhOhrjbY+eViER39++z9v337cfxopKsNhW
xlL/IfyI5HFz/j1oETJLlKyM5j/pP3DFcYExqfOQJVi6V0D0vLKxzP6vSl8VH21r3vvl7FAKsLwf
eXnmOma4mmVZmyOthfOh49o5WvDqgBk1nd1t/Iij/74PI+OdYrzbCL+n526Mv7RGQ63i9/PH1LGq
zw8QMsoklvAyqfYkhl0tjc7A6NB8wG+pDHNj4AMrwfS+Ol+kS55TMlCPURoy2pHBHSeqTatLcuvl
RVgEqgJXqEycZR25OVhw0K1TmQgdflJrd3+m9cI3MOu6gCdhBJEqosTvD71Y48/SzBiFSWWv+y91
k3A36sd+dMdtDcC4/O6d4V9S8haewW4f8jKMwc/Bxz7C8xJbRmiSBwvFvn5/FLKymkBgxDdVaDy5
+Lxf/GDyip5CsV5+grH6VTk5s448IC0lL4QYf2ytMVM5Wsanf+Uc+6ZTCLEg16dgyoZQselay/Mq
uN0u31XxU/iVXVqYEvYtlPxS2Gey9foHptkf2+PsUms+T3MT2RG0ZLFns6MS2BgE9buy8YKVS1MP
mCrWbi/JOgiNEII1JmPle4DQC7nFwwh8vAkwXx5A8A6NmwUeoozKOyeJVl4syFRgMo1gdYS/yUgs
D7cRNlQGB+e2NYHo96SbwxKCLYOpQgIG5pC4Hdz0iySHfLcDywDH0nc4xGMJh4ySlthMxbrcuVrb
6h8ZhtW7BzcsGX3g8goKsHcVPkW5jchuNaKb2A2zyCqVx42+rHFuWK/zsoof3ePhEYYQGKaR8QRa
BXzNPh/m6BxhdTn9rqtprbJWbZWGfQRie/vb+liIsUZyXsiiCq4HZTIj91NjmdMahMfXE++h6sLl
jlVsblPlFDlRfb5QEUES7bpWZq3HH6/aT5u4iez9LkeeyQL7BcrN9Rg7q1fHwNKgi0Hy/x1SztbT
xlWuAYqvq0+X8K0oGESgBSiLw3tANMGWu0YPfeeWsRk67xZu+wAlUxVz88Z81eo1lWnrOEc8ya1+
ptUiMxsD4TR+6AGalQsaf2ScWPxOmk4m1nzWtSsG9towfvKwANQl5bkf+BZED4XUYlEe+eX3aU+X
ywUVM9FhzMsS0r3XiOrbxZY/p0d/lYbMhl4JNfcMZJWDzNoWwEACpsmMY2bEkDwTX+FjcmkZarCQ
XvKZdfcT6VfYLXbc7BxabP02ZFB+leUM5xa93ReeD07xThDEcNsEVGX7YgbsmtfWMGQwTHvAtxMN
Z8VGgCMks1VDfXYsT7hOESufeCXwkSdamI83gxR/bkkYsQnQt+eBHjtcgSqTHipbkbHTwqvf3fjC
awsxkswe3VGEYdAR5wip3glMeFx//RRtkm9pC8e7iRhvLxXRQNYh9bnLhsp9y7jIXLMA5GDU5swV
r1xVUKxd+Qvam0mKN/BCSJnjDI9+HOdf3kww9svEaU917rqY3NAcj/mTDjyrIPLu8rLfASPoppH1
ufZCsM3pplVsyD/E6/5crXmY+f/2it5d12F4mAmn7rwzCg7JC/KVW4jJyxzV4clysFRnPNU3xf2f
ZgCKEuJg+orRnLQ2J+Xc0eLJ8YveW3v1Ztk+5ig805XaFhM+2ov+8fALqpc3B+xy6iF1EYkP48qP
Xx7LI0TpugrZ0B2kWzdCmp+5Ktvddjq4cAdLhNEgyoQiVRtvmoLUkV1I09krkZFjs05gfR5tUzeC
/oMthApyMInD3DCZQG7aXS4S41V0ciN9pBKNUYZSY/iebgVRjMgXWrnEuf6Je3R4fW2u+CGJ/27g
VCZv/VRePka+GxHqTqjOVZmUORFBw/ivx9PG55YzaXxbpqOS48q2XVPdm0xNhdHVTmxsZhAwI0BV
A5g9zicF3CBZRO3Fq4t8tbo+24c5/ob1dkYwMbgGKKxvTN6xrknRmQCahGR8BVIlB5yqXuuMkmlP
l5kxc4Zpx6EJU1Ux+BD1KnhkuHnmdPt9GYBzjTrqvl/IiasGofrVf+1Ca2sejyEYKMI63PeBDkGc
I9lZyWdVeYmO3Y9p6o8aYNreQQe/D122UkPnRMoLKQgOe7xwknK3GcLKSLBbpzHjlQH89jQt4cVw
+Z8SXs6ubdpTFY4tTisgXrBBzN2ocyTnWcKufiYb5D3ToLPAO2DXmwdTG/zOWKpRKekSnuOJcqPq
9JA2ysSVWyXy+r2wuBdsUqAD4q3EP1ZUKhWzRXm8NodEvZo5y2ahRWNkrGuPZpfh4BSFMYwZ9KW3
yBNR3JabBOMm7ysSHHjXv/8VgA4WGNA1Khqamd8k5zLSmvqD3hcFY3tyN3CEzm5jGyHAG2PRSbln
fUAtwk88qrmxeUGig4nSSOFB2/SRBI8iBfPdFROb1GSrwBDGyq0pKEJua69PhAWrzk83sErPaAZ0
lc/CQ9kuKlfc7+MqohJfppXXX5pGpykZC76hxiILHbms6t6o3OJ9eb1cLTpbhrCXOPrFtZWlVj1W
AlpyVYi9M84aFLYfWpq+s3S5cNQ6LfZFEf542d/aOoAz9BVm1IsLx1ePD+nVH7UqclESK3aruV/S
8yDSnydBPBdNU6z8VvwRW/Bj6m7QXn4SNXw0Kdr/Kj3vepKi7xy2oqvLbMDNzPDn1+GieGafxEVq
m++A+JW7VkLez4Pkp6QNIzavnyZYjc/ND5vNvrAllXMSNlpSv7o6CjaVakEOTWJFyFvnqrmDo9hS
XjvRWFCQCs3KRksIKo2qbKJEWLHIx+jt9By3Blemy9qgbc1RmBUgqMYmds6XpH+O7BYOUMuskTg0
DCn89hX08pF9WRrTZqGqjHYDywMVunAkn5AZAqAF4JllSWFEa1dANDa9JVs5XD1SiD8q1TfpiI3n
Pp+DcyFbTKvpH0/HHbi0pMn58AnmiOCrZxgSwuAUYRPsxoLsCGKoT1JP0DJBzIMfNRlBoULg9IQc
JWswMTrv/cAj6jxMROkIn6EUA6lfBXV3Qqj8gYUIwLG65gymHIsrccvXnfdUOa0lFUERQZwlJ22g
T9K/xSzTePTY2pvowojoEZJvLlzNZFGxnMTbLWtij9pMx3118MBdB+idK4TeXNVB7PaQFUM+2iaz
QlfpSWrlHAL6TbVZQxouDSxlIUSTWKYq4zIykmOvej/yY3AsAEc6CWrsVWGFpleLVPdeuT34arZb
VYscFRzN69ESj9qVE8VNf5HEXSqTOtVHbMwM0H4nQ5Zki7xxygp+mehsP7uijfVtMPIRjD1Kby1K
XvJQ2IhsLvFaCgoDIiBqGIcw9cKD7Pyj6siuk53lPGRK2Vi694L8gu00i2k9f133klFXvgIANyDM
FlpzFgfphqdvl1jMw28kLZL4OqGdSwyYxY/OO18VME79/OqgLfbCGjCWpoKTPRxrdcelmZfOLXOk
ngr2jl2iMRnhgu7QNoe+BUtaXEBD1mYQXakxuWcTmrDhlEoDZE4DooI/5Dlv1SLzAJb7zld7expj
LLnzFc6ufOoxDNx4kp3dadL+j3tAiCVaAthpjeWlmZvJokmlS2DanE3ovfp/C5Wgg2kb9UhdGU+B
C8lXui8iA8PB2rJHA56v4CW4DrIORi0+ZFf4hbB0FT2bs8qXZ14kHO8yYjVpAlsbnO68enug0LTv
OpHX76Ve6NORQLSBFW+W4zjMHUK1Oy3OfQNPPlJsyd8jbCeQWeVbA5JLUZWhd4t3LnWEt0l8mBdO
U9egZ35gO0hn+kokYVCTYOYMpNMWR6UpaXTkwWS2U/Ed8vhv88JdWkxufaFVMyKCo2YDsD1nGklW
1TWKTPkoLDsSOzz8F8I1TLsSuePMcqeqsYzJRzDd5vFx73zMbxK9DZqgxKel0umF5CbwY7oJqiPC
Lqq8xg+4qEVs58crNW0buVOJo4U4Km/rIDe93Duv5egkem5UB48JKtkE2VZEGFuojbXvcZfXpPwV
9d3u+CxOG8Tsu/61diPBgJob5Xb5GTBrH7Isto0z7jiXsGPF+Eb5qd9wUBdAIEUcfdM0xtcsYiNS
oSFppHGnn02yNOJQ86Y8tyf69u5x5WlZxEk0HZQOssYHbOmeg9a85HcC9OTGfQOhqjPc4pAS/41K
DIf7v50LpcWMm2HAvgcPPy4GMz723Oed3L2N+Uk4iJIMzLr77kWBaekGC0Qy0iRcBcfrkCcFB430
mXar/7G1lh+sJ9MDIv/EAbcZHJ5rLLJkICoNzJWz+K83IIw48qZAtEWrGe3/7ydGTqoduUPjMsdM
1nePDskgDA/oFYiJt0m+IzUDpFiAfBNICWFnpPM2hYjQ4Z5lPzd2wog9tPE4E0tlUHxW3jcaYJjl
7n7917tRh/MpSf7mFp5tKDN2k+wjDbsVUlS/FlFPj3h2X2yPShjAPAc5c7i7NDwjwi5cp2olavGc
htyaM8DA151ZxfzIqOgtXzAG6M59Cx93Ws23CSLJnImCh2bAw/EfQVs2Ka4dN21B12J4X73zSbNo
brjY9hAYQM8pKwE7TlWpB2SjX3YJGX3yFRJsc5e6Rb4mzaXmUv50S4Es0aHrvhhetoLX1YyaHhGi
GnHRG9UueaTT89yoZtySUDIl1SDfM4+NQka8kTSzNJsuBH4KCKDwbIrjWPlnvSV+53yufCUKdxyN
l/WOp8UI/XQXjMx7l52QJg91ZfDrHIxgI/FclLWKlmlx3pi2fItYVC4gTwpkdJF1/hfj0nn6yUJV
8IZ8LqUi5yOU6irQzXO35Lt17ma8vgbSgxnb2s0tNa54aalxJ4QcsAVEHbfgqpCECa0S6BzhVz0E
xqNy0u8skcbtdn4bUW9Ja2oyIvvz/EYZtD9UaASSO3+Y0zNCljx6Q919dKoNdAoIPHmFhbnH86vL
A2n826gOkPsErc+MkGKDYXgr9EuzoSbxUQeyM+oHKKZTeLLuI2/EL6rfq972wUZ3StnSg+f1F9nk
PKH/7yxMT4kW88Xm2vsjfffBNHt648HI++Q78OsFuT/rjHnk/7OOPQsRKfK3nYRRfI02yVoZTZDR
sEir0XmtiRhmkCkBbddvMWb+33FHoabeIc61Oqt0w2eSYtSzHd99pvJIBha4l3bMI1pB6m7qes5L
yxd6vU2F/M9loqOKCdxpwXwA33Ssy5fsmSpoaW4G2/QzPWjE55W9n7HpbsqLjNFiB2VCnNZPCgJE
G9Rh0HA+QMK4DEuFmf7XtfEcgg/qfMdXWrPzYDtSq6VDAjcVHa+UOttyczx04xwugw2ans5KrYAN
KScdx2ejV10JHlbbqcL0dZbhN9LxL+yjI7KuF7ftGv4JDOXWz//Q6E2SwifJ4rhVRCBB+zeRxewi
/TGHbFDiDBkPn8a5gMLq6qVsfe1YwiJWbUH/dG4iAcHHjM0FkqP6NW39qgRQ4Re0gcq38v4weO3R
W6ErNc1aeqaQ6bx1X8osUONThMgP3T/S/mVcaGzmLqCdSLCnh2CLe9bzZmxdzztYKBbl2oJ7DGvA
4HVSU+gbSEPnwns6OuIaZy2jH8feXZNXLokq0RGA2jh9XbZezAa/5u0K7b3GeinYwyniqtQRrrUh
kDPk73g+gYoEQP+t0HLXXBaznOwkPsbTJadQFbgxCC6NYfLUzNXhxeP//qn+a5aNsU6uzf1qlUgG
nkPTvCcYFeZUIvQ7Jan0iImAxBnfE9d1JwIo2q3XiIvEb50PC7/AzP5gaTzkWaNTlMdewQ+CU/ob
sg9///A3mA9kFmf65jvgagCxBOZNxmroUFL6aI/LUDN3UY2ou4Z5LcEK09J6uKSBDQulpthmFuK3
i1L8qEU6cvK14+ZGpS8Wbd7u+fNH+3ncNkUh687yocj+spwGvusgeVwNEdwHglse+jBCehO1Oewc
/DYRp4etpWzEKDqF4N7v63oRsB4C61u5nu7r1gefeItM/SViRKlwNP2R9GRCp97Z6Ibov2yERv35
3W2YJBAJ96fvZzw76z8ie7MHQSlGdF2lv7HNvneHQHX8wwU9+aiUIHdweou9wtQn771Zr0IHz/tB
o/QINB0hbzOu0P/rtKrTSyNSIRQr+HqpDNFwKqLtSCZ/0HkIUWTIuqV58aZsJ6/vBrxrSDoUtle3
QyqMS+JHG02WrodlgTqtOH7rHP7O4Kq5PRhpqPnFQt54TSos6Nz5dq4+uYRgDjiFrYrie8pBox8f
yXvtMDbb2wn4D9Lb2E/bPcTZ4SSG5uAg3XH8NitD+Old0gcpkGNsizhXfSYDCDGw0SLi3pyyesY4
tffbOeqINHprYNX0tJTI7Wek5ROJRytvxhvRQRNcu1MMlti63dIXyRKY8eZu8FR8ikk+MSJITg4H
8/emglGsC0wNDpRyUJiHjaDOLGiLlPJsQF85/PyhRL1LZRX7chu/JDmXXYw2BugU4rtAuTYGCWjn
jgibwPyMtBXZ6XSsdi08pQUec2Mfo+sk6fIYz7mwukMf4XmRSFDO3j3hT1kASHkXbGmeEBWvde6M
MLrW5ta2J6Bni6Dh4G4dqlYk/pGV6p3GOw6tQkgl9HVcSHegbwPCvg098BS3PSkfKgChzh31PAP+
JY7fiuQ6sUu0PD5yk2CT/eKxZ/4WdmIPPyDNrYFS7Jvm8E3Ry1Fv7KebmaKEZ3SGVIv6IhCFAKMm
riHnBI0ff9EtPsAm8nCeCKAzuCeAZPdvBrmAuzdUl0k/PtPfObcK4wF0Xu0A6vJJptUOT3B441Ty
asx58OOFPKoeP/wW1aTZxzPR6UromaaYdlbdKE8Q9ZA7FWS/MQbYwrX/z88ffUSTmS92/hXUbzpH
DQtiQzSmb8CI1PUxlD0OhYDXV4TeJeV4oNK76ug4Zazbo1+zkG1CUwrRo2kYA6cC3VBzO2tYiYwW
suJoG0JjWtYjbp5OuJuwSZ189QrmY7771akxMkubb1TVZRVFY78UawQDpZsShqB9X3rMa+1cOQ7p
fVcdSuBD2H5EogvNlVfxSJkkcrFatTWEWTzRTdoGGP/xZxkUILTtpFK4LFINfcYI1bCQW1wvI2Dr
myf0/zQOgYyF7aFJwotUXzy5eBRlPzbM4Ae4XsuD7OD37CZk3kRhmCGBciBRvIr6dtQCCmEy6SLo
uPqtSwB9vSd50RvrQmhjU5QQBWpbI03ZIAaWGh32GXDnzvhUttyv3TslMlVreu9X1PDce+j0WnZ1
sUe95O7NrHwSDUocEwPY45ZAxpobncKZZt9RPM65SFR5UwdiNiCtmoubR4CUHBbq9ok/4WUPVOsg
mdESKTY3Yo3tw0U9NdrMJLBMoEaHeud0RBDAom3aaRVuD2oJn98b8hZhvd1mseU82lsY/DHdcnlG
Ma+uPsH44maSdHjd39HbFj/fP4IjsIhLErRNhadu7lFVqBaFuMistWW7DpszFwrdUh80EsbPs4VH
kpxWNrfololJwgNcWX2j4TkeIjfigzTq1E3EYZna3gr4tpXtKho1NCIU6FBcd715E0uwYwGbV6cj
B6Eu7kcjMDzPmy1IgsJXgz+14xveYaSZCqYzaKU19+84cCaA8WG+EnIX3cTMRmnYPGINaLmcrweo
DdQf0h+yx72Yb5EERZY0aytTp9MxuP+09s29lSbmKJaxrfatcYkuSS8CMHubniWqkpsup3+uaFmt
q5IDZ5abr0ZBkO+drTidrRU9eoIgmeS85SKuaARr84JGTQ/p3ysSuwatCSTxwI4MvjPudRDDgr7J
/vw5xqxHmoZ1K46oEG3on6rQBiTrSh5b2JvhCemMr4ZuvgUmOijrbuwK//Yd14z0q45aGAwHGOQM
nzztiOIwjZcQ50tLfhMDZNXm6znYN8xKpuiWn/OWUda9SwKpJGHeO32T9w30lLipR0D8aNOq/Jbr
VBUTjo3SmGA8OjopTq14G0yj7gFwsPSRY4JwY2Up4OSLfIsDYWQIsNgxBj9X8GbeOKy1htEIgpOJ
cIk5L6KGOHcFyCjtLr4XIwnDCVjHDuRjlbWwdjMaVEKH1RTZnBmbodmN/VNNQj4RzdvLE6TjT00x
zBsX00VH/+j7VWt+1rX0UjLg3OtGTT4mMoFMTwZHNTsITtU1TvOBm+ley9/QfHuu3S0SmjL55uW2
5i3AssimScqsWY0dAJaqnOP8iPs22wpyeS0qwUNP0vEDvsiYG+ocShfOdAim3ay3nwOgbYPwHXMF
BhbPRA4cJrTqj1m4SL8S5K+OlOCqajb5L7TzxcC0RxzYonf8i/3snXE6JuR3/5Y4u4W7QnGKAZhj
Hwx+ELxhWsJAhdTRWImW7qkjmf2aJNG8K6qoc/DsKNWOT7vhSXiD0gUI9YjY0o0R9JCbn7W16DBC
Wk8f2GEbBEo35HPbLULJsMEj4LzzHSC2RD8kEDzFusq5He8GeJlDbK2hxpD9X8x3PeOWINGj7byy
3o99+6NhmwY4tsws22MedZ1gpM9fb0AVbcVwn3ioqz3LSIArAAtaVQidLmgdhAMsV8mGLzjPJpPs
xrXYl5boA6nfzg2tGzCBMRQ3iIr7N5JBdmun9dT3wgxO+yBKkfRKHV8cLHPI6sD3kxr3vNEL0Xmv
/HcvUVbn22LaKUi5v+cD0ELFlLCHAeBLSf4B1+q8VScJEyhJzY6EkRJwWthDqpoFxqC7rSaYd4Q0
KX7C2c80gBadf+d+trppWtb5MmtzWRpF7/IvQf1SSL0sqGuvsFctJtKxxiIOma27oNxikoQJ/FtU
ClmfWVQIUUTTSr7qRUxroKgsGfvMp4titgGZhKdu9tuiExxyaIVdFyCCKBZXFyelC1eBy4o/VWtw
lPqUJ/e52YFOFyrpzuJDvHvqu+RwLhAioc6dX/742rbTCSZsg63anZk7nuabXVk4eoliVWlu5N8z
GKaDG3a2swjciYTYF/j2Jfpxh0Wy9/OIWhSYH2gx5Gj01IPRnVeSAywctWD6/7yFb/jttfTOFIZ4
fHYypt7dso7Lh36U5rziLM6P8hahhuRwHWXhlAMhlP0wnaEZH7BOHXN9U8wF8+tvL8jiFLkMp207
C7MZQxnRN1ZLd5RlKJoNR3mlRo0L8bk26qseYKAfxYBnXgZCpyZHWokfBydeOwasJELUSwT6Scgi
R0GMhVln1wDbrXHjagh1ewDNHjoC2QB39AP8EsxQxw6nOyBDE9N9cIPlv+8L83iUwlhslIp8A3oo
/WxrXzTDfrUiUQBk7jz+WBHptEuTX9RY03g+ck/NI0FRZ9bBD5TrHcdjghqvY9qcdcMZFMSxy3H8
34Co5W9epnnj6iOQo1bdK/bucZKGSSjW8ey77fZXoJEefRXTBK3H60O+dhNwCFkY3d9yYFUjTS0U
oFOsJxo1RhryzIgXiXZs9iQ40BGbpxbdk9oXWn/udBpd/rbvjKQA6AgC2z88rILV627vI4WFoNUA
BJL8FIKc6GqQxQJ9y1tF07cQadSaZpPo2SbbCq1YKzvmLrmyPrOIl2N8pW+/+7lhs+hMpks/lA2d
Sev1y6xvLjuwHR7Nc0FQ45IGEiw/CojZCQlu5vAZzqz5Hz7vhN0lWRVPDEO3fO/QX74zOQODKFOg
Q9UK2HFXY+qHn7oWHdDQ3hEJKOtqPqbp+gpd2eHD/dN+b0RNNfOOoEnrouzBkb0jp6kxpJ1pYYzq
gfsmkv3/81S3JNVt8l7+u2xRe2xwXXCOyjzr1T9mpKwSYCe33VxlwMsuctBAbmGaArK78ZC9keaE
zgvre9U3xbFBZLbkL5D6CG9m8i0oN6FX8lq5G0yY6EuBGvmUA+V0icAdX4owADqPuH4IrE+GdZQn
k8bFyFOwbqGr0USzXqsOgZaT7ubNuAsAArl3kyqyXeQUDP+y7NJgpdfIXU1wyZWBM6wEB+tGFtFb
SoepPEDc+xK6AhWp08B44bAp0/iAJ43eE1DXOnRDl9KKKuxPjaD9TLWTPxTy5FO0GJjv44/oY/Qs
r9E5Q7vPM6D5L31ZQmXf9ATR0rg3M8MX/k3d261B1N5q+uUIMZn38+nd5wo7fK9aLvpDZ+A7lG+X
t75uksr+e9f3w/GRCKY4T450+5OaEi7S8DF8iVy0+SneGDWP3jFhn2IeuMqSbGWpiIp9hmeGeMRF
UEWXYwjI7lrGRai7f66Hs/6y39C1GqX9k7TBpJ7nt1vuB0toZjONrOyU58+5GTKmFpee3NUO1HuL
01XXy6lUsFg0GQZNou0OTyd6tN8cRFIVe+9O6NwZSZJK1SHPLqLJ73HVBEm73ypF09BKlB934Q55
mgfa/wVpHz3kefPEc6zcCkNj11qClQgY9Ic/0I+ry9JrBfzAHtNWZXCwV9Bdmu3O6W8NJvGdg4HK
dmAYE6twjdoGtRq3gevZQHeLBjVlW8gsKm/n4Meo1OvGPke9dYHMRRIhw/w6+oKbaW8wERWAeiEc
i9FrFB+rzd8xS6hrJbR+F+8RSGrZ7Pal/24cF7AGeo7yU2dVK1u3ApvWAOxYFWL+OXj6s+OpiWQx
A/QoLGVln7u5BI84pGwZQJ2dplV245hEoA67bZAFxvt8IIqfOcJguCh/fRpBTu2seQKQPzJ5Umd2
fXP0mYUWpPa4zd3o9iqunLY2wh3UhEP0ACebBGYoJeh/kRLQ1jq2b5Q5bnWhp2gUbBrt6u/CWXWq
YU79NdwUL4e+yRTVEBrldk/8UkwBUZU9HSSFXWCN2FYiFPCT6OlcYs702jMUIBag92cic3hPQDlF
X2MRQyUaPtU4JsJYYzvsQ6hDDng8lS+H2EcSlzFwD/IklgM704q2tfmN6nEobyEuJeiMgGCKnODg
Hl6BVGe2XW/f5qETn/eERas5aEHCnT46VJM4qcO6w4hcLIQzuamGNzpgxSLtHXPkLaJoun2lI6p0
gOnCNrihfdHg/sTxsvaEHR+S8MUa6c5yWm3ZnLHR4xhan7zCZhcUbpC9sp1JYKGTlKj0qesJ8noC
434EChRLLALd6Y0yXMGLgStysRVdoZNLNCu/d03AMmyWTCK4ezwgm4hWfsEbWg+V+hlIKA1WSBvE
gVsXpX+6fcELWsJr9Dc/YgmNrP6MDfLi0AWr1GbE9PsOgyclRfQYTqY4IJCQqIRvd4SZYugt1z7M
yjhu4XCrrfTYfeQuFY+e5yCzaIoMWnk/HXhkeigrq105lfDbQ4G6Y7UQrgd245CrSZBiO+5Lns8J
8H68d04HpHoJNgnLL/aL0TlpSgIuAsYXi2BYixdEGLNGRsf5R7vrdH/9sAgjR0uwiYC+O75Evs1Z
zClMiskRsZbgPU5UvADT970f0RcONOwncvJKnTDMnfYZHvnjhm7K0CaF56jbqWbtwAo3hHiLUtWv
Xrb+5FFRsBmCfYbbb7H4nR1A1ZMD4MtrrPDNeaAyzJHFFmLKUMt/qoNOKJ3LEolcmU5spcfDgszV
sMXqDb4rtrrkykL+UhiraRZ7C2yIjYhB+uoLY6HMi8aLJYhxFKqlYAD0FFfjZqccZsprxbfCcSSW
U3xV73EncMEe4HYHzeRLbbcTZV1jNT11W8ADy5rBT75V4oPDZV20ePIYHNVdhMg8mjUT7ZBpeYQw
vU1ZzJxnFLLqjkPg5OlZSwmBw5kzp0TpfSHsDu5bxrRAGK9Xm9/9DnbWLZHu/we8qORwYh9hXs5M
oAvZUMQwNEyAj1+3/TQi8BBR/x3BfceiLU28Cwxbr1sHGOK1F/ua4g1PeWWf/WCR0AOIlbfV4/TW
JLIAGokYBMXVcnbr+Y6BdAp/DGMsH27bVxfba2MzfhqB5u8ZHMsxd03Yo+7ntZHanGTv2GtYkmr+
cdn2hTH10b7jKHg8czIqS5eHmSnruv8jcYVqgmNB1IB289ImTLEc17mOke+PdE2vVg/VKqQUVxwk
oV6dSYjNf0K/FDJinj9SmDbz08hMc19AXRpieU0f7ZsAnmeyDrmxA9MnETcp8D/Be7kAodfFy2pZ
OtSmbFC8YwxMAwC3dO5H+X+1DinKjC6yfELG9ZOG8BMl9YxVTsFffw2e7TXH2wuv7PeQY6/rTb8n
pbQE67U9uQgMQrwmDrq6HTL9bQ6nWweXd1+nSnRO6PKeI0iaynT1p/jdWi5XL7qBFk4CdSLycvB0
/BDBlvFVIuMTcwnSf52yrKLDxhWeNb2pSNk/nnZgwF+h02QACIRoK5fMvCqXAV9AHekRcc0JItUV
ikCqMZQLxz0M4xCj62Q4TjnsDpgDcY4haBuiLsvqiHS72nXtlpZkKQ0ElHkQd/OtMCzc7ZSePkfC
/Wq5o4xuUYkCK85wI2i+g7gSkYO9Eu6LHugKFcmuei30Y6HbSkKTA6JzyFer/RK8sUjrkTc+ApyI
PLErJG8+croxoyMbxJYo3rLop2ZUM/y4Mcsh4q6+NbxUT1DKEgFcmXvPGGYCw2ieFSF0e6efDbfr
anHPG8tnZ8PZfIfm+rEujfUtndivWp1a8F4ZObRpBS1osD9QtXBRz2zkfrs81jL0s38pz99BhMUE
l1qYsk7i6hZn0koA/PXFz79AqTniosA/BuGLiHTkcQCryWIh66hNz7QXeHVu5bD1n+kDShR1KBKw
Y/728XGNKfPjOszlB+DzVEE9wUNx2ndhP3xEi2HicuMrF6rExbx+KnlZLCx6xnxZKigIgY0HoEpx
9pzyY/lzh9i+oNH6ejbTB3b5KotlfRfBtXniKoo+LRCPHbL+25QQgwT9r1Jmi3/vz9z0lgld6Uz3
+1IjjdAlLaSKXN/6j+S3uCXXfuPtKXFnCInFew4TXaT5wwSPP+/FdUi3i5s4IxWgOTC1bDMRVtSU
3K4PgAnC9c8E5FyoqUWW/p/vWiv3kda/5QKMPrO2H3VVngs7PKMo+SNQX7UhhYjOrc0NkBBIkj6n
qrOyhQST2icgp/2qvwMrzZPUtpu5vHOGTG3ROHNpSERBvui8DQBjqpGoHvUcSyDQE8ZwOPyAVH4N
vBRtp+gabFOp1qecU3UI/7vPdmLTf5AtUO0lqpGip/KBz8DZlwbRieZqZyRLsz1nhp5C2fal0ZZn
87ws3t1BftnOqkWSFW9n7ZwVi64wdOLfvdG/2sT9BGF6POQVpQuzHdID5gxn32e2SzM87YFFaAhr
z9ltztj9z2errrEaxH9+SFG0QxNyorH+/wD5dtRow8PSJmyY2PTXdTYXc0umMc1UoJrIYDN8TtpR
NK6ZUGFxNQYB0WHVIw93EbNpsncK6zf95hE8qz/scxYTux74lAoba1CMLA0VNAZClAqhFZsx1EZw
bPzfkgp2Yl4AsQGDGnowV2BKYjDFCGy1cLJ6y2Re5tRyQvuoxWHLVCL2kVgrAbD3q5otGHFbPa7d
H+I9S7RthryfPpn1iX1SGJ9PZFtBzqTl2eGvbdHEIOTaMvT5Osde2TjXl3rSjXpB6gDH7TSfonxT
JOcL/44LQnndzprq69LCgZtOagwk0pL8yaYfvmXRonoYEVL+U8lF/59Z+13JuMj/jxdQqUb0SSZ+
DjhALqswpPiZB38/1ufuXxZ+EH403itriu4Uw5K1lyr3NKfzsOXt+RL7DhiBlV9CotbheQuSOMi+
bYCW+fISasSF+LStLlIUX3zIXJ0JJzZmwms5/EqcNV8i9brTBFi3p8DXXyI/ESzTs1SnL5/Rq5lH
Y8NYPBp9sHpb7IvqrWgISUPMpaQQlfPLuM8ZUtygVRVvw/45u9OEoy92Ju7whvak5CXON59Wb/CN
xJ1nTGHAeg+zoWPQELcjYqx5cdM3PVa7hInF1V1ak47JvRJxwDodlKy4YcC1r4xhlJbzB1aebgsY
B4jNVvrzydOmbismusI4M1kPrwnsZf7XcA0uHxVYM7SDJWcVs1n04Zx5fQ6IGa+GGXS+TEJvxzND
GlUT95OTjdO2ITGYWo/hGwvx0hQlV9wbXiAk29j5irtBQv4O0HjMFXXRNOWMuKXFVbqSgbQjrw6A
Zb0V12ACGR1pevi09q36ArFZLzNX3g34ELFhA1T8VdyyOU48+EoaBV8hOHFMbCtYHp+NWYn0XlEd
UHoYbtzYVSOUEEs8q9JKXOWLVSfRlcFLhSjz7aBkibiXTDmwgjJfB/mljxBbpl2OKz/jqg9MOwQX
bEpbBmQ1W5RVqq40eLehv+8rDnppRAG081hTPTCZxRYE0f+HGkjc77WZ8zg3TW4lEWZqhbAhG8yL
9D+D0U8mKqwuGa9beVzgiWYK46mW9fxY+inS8Zqt4HG5i5PkicGjCo6WcwLLvx75u/CDBe7XZmkE
Yo4Xdig5rJyczzeOlUDEjE7dlZ1NA4W3oaROTKVWWnMa00sF8aw7HQ8KFcUcywYiSLb7xAsYjIhB
RA0tz58aVia7c9F5Ee4lN+9gV+ZBNyA8B+C9nsB+WOUr5tD1mMzit1FwvbtgzV3wIME5kwMFwQ9x
U6fiMCxMRb/2My9pAuW5aZANyYCK/y+vlbh5BuXUX9QvCHYL57C9ALLgNaFYz1lgCZY/R20Egr9A
sTh9K54aFMZshyrMrBNak91ec1aCx3jtHFgVfeWyh9yJAq1ZgKpVPES2+EBvp3YzLbABsxgyUchL
dwKlMzXsOtP2xqVvx3bZzN/Q0LSgKdYnuAW4fPA4zJA4q7F851JiqvmRrsXMhgAl1lWPooC+4Vlm
AT7C4/lac97dUZVJJAekyRKiuene5IPUkkiyi4I3w7V5LvD/8XRu7uv47sthUXoWhAsgrGqP4AhY
LwS85RKl3xzPyzHglDqyPEsyeEWj8ZywiGDouAd8xitwaJnNdyJ/P1aGoY211eZ5NGDr35JpeGZV
m9esE/mt5d5YHi3gcjfSR4MAzNqoa0UgROnBNcrIUkW2zgcK2Vldfc4h/tINmg1m4cOH7bJL+mua
pxC7Q3ddle9l9YNun1Xxv4B6GNRWFZKTl+Lfd2vX4fCVwLCbILzcTeg2hsbyy1LOrcedUDAecW40
eMXYM72tPpcVIDVit37cONjDzrh+g0cr4tC90YO8AE6GIFa/jzMYQx1jnkAt6H4J13xKzbsbQVVq
bJJ8Qw3G5COz55LV/TFPVjZczGFZ8oTFDjcdJ4EhP+ZilzIH64I+bhsrUKWTM+Voj+KkWdYIMK6j
ErooqDeyQeB1cOyvKehw6SHt7cNozsWIAcf9Sy92ywRMGPFyuXz5GJ7P8U95dDPR6+TAOQneLAMQ
sWit4BQLSn8Hk3FoFGG4SJ5xh1TMfKrXLI2IoHojipAEi3ljdI181rKiQZ80yIqPv8F91RH7ZXAJ
4iDZpyWrANj+Ah6HcrnD2xsFENHZcAIvOVoOnUNJ/tk1Y4qqDs/U1Vv+nH50mXr6ec9Rkzi665n+
IZ1oeb+jRT2SCWCmTAaa0wJvKWe4LSTY0vIVWO10wmmu4BLAQ9bcxJotZy/o+gcnb7LJlQE4+g/w
1AqEvjjCdU4EVy5vjf+n7meALjR0GluMuZfzy7tEASbI3Qgo3nlZZIKF+Fe+B/NPomGGd8DR+JVo
Nmh6/JAdjE3MyyNppd8YnFNZF8nE2bbauS5uj2DG5sI5rNz1du5hgT/60xiP37FvMciv72Vs76Sg
lsyxm1z9WCObQ4boPay7UcV8aJGC/KH8bTHxGAQkt2c0odjpprAlVJS3Sa6TKV6HtuOARTIF9lH2
bmxSdv/6DpllXrQx5B8x23E/cIHOH7NkYv1L7C3zN2SQ1tNfNrNWMkhJnkUbFyNI1sRRHhDJJepV
NFdkKyn8TMa0Sb3k4VI17Ei+AVgzT4x9aEHW2ZpoKQzZZdJcsEHAQKGkTQzMgP/HhUuXgucC7Ei9
ByDl6QgQd5mj7reSFiG3purOdH2NKrM+ie8SVUR7LnyI/OP+yI1e44deTgsmmQITBm3Xa1HhBwL9
5gIItaEeKe7irPyXSbgLgeB7GIAJs/RYMETLF9bo0JphRy8oDfC8e6MCbIX+H1By0/NYY+IK5bi5
E9/xSg0IHCWm7TALGi1f9VdGR/lrbP+GyLei/yPk2I8SovBLHI7QptyZcvk0gkG0idLiLvck0RAv
3pjbZZAfKyR09Mt1n5D2agSwBHK0EI6/Ao9/riwfKSCOd5HdohpsZwJon8Hclk+0PmKYGjDC5fqk
XKRd1pezD/RhKrJ6NsvAiuCaYVU+7gwvspGHfJXPhoDVYlxCNiDQqFYa4IulsgkVWT7OjRqVY5xG
PskhhyAHbZrHsUF58uLQZt+m8qmvuXvkR2qAjlYk7Gbu26p/sLbD7TKbYuhH10xzx4c6x4RcLv/C
ZvPv8F1NUqt3ppKb4j8BF1jyJuWNfvy/92BK5ZtK9DVyoxt5JnV1ur3n9THOLMCFj3Fso74YgvTy
1bm4/TFpwoV9SzU2UM6negio0+KO/9T9K55JmH5zHO78rcRET4VuQUTUIXSeI9w+K0c/DLo9XyWj
G7WOW1zwd/67p53vekCD0FilIAmRWGBzgKIPLj6oull7UulyV+RgX2b7s/9TJ2G9MmjPqGK4bK7j
qgh0C0taK/plToJZys8OwbeC6ijF2oqAuFZ3Ugs3B8iYaoxvsIj3rIxveQtXtfG+dCdmOYlATg4P
ITiB5kY9x/Hjimj9Z2rYC2wuIz3el6T9HWialMtzlsfSUk1peudOOXHzLI5HZKUGe+AD6+zHIaEd
QFelD1csCer5dHoVa24TZpmtSYbjxDnc2yJZXLCMwneFe9yqE3lOegbiwkMTo4U42/FULme8toFg
f0rDPMqz9XvDF5yHq6JwLvl3TLPmUz+THn26fY2RL5cG9/K9Ba62hq+uf5r7t75nQYKI4jEUC+Gf
EhMDXwVLAtzH4TOBYu+h75pesmr9NFnI2x1cO56ag+zptuURQV748ATKxqEvJeIJZUK+geeN1F2H
CDZoZB3NOS9B3YiBCGIqOLnUI7JsrjsuHTGRpa7XQ33hiOkKvcynBnPUwdUUuTN6mVWEZdc+uNfr
Yam+L+nTbjIXC4fGFhEC+FOOCcnP989C0C6SIvDapvCWsUXFa3k1xAtA3mDmzFLTbEiBdHwrvDuJ
N0bDrEtZXbatRErpscoAv38jib8zY2oc4MMdL9xlOCOzibIkj1c1DwCr5JilKIxRi9LkVx9aPOOe
W4zzbKqAtdikY6VvLsWWxMXmEmJfnZaSz+m7C8ScIHsNfNVMOhzw0ExGiociuQLCoH5jnd47Xsi7
wIYvlwXE7OdLrOJ+DI/Fm1uuRc5UTnXqoHQC9oWcKbPvdBa8ChM7l9noblmGvv2pFPfAnY/wXk0C
4vYGJzYCN66VRWHvR4MFMMlpanfXqUvtXIRwMVAIegrTAgi1r6OiCSTtVjYlHN4wY/eT1M8gO/Gf
9QoQ//9RJVp4pBHuUAMU7PD1DVz+JhU4oCmlvdakvv3yc6E76O0lQkKvIoSioij8SdRw+IcdjjCR
HQYKLVrsyzfs54DoYiqFYtiqLtup+ugG4r34lzXcr+SaOFCcyc7Wxv+YMC8eie+r8qyy7s9QhYWd
78j0jfMnn6iExjNNVs0FHQVFJYigY5yy6zsTYUVNmvpBl5DAJQ2GZk8sJWF3oIiGbZoMir+dVQQJ
SCaRkDls9edZ2yHnqP4eG8kiEXu8ZJu7wy8RzlLxQTytGGqin9FMh9JwA2x37MpobZehm10JCrIH
TKeAb4fu+USare49A3uOUZZ8YF/rjnc4s8/yTUOkfZm5LVFjiE/WD11KfBU1VRUGJ+q6ZPSNUhXA
CIoJu4v7/w7m4MG2VB+jwUiJ6JJ/CIyiPqM7Il3WbF9eY+x2th7BWfWzoXXlfnXkA1VbxO9kR5Qf
yQOe1XSS4MVExkkDHOOaGSAGNUwmAGcYgt84UdLHSpLJFZFpB8Y9h1BB8HPrfGScQhaN31Q+Qqam
7o1cSNILe0QOJOZl/C3TtPoepcHK7+9G3q4DFeJXTvLkETuK2fgAEK3N748h1Yy3j1kTBJiB9bug
IyZGms1ayanMGKh/wvhxvXP8aI3dSY418o2jFn2WBnG3f51kP25qtXcI3Y9UOpDpiNbw4ckdNg2q
WbjKQZen0Cejm7iDlZf80nC+QVkitzNEFvDAAOxUQEqi4qUzyqlHWSEDcxRtKGxAWAYtsIF3xPAs
0zhSaU1ZMogPLp0Kz6G8OUWCLSnzc2fNS482gEph8kRwJ7G8/vVnl4Y2SqFZvuAcen1MUjEUjl5t
edahSasBrIX1VsEvzsdhgyaqJiHm+2ucupuTTeoYF7Wu1R6Aa9rUKROfKo1t/9+1cHYTgwTTIpkS
tbUAXl8kGPdTsDgXTY4ksUXKgxf9yqOZ8nb3Dv9n69u9X8dX1+Zb7f27G1C+TDpG9QYLUC4+zaN2
NrgLde0Z6fARiuRRIAsi8prghkajjFhM7yEZCkGqYDvm8pClv14Nw1r1Ac1L3ONuih0Egqoa5q4d
oVrEwbbD9j9x3tWzLF1x67sjdeMqJtt49us2gKxLUW/rB6Z4F0vk6hi2F2pXeU+kUVq1E6UA4ckl
DOz8/F1OVC3abEdDdCoQwjegZsklZXiySEo8gmJ7VCXgQtImOZllNMqIhGpoEy8RvwbZGa3L72gH
o/ww0XKJqR/BbcHcxNMcfYmuQTi1pwycCcsjp3xEKxBX36x6NRrC/SqZ98VUW+wM96GfmEHr3zey
gGEA+JG7U5CxJPgwBznxr6UUNpGuhmqfrMG2n+OclfjCIMUWM0FodzeuTTpmgZm6g6Dt8Z7zYSAw
pO5adIV3mdR80m1ZyVwo8WIup5pmBd3o8aaRVijgIfUNUZsklHJvQBlUesu63bqjDTiAaJ+GO5jB
0jOcJElle4FOWhxrrUKazIPbLQ4EjPLKJfRtBYIkoOAGA0g78z/CZIFvXCCKc5uRlF2LfbBNl2Az
Q+k/w036d5AjsPqWzHxDmiTWrtC9tGOCDuuSVDij6fsGbxnHHD/iezibfuglbgIYBGMGA3OByNbA
27Z8NRpI1Ajw/dS2Lg7UC+MgA1TxHSLIObAZLyk3SnegFXXRUuByabq9KKnc5QwDnxOXTY0v1eSA
Zadt6MY5dYN/twoPzGISWJICndvXn2sBIMe5quiuU6s8KkP3tbOi6+ZLAbEMJM50FUaefQrA+zzy
PK2ypeUQxhS2Cdw00krpV7WUouXXYiCD1Q29luphJ76UGJfzR9RXa3kvRfJLC0LaMG3n0oEg6iaJ
3nWx5ILulntl51IHx1ekGOfiyYFOQCxEbHpUEvypJFKcE16sryAs5gTtpguhTUePCJqlG1eUHvfL
LE8k9pX9BuK49udjVEBkbpuJ8YVsgqIqhulucIDI0jHiblOqeTUIdeY7GR26REL2cL8cQXWn74Vr
jSbxpK/mPBdwkHdTcSMExSYbXKXzpemIEpajbJWJ4his00I+bsg4fHaKSOch2ZZH09LkQ4HHi6h2
hkjjgrJR1oXykOtC2gjQyAHQqIhIjuaapJhgr6b8E1ZX+wSK0jPasYkACsE1EaAi9XDYFaVmBco/
rpJUC9CAmlmsX4MfpqtvRIkFUcCTkrQ1rz6spACF1lVperQwBwg8x7ynyChQexy9jLKz+kXG/IGW
A1qwF96g9GxIqVRd6J/qo3QG5BeZfnWxaq9cUXotUMCNQN+ZB5PjZu6WE90uvwbSzCKeUYRDkKlW
29OghreCT1a+d8fEYpaAPKqbRw6TD7EHUi0kTsJa1jz6R2g3hUgZvslx4fIAPzBjZYGmTx4FZxMm
7thpO8FbNat3KptANmUMgbiu/YdBX3lnZQtiFmCTWkJjHe09TroP1YoLAW29cjI62XSoTvSvMORu
qZDyVCBB61iavFm1n1cLEDppA303bvcwm4QS8QdVtoHTZNnnJMgPB7ftxPX/8slbAzqroweEuIED
abCboh5Zg6qe4uyKtuqyZSCZ0DyAhF4O2yXIAePJsCaIwpmUBGm0gF34jLDCDR67gsqDA6R8mjiM
OF6I7joQYgip7TTUa0eWP6f6N9Dv8FR1sorDJV3B2FrbHl5YBqkImR53a8ku9Mv309Z5k4ze3xZQ
Nm8pzjs4uKSNn0iIlHARwHmlWOPngASpr8wl+7Z7D22rXcgjSeO2Rpe14TFytsG4Fqy1WVVdJQOn
zp4GHgBwVtom8HOL8ouEWb6+Rjy/lajoBD3vyOsx17Js/yHEPIcaSuyfJaTroLXd9HUbjc4jgZb7
lXsbtJB2DYas+Li03vs+IA7B+pC+Hr0xc7l3fnmN9PI/A/CrKvUdKtawiDUYHmVSRz1rXFAM98jA
K9M8L7ctBftC5TkCgGE9vcXDMuay7yLXIGo5pKbnkdghZO3D6WInMRYUOab426hfzEyJxdNIk2xt
TD+Kls2pq5Y7FY+yvIIBoyjhkt0ALrXIcwgq7urSh+nLWjbqeLBfi8YHvOyNeGW3+FH/dqByNIXM
pNiQ0sY7a38PPY0TdfaSXZgOSccDYtKSHRNxuLca4p1eHvX8at84AS6xMlPsNon9kOhHhSOlYxfj
0ZyQc8wAhZbhlC4Z0p3qkixU4PE/dSm9UsINJ04N7XkCp//g6aXS8ch3GGWc0AhQYcGZ5PWfRfhq
eNwEfmL1aZdNe4dkrZxVc88vM1CXXpKFNrzNuL12XlPL/oZu/2/2mcRZTk71OPwd0qPhPpgCM4ia
lsJhsNcVgll6tJOQatAGtsKFy8ajOO6YYXYr9yJGuXMirvU713YRIjPU6XkBaUFXI7XtjJJLtxPu
E5TLEU4SUpLxMbZRBRbQoOBFaXkoPGvLHjryKxoDcyxixbynZWI3Bq6lvmHyZq6OUiFgezNcEyXx
zCxSWczfBZHLT+xDHmTzTGdF9GsUl9sJLWzYIrx4dCK0NxvSNJErm3UYU/js2YO0VDyPO73AL1/k
uW8eG1SEUiNfaENIyPKGyzJ73qCJmgh/GBgStdOYfMHmjcSqXIihWZGRZbRlqpcZxo9SxI0yqHby
B9fKO94QnCoH/3BtN3vU7MI0yABxbNJ4FtuMx+fuuI0tSEn9f7lHIFdvEzVYYcAUmW32w/YpMip8
CSD2HW7UkeNoZ3EpV57MRyjRCFghBr3jaGDa93iHOZxyRl+A2RsTyxOogX0Y3exnRJaZEhwFYcTs
6jMVzSt0yrfCPvI4zmdgmJ6DKfNq7USSbF029prd9T06zbWBffa3JTKWb+76cyLXoXIH1SoiVj8I
HmmetHna0vqKi3rCTwdBW2mKk0PGIQf0BZAIxB0XTCXD154a9Rv4b+M08SeFQtOHKBhSu6uEMzb/
4JmXF8s8EaJMzWfZXQ/OIeFpGjcT6Lqi9KVhAzj6ypSu98QSE2Tb7cSAQ7QBKAQ1xjW/Y3s8le63
ljCMeHRkh5m784AgZpo6Z662o4jWOqyXKKdzUWo7PYPPXiL+P70+fSOv7t6qZvWJlc9nFB063gDN
YDSYTDTPeTf4orjUOCUjQY/8QtebYbnAumgivFvneql4+a+bs7Ty1pN28voshlr1k6hVXTJCWsoc
r5Qb770Rnd10+lg+/aM+Air63O6GTMCERxUlp5cekRKqUPlPCYTJSXqJ2cZfY1psfR/jdgBeFET5
zyTtTalBkRUbFIVDn7FV7epJctmNlfaEvJX2YbTzUNNl8Sf6s7Rbs4fOwBNTYH6lMzRkzNUjKj9y
395r02Tia3SRoyEhnkGmctpVvy5/p8OEtDUfbZdWekGZDGjtSD/vu6KAojru5pgrw6pKck5Q+TfA
rVconxsgaBJg/eUQtiFE8njrR4YoCr+XZ6n4EBVVh5UL9Z8UBlZkJhAo3AdwM/Y5nQI7w5A+RXOF
QpwkSM2JXRwsXHwmMXSCvUEZY4dg4ogE3EIRrBfiUZ48W14F/SLdJFHbLvw0WuBD03kPnZwMbl2q
wsuPm8zZCUlqDglG38IKdIeuCFO/lkGJGuXFZvYaRflDzxi3ARGtmUugzqG2XgnmgskGMak4Yw9S
sqoTqTQo1buqxBL5BNedbZCyrVi12rl6nq0MP02N/58VtTmxtbC2rli/jfxaalrZzvZqr3VzwQ10
r8T/+L/eZ2FSSWTW7zJVN7852VQ3YLvmzs2uQHr9tukWPxo7Kh9qDg11PRp6nrt+U6amYS/kLroW
7bvgxfvm57LlVz+Noi8XfZ4MXb09riI9J4SFKu7LuL15SHQrfUQf04S/f8Lya+uOmriIEWe9C6Lr
NGRFRom1HvYWCFwvQwfsvhNjXPGPWu9d00D7tpY3TkLdN4zG1OdS7C67Q3A2iUqcEHZ/vbBIyy+g
PmBwLzyoge9mXJKt4FQUaWnnDq4mis338vc1nis15/UFy0kW/rhNl1WYKYB0xBB6DViyv6aXYVTv
vElRM9QdxldHMgHiGgsNV+uxtmHYnsIikdUJsxs+OWGhuaQa+FPPN5itExkF7nwXMGXL2HYh9Rhq
N9sMo/chOdmIFQvHKC/+Fk+NwEcuxeo7V0ZCfgmPmhrb5wEbAZEievXU+kLVVqRVE5bGrFJIf7ui
Jx+GynEwSlRAmotgPzDZM+PgTb5qB4VkavvQ9t8taaKQTKrAthBkAWeNvPuiqQBej2lVo86RZMVB
MoSowV1YhTdX6hqgcJHBR+29EloyKfq2dttPx7+c+Ev5zVgf6gs/IvuagKwt+aEevEPggw4YYSUw
JBZSfK4yx+8WGEh05QYG8ppk1ntcmGrmQLIIlwHUS08inLXKqr2bZttsj/b2AzeJJmHoGyBMuAFz
KGdFZFRRDZtVyiWCRUGfxp0DHQCzFrrItcFhihc4VhCOnFQ0BCznqaH3EGf9e4VgcHl9KaOwS4XS
5wI9lKGKXlIWG3wRaglopqsP0V1aPYhuEVnYhAU+0ZRpI76wi1u2Dc1tSAAhY2OvQVABZWIYe1AO
mcQS2m3kfbG3UDy4KTVkwtcpr9OQ7DxgUTKMpecUIICFpRnmej3zw6IJKwxj7igq1ujL/q8U7K/a
7ZU78ty9MNS80N1PP2n83J4zbnbgxNLTNHOsneVte+1hQ0PGYM7mboCMqR3Le6D5KwnYGYITyM0U
J1q1fd+TdoV1PQr5LlLEg+EEs+UcENkCXvmpdBExG0QYUSDWQt1c+oWdUc3URgWCpMeuUUD6Gowf
eYkEz6Jttai6UYn7bWts7jFAJ00yLHP6qYamGUMP097QCMyHvejrLGS/7MN1eOTIcyZgR+N62HIU
bWnIb2qJYhiDc+oKyT6x3e1RB6S1M3vFgOfT5yOEHz0riYa8ogEtZEGsKYdCwlkECVPoLp+yUhMR
oCFQMOd5VYqk6fBbhbJxKu8ZHTBNR16mFH/lOy/wNUwOONTn30M1C5WfzCeOQcD6p0WO48nnWOgq
lvEvcNwjvBKQcxtuaCa+WJ4psfpNf7+JNBM2tcAUOTbQ6G87+1su4OypHWipqmKQiNkXIAUKWT07
ywsl8Jv8DLt2tHW7L+bqLaAK2JOBxBbZ6KKdsveTe7WhVtN2v7cqBh7MtQEWuZKfL/k6cYCC7qwC
XxQQ1yyuTjjx/a1YBB+f0jlNXtjTy7P5V484RmnWWroTB+nT+j69Y4/biNPGMwYEedX7cANJzF1a
q1NZpDNM08z79FqDkL2G2+CqV2A1otu7eZTbp32NpLewTQnY7wSLAhteknxnUGfZ27ry8FImbq5H
Em86PGCUVuaNfBpdIy/4IBBVjnhDm5MbAIb8FSj8x8I4YCubv70uF8b8Sra9FdcLXvVydhDF+HBD
quIDQEObQmwukjup5BA7BBVyHHQCSho2EMx/fF9YXUQm1o/jbOwVV86MzH5Ia0LCQuO/VAB9PQNy
t/m4NAWO0XljZglzevevkEGGn3ldnvA5QBUnw981cX0Yl8Dkmbltd2VO8C61AqFvk639ZsVVow0n
PP0s0JySafLtglVoCkBbNcogFWdd/Ei5GKpIc9gmm75jlK6HI+pEwYCC+f5Ik143XbQQdhQiNtNI
wDbbMH6TMwbVNF3SRUTFprOnSbAFF06+ET7GAG7lxas1CipavM2yyxEMVRodiOMiC1qA+dBrwh9j
WfRzjTw+Rd5h74LGj/5+18JqniyrXez6KqxXtgjov/VvKJZQjwG5kVrGmI5CcrrnScZcIZfbgzN9
VX/9hHs2pM4YsUeZHQGv30pwiThi62Uhe4XOndtrr+yF4i6o0d1hu61Lvxcub1c+aHuMktNPj73+
r5NI7hNQPtYXZQLx4H9EVh3tXra2KLNTWfVi1QqNceJ4EFALM2U+WwJPSutMCAIpQcgdGDrV0oc3
VDoOLPLeuHqJStflP5z/1VWL8yZ+XCeQbL6U5f53ryjxNV1KLag/pfZIa4S2Sy4zcPwH0Aa6um0s
Xz3aYXmfyewbnN3954m0tgXbXaPjPE/EqDrggqmDL+98yiADnZg3MAY+3AqPJot866BSrVz3GZSy
FCGCkQUFk5rmzl/yH7O5iBvOCYtPG9iKT8iHs5pFpWp/jhfg/PnXZ5p+z9sNzBbZ1ugmW/ZphxlD
MRqnp7HwzLAkB6sTIP0gGcEs3zjSxnYBe9StDGgTh/CpCyfYNxq2TEx9RUjKEsImZzMc1/Inh8jv
b+/sNSZ+JPBh+k+P+ep+3kZKEjHRkjDSjN3fTy8u+DyDwAMI/EuWP64Krw+NaClK/6tm8jO0IOf7
X8zkqIuxI1TeBxgauur60WvjXaaY0PPc8fnYcdw7FeCxlfTJoLoVSpbcdpZ5O/a9ycBXi0KgiAoc
sLqnbKZtzV1xHBpcNJA5ydgX8diDDqA0lJxsGYHQolG5rxbdluNq+kdU7qr+hA5dBRCIreMGKBq4
pxAwlnR852eOu5DzwDZk4GALJpPwLOYa1XxseXk1Nlg/2jjX3WlKeoDISZSJ2pSpus7tXUInwpeV
Z4K8gAsNHksu5GwuyVwQxKSdPChaAs+KmYob1JF4BXNgAURLY5+YMu0EZB/fmi7OOhF6nWUB1ktl
Xt+K+aAU2y8yNB4RMOw7aJ7i01tn6D1wWIsR0CnQvMzVLZb4XrrcPF8TPiab3FrCdESrUQrB11vf
/mg99eDGwK0Pq7slQ6jQr+qeFRamyuzoIjFOOyTQiL/HjF2ZRbjcKQhqj7rHPiDhUYVxPlsBNN7f
/CrIL2O3Q77yJkug9vG9zzv4WeovQRLrP06rcOFNeVxmnzdTSvqQDEWvvBhSLAYRG9oDKNppDEqv
UV6EueLDPGA346KDjpmsTMFjSO8wNzscNg90RMT6gVd8gbrJDcJlxFTrI5CQ+PGADRmvOPSCYllE
nJWAxhJv1dSlk4r9VEYceTmchPYelC+FezVZ6D0+ngibzyPJljI97C/HlExaGHZQg5+zRUFLLMx7
fBx92L6ex2hCH3tAzUPAMhsH9TlQy+A1AHiq2Nf6i1fU/U2K1rnkrnIbVTMmQzt6EEheKvBlBMXU
rZiw7KBvFXqMVE6WxP4VaUSQfQO7RFy4kYztDmtkT2KT+gFMv77+DqtmOkotjNiGN6ZpNd97s7cO
pnjw09foPWpb8mzBAvY5vLwhIPFyFEuJxfffg5QFj90exNbcX7uYAZWQshuPaUbJo6t/7aj5XO+D
+00F8YLSN+znDrmYNLL3XBrNhZ/pzOumS9ScokO+5jXWzL2LuCeaQEh6ab2nvC/sJcBsdxtQwT3r
x8V0MPqjf2JpAVCNaSNm9/k0ZAHf/i6ZbzmDiyXjJwA+Kzg/FA2g+M4j70HD30ysdQ164lqrbHCN
XTLz0H/dG5zePRG39Zs8dtL+U2fmmV5Vy+0PkO6vdpHs81nnMjh64pPrEKp58yVxjz55HfLwp6pP
ND0oClnUvScHDxSsPXjkSwpWy/k6W6O7KiXtqpefilPf06I1RFY4Ytk8DNy+pwwWM/VhPHWLVB+W
4C/OmucFNjO0grNr4gQMWpxcyT+/W3J4alGJcZFOiAskC4vIWjlz8rEPBitEU+6Co8ZUFgIw2W1T
1ztvH9+qbU+bisp5hKNfjl/r4/wnbuVeyRIOg/XCKO8y8AZml3UEkZaNs3wlTL8B4eWJQuIPebeq
AvLjUVNd1VIfmnhDuFm09coA8skCTa7EtPcAc77HH/OYvGFThP+YwydReqbmWpMZTRULL0LEsdGs
Wog4OXvG6uIKd4fmAf6msgofz16dF2/+rxD66CozIKEcPP1MhRN82uE/zPle3uzVm/eyNVqwsSoj
9P9GsRdTxJ/Eh9MlmNV8KAvCEy+7l5TdaI7UMz/2fClW8Jyr55apPOjAGnrV9RpKlm1yWdSgp2jU
jOP+sNrzISAs72WIe1EV5LpFBfGnkVuhbXHseszPP2pTElEl0FYddzQAPcv5558ljoxwcL7vJj90
p3ZQdK3isw/kaIzRh53+4NENpco3IezdIj27CfPwaea6OoWZqola9ihdNPh6yKf/FFJJ1U10VuvC
bt2EDZrBF8pcwmZK5lX27yCZhMkauYjMoRQ99dWuFEviI5RV6J5wX09UExL5Lbk3RkooEW4Jiiaa
R3jnpheXd2SHfNsf9wRtDl05SNX1oZKPaeHYIK17/Z/Vi6b+e5pCXrEKcgnj6icECvW351K5uNAS
babsydFAxdHXka6+n/YDyRj0hCypZnRbHCypa71E/rgKW+xHrgVJOex9MERD6PCrUVJ6hJ8ofoTE
3VaRj5Fr7IwbVm3V9XZBWAQ6IIOBKdbH+A+VWpiq0fA2Qokg0TPXto3fuV4ptplyCBq1PEqw+1DJ
/HvzRPGyA//iUODJuU0QsUwYNwk4DbPrSxX3SDIC+Nb1y0B6RLgXgE+mc3OzmXlGYLYrVZR12zkz
mlaQBJo+VV4lkLrh9ylV0+geshDDhRm9XdWOM+aM3SjGLD1jiwIkFRWwD73L3ofGk9iQ9FJfxl+M
oOzdgZotGNg1oEAaiaCSDCMtNrIZ0MHwt3HmWsQJSiyZ6rzIGXssRiKY3qunt6q0Twfb5DSjq59g
tRZS18MZKsGBephFz8DQav4qS9VMwsldTzZ2TLcQ6GrKgunwV8Iw3+i+gKJytyBOQLn1554GnMF9
cvv+w42GQLtROeayFQdVeD9HVNgCgBbzkBLwY62tQ0QJdVv929K9+cK6J3OSTywfgRIWexPF58JK
f/JuyBeaiMO/23KwCioP809EFC/1GPsfWGWxTEAdDtkIuk9OP9DrbUmQ4tykM0ECBKEeWcqG+vsm
KgzMyAbHRqGs1KYpR/FXFVBebUy01Ed8zaJsmplOqwUTOcDTD7oLzCphdcW0pBsAwlfA5PplXH83
O0LGSSFe5utzlG0kbZzRW+rOCg5Vs0oF34WuG46KQnMQgYfnrUZdr24QgefrrAHj1RAYzoiteUEZ
fzrs5XJ3cg7irThgoxbdVD0y0DEa/hmA/2Ntzm2RR6vToVokXJfHpPRe6JhpBwL3rXp3dM2+y2MT
rxBHcyXStcz2E2LRJl6hQcCbJFhqd6o++oEiew0vlB6bOLmhZmZiaKP2VtBI7lJsut+u+LGE81vY
Le4/GViEmf2cCnLiEbKehrSOh+nmXig2h09Exk1/9xgsd94LwDZjZVzw1mIKfnrk6uV7rAfGkygL
wkVK1cKDXQ6rS2WabzmWtM0r5aD6mSRfVS6gG3coDSpvbcVUMykyoi0AeawUzBzzo7NHVnpOk12B
bqzxXduHdVH5Ajf+Uf2M6lwSZcvmtiyrN/i/452JFFHmTiFwYsU/RP9yJwSl25jqqaIw9CvskOM/
xTTK9ZZBWknzggxvSliZOxU/KAsTCEVHAQYMl0q0N5oDlStUj+0OHhC6tTZVYOC+fJWSsn87kdGQ
/HGRNZpvftvg2W/B1Y9g1zJZIdond+1gVZwvqYkWT5PgfT/pBLiiIQfekj47TuL52yKLoTMLnbCY
klA/jbPLXSlOs+FsZ2fHJEQRG2eSBKoUcnxEIWyDHUoq0CRzCFPm0wrSdP4RtbdPwmFK9Mb6PLHw
2huAyM/D6Ftytue7JGCYQH8w+UTMDJodelWB/XJcW193YYpGvzZA+R0bs9YuxYx3qdq/ha6cItDU
MT9wcCPO/GVEXCozgNDbkfFRC1nGvbx+jIo2Mto1Z/9F/p92hvV+7OeFNbQ65JlQttPsD0nR1frJ
rdjfU+EpVmlJTsLzPsEpPxxEWHlX7Vo+/tAstVzp3Vq+VB5ZbiTSp7LIcl1Vt/oaUJYBCCiQNfbo
C46rrjCqG+KaqzRIKg5Ftj5seoZoHNKEUIUjGYO734B6JHN8zBPDeJYycSdzezLRL95SgQyRJ3eA
S65JZx5uD8SbkWXsT5nOdKbhv9NNEYaot9VQY16KTpYtqeHrICU4FXGue0WXuN5ecPdE6OIZ1O9g
H8+EuAt0vE/Q+P/mgN2M7/JzLFwmN52uNLT2FmUXlFir0VRAEty46kfFHWLTiPPtvWh3Jb5RID1B
T3AyuKsqzcDntUXQnAs9Mdaq1AZh8vrLjTDJRXFqbWb5objFZo0Y8gBbG89XU5oUkuLfY60g+A2H
tykw+vLKMmQh6F+v4yxNQNisRqT/2FV96rf3e4JwzSwKgGiYA1HkMLXJe1hCM8w+DxoZUZo5fDia
G40ERl1fL0bGn6sevyCbU1b3qMZa4AoyYws7PLj/quixOhWENjnRLAcRuf19lSX6Qb5b4fHDPGzD
9k4OXIWTn1aH79Da4QbgPmgx034F/yy+fSaf2tQhnJTPKtTPaqr0MaKDmUu6pKNziNI1hLlHB2YW
qVYTC6Wk4IkQcQYR9qtJF1AWfLgNVO/mN2vt2SfKp0GWAmyXpOugfCREsSlxaKbAfGnDL7kXZkG+
g8LuptJQUzWa49uKDQWWxDbg7oeuhsSLz8Vcd7l/S1mRJCKe88HuuRCrhYnVBE/E1D6bIV8Co9va
S+PB8RjmB2XlZGcFq2nuXkgQRqR6vl42tbcenWUIZmUTwm7NtY4FgLOexgj2qli0GrSpFt4S3KCc
QqKhhc7MMjiKhLCyj4FLbiCrJUSp5ixErTOlQqsVwlVe9SobItkDTSwcd/TmJP/4KsTC5N8sAM09
ZBJeEk65Vw1KJIB5uwSbX8t0LCXmQwqOK/fVI/jx55iSE5HC76vnj/g+bcgtJeYNR4KGd9Cb3Dbb
9NR2dntV/ZT2UXDc7tBsgSiYTvOb43RN9+zxlH38v+OXZ27WHFDdz/izYapV50wTlBVdrtWMAOux
8NuwPxSOrWhuYX8Cu1ssCuWQbrDe9sXOWdH0uY1dAGF51vbapq/u0VkyCtINTYCeJ0HROaEC8z8x
SisIacTB/J9Fn/fJhgdadPuwleqqQuyToEna6s1NcHrg313LksXhCs53eHIV22eiPp3KtK/bdVRd
AE6EWRtgfIstDxDa6TftjP555UX6mtI9MYpmUWRG8C0F2EbuftNYvxzpXahV78jc6xt7Wy8tLEf7
sO0uwWim9Z3vp/uWMy6Xosb88XMAy7DjflDXISOLWoDYctzcIf5xoX+/q+iYqFoFutYj0Wa1rLh9
SoyngVVun1ES9uFQ/HtaIj3O2mAjxsE2E//6zygjgJRCgPDP0kHBPCH9xI3mgeJxUW5YHaYgIC2v
UC8CRwZwGDju8vXRMJILIxCEd9GkZWZJ35D+HeZJ+rSZbMBbW7RYSPBg7UkX/WMyhWVIDLLQdyGe
f7LidU3dq+/5W0z6N2wWHI80o7+WoLsx72+FaU/KSrMLDhwaPsi8udGOOarX/+oJGs50IAARKD+B
cvI0p5qW56XE2Kv+6WzrN2rKny4aS4Mi4N+RuFQl1TgRH5hHL6HQf9gddduI2dm7lBH9J99z2Vwq
kq1KuxY5YQ5jxa9I9HBRjajI2UybtPJWEzW3KiQKNlfUPsjTNDGrXD++av1bev96nty3aEK41xO0
/1Nvbzh3lse5VxHGNQBgPY5PP2LOVZcYDg5VEKgMXpISCLxn82fr79ZVNRC+t1zZTlfkgqJ8PfUb
wVTZT4a72fkKHDr3Gw/dJwPmS+C5wWKgcKqCi29ungAvCU6c1SN//F4EGo7eJOgf8+I7rPmuH2rM
iUgMgXNUgx9JamPJLapdgRLrBk22/9ymRMfzqt3WAruGgl+Ysl4IU/cVqN/q3C26snJ8JSURF2dY
HPeGTAT2OVocluWL42oFUzLbfd9Oj3XdqxjsTPg4nR6ZYZorEKCk4nb+NBjgpAN4KvcjPxE/OfnM
In+SXg2N8b33E4O+vmhcajEcSSU/Kl17bAABZGJB9Y5SUhIiTaP37bbSuE1t7DMzmqoCAlYYR5I2
nLBqJawLSS2mPXVtgN1okQZkm+iijfBeF0e+8Y72TvNrvs2POT6veOzXigt4ul9Am4mBgdB/2hPO
a/tSne+hBv6NcCi+JfDjLQnENvzXbcgKnUtcNiobIfdbRV64AhTjMOaEvbqA/qot84RxD6yvwuuK
vVEOIKtfnkRapBMNgxl+rpa6WrnCbVulIZYlU8yKsQhrTfEMmOY+ooAO8H67ToqEUYPtC81y/ciD
1PSUWukovNhI1JZAaU8YswemGjv4+pDUZmkF/oZ6mW6dtg/sGYbpFkzcaq2ihmuEGHhv0/F1H5G5
DwqdGvSV8/Dt6C4DNonWDvxms2UZQRuNiumBJVKE8NgNCCsSiZpfRi+i4c0VleBnuowMgkLg4Do5
wBL7i/YouZ6kLnIb7gbPDrWRZ1FFYGSiUJO48uXVVgfKJYZMqWO8Tdcg1S9uYsWP9zUDzDiun/xc
xmB8+ld+cEURYLDdKlrO/zZzFyezF4oJ9NYkhIGuf3epF0AuiXZFkOopIByu8kvRyn7Ci6WPC29Z
gNSdaZqC23Anbo8c7MY2JUTiJNogsFv9ML+tAOZvbScSBDRRuM0rKWCJDWPfw1JCmlOqlSyD7NtR
zQEpTo1tkc/qJ0hOiVcZJPs7tVDwZ2Eq4wYqbaAah+ohlS3VaHXu6c82iVa7ygYT+H0/m62BujhZ
oZYfGtvAdLShTp/GOeVVD5Wb6dGJkRszGZmaL5XJ5vqvK/PoMTrpyNS44ZnzuC2wRz2kq8NOFsfc
WyV7LsYhyg9CeOK3R34foMzhfd93GoKE+42qyyz8xbz3nsdNIIQhcUB94FFBZ9yXxLPyMlhkPiJl
OHpnBZ96+42WDmC9RrFGsLZMzKEw5L2FDXNcATcRTMrFeDsdrvvSG4N3sYoSGdu20wWSFacfP85N
KsESufZYLw9gRAZeKAxrrlwWUYwHvpE0ZODqu0NJ4VRsV+36m3Rge/WyyRxFPt1kN0ZNfGW9g6oE
tzHugcZguQ83hI6CvHCDAvWMsHtpQvDRUKJtLXsOgngJm1hsTwQv58jibmLj2wx6zUlR22y4e3rX
OftX4bJefwBBv48ZoPHkPetRWet0ARYsvLrczd7pQe2krqLU9v0kJ493akbw8HNJbqIyObUbXY97
+I0xjLLJ6bKKHEwrkhIHeOQWshzFXMbK2Ptf1mrPR8tk7+z28dl7XJcb11YrSavTJiYJ0Dde7gA7
a5u6A2HTIk+YhnrvOLGMY7VFHNgfAqlr2vWywbDPUy6ZFnTpu1CD3pFt2iC1p/CrOPC8xR2x9jnz
ATc1xdonVyEqDQaXjB0bGyMcWlAZBbTuj7V70ehzU9AWC8/UB6JOvcJaHnS/lLLIArf66CbGc8aj
29q3opb1gywMRt1DNc+34FbgSFZCQ/IlqUfMY1/RqVNkVLdzOuxla2LRu9bx6XM0S3ojdBecf3o3
nuorj8BQ/OxUU6MG0L77g26PWRNk/7lYal+I7q6Vil0NWerBhxmZ85mKatWLDhlm4Mpw7J6TDHvm
QZCh2G9YNr/x4svNWBLWTE3Za5P+yqEV7ueiZtHXqUuxmUQJ1wzv4juDdjN7YTA1ZNBhY0ctJORu
tAe+db1CwsNmEf+iYZaYnFTcnps7DUPDXiiKZrMdkavUTdgFlGraZ84nQ7rJtASlqjqQ6ONUARX4
4IC0W25b2K3W5GfBR9GHqJYrqv+7gZ5D3WLj1wiZz280VeSXlrKjdOcoAD91r7yMxTowX56DrBnU
+M8BOVDY29J6VCSRg8DnmOu04Cx2/WAsM+lkQf6jqBD0AQ5yyKboyVQTm4aBpxCZhBG55op9A2Cv
Uv06GkL2XcCqsXfJo63NFCXru+gctkC0nC+Y/h3Id8FiogMVvdjxFA03jB7GY8n+poVU1rcAzVrr
rsFMU45dkLQESLITTNoKZxk620SSLV2eVY90D5ltv/hvovZLBacEXs1osyEGfF1hyFmh6KRbGAEA
zK9RC4SpFEdAHmCkf+08HEjFVceTtrrK9nuQA8EnQgQWE7CDpPqqNdHIyk0vWw1xBl/xM1FFhjeV
BgrjVOSlqoR9/qlncrVeMkcMaHntaHG6rRsV2cv7eMDaTVUxovBcgS05UoQzp6nmq+i9Pe7EA06z
RM4NklYsUv36OS/hg+duohrjcEAPKTxZoziUNZn8JiaMt5ZCsvq2Lm4e231RdZ6AeIskqDi7D/92
+vw8e1v1SY+XIq9nzZKEP1lz6aRAHjWeh5a5BfG0BLVc/XCE48+GMmrBD5+Tlrx+5DvCAOcoR88N
j0ClEuuXEKIn8HLt9lbJtQ5I79W4vcyw6iEypjc5d69RJUlgZiWhRSxOFc9AEnfV2QgAIDJDuiEH
VSHHuxbBj+1fAeAKNVRhZc9BHKtC9Ob7mdenUbUC55QcOIE/jCmplWXrFPD/noRnkmhciFYlcv7A
aKdROvueTlpI/twwzjrg8o/ruzkfZMuwLMRu/ItIrdJupSfzbmYtDi3jy1bjYr5BSGwk1kgqXHh2
qSf7fqxreZQ5rC1AKOgd2YVRVKIciFGp9xYb2XZeXENWqKItWGzDpKrwNT8XhepRaFvoQo7OgGBC
hTpdiLmzuUF/HbhD9/qiPSVrkEYBjDxmAChAK7oU6Irw2HLvsWjsLHp2Er38zHgrVPU54szJTEQt
fDiEB3b+jz6lxb4eR6LqnzmCJrpDA5eDeML5XSbH3/E9MppWvrwYZJR+OIZVm084u1ZMZYaR9op/
jwkpt8xzN2NWJbNttDMC4LTGDhEmaiWp1mub00T+uRfg89MU8VP6eY5d3eXynKNM65KVxa/3d5k8
WG3lb0QmJRAEpiJD69kbIPhDhrdtagjVSD1ylcn/T+k4R4W+ty62Ej6pthFeHD2+RnOwOT8OUw0s
z6JzMfMvEQV7EItEFaJVexIkJLauk32oiDGSEPx2H2IBKxuKS/dxhlDYjAsJkiVPGsUTV2UowqFg
IqyGPhHquYczdCTpCll7T/g921ONGsLYTNQzLFnZwvJ898K3V4jD+5Mf08zxsvPfOVlAPTox7aE7
4WCTqVnthE8i2BWWjSZ2pHLqHYmUucH09iNJ1ojlhRhNkc5s5tRMqawOFrg91zompn0ZttoMMJZS
vo0BszwrMf0RaVU8cROue9MV1KoRedPud8gyIuWb7afqoZOF1stGsQx78Vn9GDvgLE+plvh0bl6y
A/55KYqY84+Khq8iWMLm3O9c+VaPf1Yc0NyiyweflS/l4FUKJch7pX3FNp/1cxkd/154XD2gYbRV
qrn3AbXCwo46TZDPtbzzBAetstlOqrIccdFHdo1c8Vklrfji+3V84kFe5ekPSsByZNv7IqbGHz9Y
LRs2jbpSaKTrITEnpyHpbCO8l+qYjEF7O3mehtZkkCE9rNcnazMjMJ+Cm1F9VQHKPAiQnaImchH4
yPoFUIQbTUNfIWdy819jj0buQUp5XIB5p4uAEoguKes7dcrvfkO7j561JLgyxkALvwRmvWX+xrzU
hjdG8wGK3R5tNdZsIFieyFtAAOHBFJ/CJHwAY8G+W+W+ynGxe+AT4+XEtLUoXZuBm6aywgOScilA
D68aNs1XGsApWGT/IZKzSromCuuoef3cUq9i41TKCEi1DGQrsBhxll0R/oOk/vsOsIkkhKvrY7Vu
1NtIFOi4qD9En4N3GlMSz2BfyM2+e9CbovyfhDGxDf2ZV7xavz8J0FgJcL6t/PFepEr7uKei1TZp
QgQgeH/NDB6iqmN4nC2iA3m2oIH/2pGbSIrqgsM8rgwP32YQsEL65FQXEEQDMropOxgZwTnXyGSj
3D5crZ29u6eradiuOehHqruBHSW7XRyZiaE2KWvUYF44pr2nvB6TFibffw19rv9oTA5H63DMw0Ta
HL6Jdo/Ck8MiPpv81vruW+xvLB7CGUHjm3E7GmOE3CYapc3mhtEoncolzfJJwbntcN4Ti1gnvsmE
3yO6ce3RZDS/x1137WrwTlydbIETKFlffrKyuIMG6Ft0okJLFdDUV2T4IgVmh504N9P2/3cl6qAS
MnzrghhKdbSS9eVnmKu1QA7uNbD/6S7qhB+oD67gYc7kmwhQt3yxKslvQ5zVBCjjiVKioejDi7mo
ng9Lm8DySktbn6ggHS3Hs+vi7+0sed12jqIbxbQn2pAKWwnBa6joow3wEoBTHKoOiJqku7mdsHT/
9+H29pPIzBETJ2AmmjNxHBymuGWtU8GzufbB8qe/9+sAZCH5216rn3fCcHE72xhabh3OUn2dLksB
dECrDMMwG4XEuEr/quawhLW4fxLu3GYquZuAonwp61Pc9rCE4W1V6qsR0PrS7e/i4q0VuxeIcCE9
ToEQ50FRNhdXbYtNucTHt96o4zEsBRWuHk9plDhOX4qhhQZ2+l1fWBys9b6ozDkBcnT38VPWwXRY
SmzjQAG9N1YP7du1hvAMOxIf7ZMi3AX85WkPoNuiPSPHNVe+K051pBihIOe6P5fg3HmW2yiob3rV
hWemMFkvIKVNjVXEKeXkDTPfm2omTRK44gJpdXdPb2zk93tK1GB4D0yegC5PPfA6YQi0Rw2pG1d9
EkBIW70VUKJLbMIEV5w06Qi7Aw6u5l6ho23EAHpcj5lHzN8p05HuLJiWWZTnyg6DA/6AFzJgQ5l3
0vLSsyDqrCqV9YJRvPqpz5VpbxDTG9EpzpfDkExZZu52lV9VGU1lwx4Za7fKQfMBhhUluvYL0R3L
Utbkt3IZGy/xXJnelfjVeayQEw+ht3kiZltsWGXxO24aprqktjj1/3OhHQfk7Op+71ljnDqUYWfm
oQFXR9qWEultVMMlzPb+G/B21HWGrCFCM3j5I97zuIk0eC9nnPWkZL5DM9zG+qIadQV2EDrHLEPz
4SwvJQ+XO3eNuedsNdmENkg0dmPQzfocJCBJO1Xo9bgj/MDYgm8u0zYnJPYtFP6oWiqJGUzAQlZu
X1RFRg5w0YHhiKRijtTWLWpROwojJ3q0/Qk0nFgdCFWcevJRMV9O53WkiNDJKG/2bjV62m7MnJUa
zkGvBSOMOPZYRxlW6g+BUBDBR0VpYD4DtmeXHTbVbliUqm4t6zPh4OcUkEEW2l4fZBv4YA5+LTyo
Ek244ktUZkIeazRG0wR2m/oGbNH79a4ufHZE9HBioEENJaiqG7beopmV0Tk/tokS73FSojVKGyGf
UTAUPS+m4RnxaE3gMT6/ZnTxCBJ5laVR2+feWdGih8Eez+F8q2gcWBr26bPt+FLURzJZCXaGdYGl
s9d0ZdHNmqCiBuXAQCWDLNXwanTjFtsGst3PUvFlqktaLsUYzrH9MdLCmb+dwWqKji/VcnbpK51o
fOlFd6SSwjSSLaquhtv97YVSnKBfNUYhD7UPzu0z4plGyGaabOtJsZMi4rD8O7km7udmxcHf+2hX
1dYjXzWYVtIp7DRgKSyUmMgIaxfVSvdXtR3JhaDs/xkkzqNTPiEkW/R1P7Vl/Z8SJWjbplZsuM+i
2iC0iX2dWuEOhmgCuoV1/yCQHoJClbyxZht6neXEMeIhdWFsIc686j67xSqDEwsOToKUmCzYj9I8
gbYYDOWSK3hpGGJy4HrbDnlrHQ6bRhLYalDGwSYXX0nfGbga6S2vSlqIyRB1UmVbM/gUrjwB5B/I
EJU4CgABy97v0kgQs56LdSj2WXbl1pstTMRgRq6Z8n58Sa8K6DWrD1rMnBrMkrsRy2nmT+zHWgjy
BSMdTn5H2Cj3d7qsmnE3ltc4dUUA/MzxlpyGpl/ZdKREF2cDwgNtQxcc6CfNlmWBsyASLcLTKBAx
3BKzDwMB77n5zMcVWulE01OHftjrd+s6Jve13MNxGtSzFPN31L01noxJDblu9Bw3TO3BG5zwu1cX
xamN7+v75POj7jpbN3lBqUR0IPHmaysyxV+Y6ZLYcm7FHN1+K+u1xcuWFPbZwhpZ4o2hBR1spk0T
j9laMqYZPwW/PG+yjhSbK+JSdEzy2D95gPIilDtKz5X+FIxeyuFQu+PJbYpiI3DXE1yJguQUaoCb
8YbvDL9s6iEZ7PCajGnc8hosDtyCQK2TLD9BK68ydU/24oLtBc9AN7HLRSptN+IrK3PZ9Un+VsFs
kr9wb7Ixea7Qpx7VJpyVq599imfjnnOhF8AZgPhVtZyHuwSwrDXE8SiGQsp0sgVkPy1551ZuV0th
0OCqFhDePSpg+F7rP8EGABAsh5jjLwOpZZgIC5LCknNkfQp6MPPx0HFjqcMMP+H+WLGnSJ9EAQDK
zMYCVx+TigBdB8a3/+BUXAS36G91k4jq1hreyns26fJS46Pd5ug8hznX4NBlppDzhEpKtpVJYTct
HIU0un1cx8NFF9aL7/ytBpCroWNqe/M5odyZVDx779kC0MXV4qlcoietetCmATBmh4CfpgRq09+g
vL6DgcWNkY/iSderg5QFH6Hr4ozDuvDU4qWMRqN+MXXaocsBCuDszQPrx4kDmz8CFGRBWmbAYalh
HDD2zHhRLCUahAFMwfp5w22tSRLlBemhQzNCqdpoiUXyn0OhhGpqe/6r8ZoCC01HhDNnqpZIFIZR
mMQ52z+nkNFaRKnUW/Nes7CVLO+dlmSmp0LdUlKcMXnpxWWsoD1eAVbyUamT3DOIQrXXhk7/hDEW
BCGpg/ZhZeqKcMQChfSKow/FrILInFQ4XyWaPcCGqD9RTCneeawwVXbO/zcNbierpsDI9ENcQdLm
ucISdUUbciKR+w2rpw6s0cH+mnZUHq7h+fWIvXIV7zFKIFBsMJVW/z1FdEb8r7cgcE2JooNgntTt
GSE4BuZobHLIlm/QxxnSz6VO9QT+CxJ0FtssuVbPrsbDA44aU9FMzrs6iWKjo9Ti7Bt2WcVI1uGI
/B61Y7X6Xaw+p8pgfsW5scTGMC3ziy3pYkb5apOMbrY/P3pvzA+qqAYUoIaBRWol8kQEWt96JA27
/rPsgyCIoPlOp4/+6FDe/dnr6TnbAoNO5XkZL3UBKlWW3+poBOHc33f9BrsFrGs6hlZSRhcY+Yfn
Vwp1XqQoQqmAmgq+U+KZnmfcY/+GUdzLS0Hjy1zJ8lK8CAt4Ibhj7kfOmJdeoSlUZQ19Iu/33hoM
C4EI9qJ6wzq5fTah44UDcJob1SjRmZrv3ArEa+jv5gsr9+Uk/YSpAydiK9GQmwdbZURdGVIKHckr
8paE6CHb/oB11JI1PeR/u05JOpznekstlanrl88FseyTKMZwX7Eh/tgwVpPBMzR6QMb0p0LsLvxF
pbQ+JGNnrLf144741NFSIiZiEo4bxmEmrIpFEmI1FgU/afV7CQ0gjxrOxEyb0S8K10Grq/2Cw31T
F094wA9wD66ZCIgI5tTt0ZXSznd1Rh85PvgWNdx8Z0gw5O2kpHzwfdMWbME4rWt0oiqz+Y49cGzU
Gad9D7pofKG18yOpwlj23iRMg8DFRUWCPFl5bUMJLcjRxmlIS0/nDt9Ja956vVJJMtf4X17pkCHI
F98rlxx6odNRJMiWMQmeOTsTX8jCPvOSF+kIbJqA9krHAkjTABtF7c7fiDZ2e0P4rumE6phtLcn+
HSebqxxIknU/TkyevmPPlf/2feMkDEJ2AQCtDpYjUgykhpyFT6zULSPd2TIlPA0yyqsOpR38C/J1
3ikrd3sdiSyw71qrRHRtDOwg8d7q+8ZpQdwwfX2DiL1sx9vl8vrXAF74wAB2D3YYcY28Wqu2VJFa
oR1xsIRYuPQZdAjle4Vs58Snr2Nvy0eyA+AqQewWQ64APp75WfH9/5djABI0CfATemtEmJ8cvGMR
b4mKh7rr1gQEM+rm460aaO8R34znilC2MMnVZjpInYmgWmJKQEnbK6ZhTJ2U0WczSVeanspoZlw6
dGJzD/zcUaxXDt3JJgP+dOw7GLvjWjRqX4pbOzjLsPqF5shQqIEyI9P1HbcBFNy3+5C8aofSclcQ
GKE6td5meUrYlV+hb5MbeqVwZA0LwR2GOMgWcRefNbVD5VtdYiLnGkMJFV2ktHB8Bwa0QJtpng7Q
sCjH4OVCHiSbhyatRW4IIhHGDVC0LcYs9PprT1StI2o4pUBIh7UopIGHXEmWYtPc/IZbWHNf7FVt
WH4SOf93NXjJjNTkOs2VlbO6shaV+vQrLQsMprM82Yee8PSwcWJIo2p/USihf60Z7IC6AdU56JRX
9/tok+cnhf5rnHSrK2uDGur359X4lCMAidyWFOyuZ5ifoXvqW/NBHadu3la3v/nzjIr/liDaGabo
C3FWTUxpJEqvdI05E3DBP+tFbUFm+EZCEWxVjxeGfO84o6DMNH+OinKapB7XRxNqkGI+B3y8w5TU
TSEWgrYdjhvw0qscZ9NVZNs/wcVhN6T/r5sP8dkssF/pRr399GB7HHKVBYaCLDniISN8/Ks4hiSk
JQkgfCsrHH/dnqYvi2l6E4GjxlNTqdbVKEpTINxKFft49oaKNxVFmeWi96DMvuyhPgEW9EbTYTfO
w08y690OyUzKNvqycoU4Q0eJoytPNVChiV0CrT/jUaQrgNdE8Th4rneb+C86opkAOfFFT8M0cVnM
VLgb1lPCoSB5w3QEDMiOyCxkk0Va3b8JHzxAdaSosWykOxnmvtKDTyKWQ3pbyaMB2aGbyrjX1xhA
QslBOqLjLPtYmVxdgwQHw9tcDkaY9HeFbk1oOuXauM3OohmLC2wm3fmqksvEjQlWM42pVq5zgp/g
1p8FVYIsIoM8Ee8+70I0aa4MvrpIE0/B739ieZbAHtGjlpYPNF2xSN+kuatOfMEFUnvxBtpO7iYX
9Mkg3VFWAnzec5NFbueffjeQxjU/09S5PAZiBByCsl/EELqoCp++99lY/YoDH6mUCLdrlPZfMrK4
ToRrE2HaatH2G6B4T80390KUxSX9QqHCI4+1E95OfEiXQhoDrC2G2bY1xOnOTqNYEeOBE5u6lmXp
qnIv+DEwtXdR8Eijwu5nNtZnVWC4gXtwRYHI+ujKFJX3DxK9BTJ1lw/7ldYZHKXXdvhIzj8SaaNg
c6jheIvfF2+cbl+YJOHWBa/Dyvs2aryDZLfACS7idezGAbo2G3VKJuCoczrsJH9HeSGaquSoJ3Dy
M6AtuSIEAbLmlB4qTlD3UkGytbxnTGiIzt/bce+TJt2jOF5SZBSVcTDmdc2Cn8q/GTPfnUcECDTx
WcHYejxFEBzj2OMRPUCd58HNNJBdb61q3OyqQ+pIogkymAMs/KyTdupANoSFF31nKFvOZjPXIkhD
iORyfDawmZyd6TO5bbLrn6Bbz3AgTEqt0uq4GKIgwz/9NXzM/gV2dOUaWmf8fF241QQ7IfsMbsGT
8NM557cN4DI4Ik8AoV99ZU2/21BYNHh2R+lV9u7YT36vyMaRBhcrIoHCWQmnvVaJ5OXkCIvIat8j
QrLxsHkX4KhUC7A2TV8jtt2cr1z4HAM7KhzXi2SPhwF6lmytMHLMHDwA0Xfpp/82dvH4mG8GnfqQ
QOvBjv2VEow0vmbV1vIAEfzEzlDGI2csx6yQVdo9HlNn7UTSGpJ8tB1/HGq3vpq5urSu8poVD9vL
bpwZGkYhs10PQuaW9XHT/6cqQ15JVzWg8Aq0G4NSgpEhI8B+3Mgb9EsRtM2pKtZb1v3eM8IAaJnv
YTII/khnu+tpq9XAB120iME0qWnIGtp3Ife6Fa/EL5VdW0H6MXFq4r3dl4l1nGyUoJAWhL/7T6YM
HvqEcPhrlIWWqj6yMZJ6A8/lUgwFGqsNJPccnsvSI7wKHdcRRPOCKi6lmPfXzesmAJm3BMOXSQhM
PHW6PH7qYPvDFUuJ4q8FcSsWwDWTfZ5s8ZZgR8vBTOWw4wzhh1yucJsLc6WY82jKvwI9F68NDQZH
i9s+RfzYibLY91zYL0C19apYti/vA7YJvRZgV4JWHJLHvylDaxm8HRz0AE3bvc8sblcWlAz3d//p
VSMfpo/RkaGwO8+rfEECs5I0Rcz+axi8Z3Ifj6OECZMXH24YLSr5PiZpV4GaPDUuWhRt1sbEyu+Y
+mVQwkLfybaQtP1/G9eEdcn/JC6CTbMsOHNyO8WF9gKMm56m1myocXyMgf2Aba5CEBmtkbJHpekm
j1H2QB+LLRO0eqs76OkaA2lahM5Hoe3UcdnLThtyeQbQ47ruQow1p1Od1GMGFFz5KUcPHBiVRECC
y2BIvYQlOaE4n1M10oe2RIJRtIH/fxMkbU+6DDXyYPOPcqy0i2WSqyXMEg8y1+m3ePIEDwGoVNv8
BxKVYPjxATVS/fKIz6d+v3M8rhQuzd22YC1SNYoI/xhkwfYxI46AItAgzCNex4vy+w9scNFoePqy
5dxENkf76DDJVGp/P2GzpAsKI5iANQAFPQZ1pNpR0sUG0RBXOwAocLe0Va4/NQZ05B8plHvl7iQJ
SGjeS3J4ZlPznPlv9pLucKr8CYKWQwG5Uvw7HPj8uknsByVnegS4MBSSl8bMBVdz35WAP1NwGf2O
DCtRcEUPic4bmu4ZCDsurtcLOp1MtUBtZKZOmXnTtzUPOE0nvqJL9n9w0yPXl1E088ofvXMezdKX
4OWpRuCZbzNTuiH9bDR4/+v6AxSAnuLIQ0TWIuRKNO0QKBUukPKa7GVXeNP4uSSv64KocgYaSjc5
gLEj8UXSZSZgOutHb4O8m1rKeYewfnjmeqZFkY/FpQa0EoZZDi30uwsMNxkhaF+ppCTZ4+PJ98oJ
wuFfMNOo5+mnfCB5jSloQFQKKzM4dwhXMZQ5nDrac5FmavgEt5T5widFggbvy/Rw+A835260dJmK
xvnc/PrdeuOsgXnT4WoXW/E0/qGWPD/OXIYaBUTTYq4DQUxwZY2dwYKUKOO7U5rjzHuJjs2QYwQj
/ShxMKVDRA4UIXoP0dKf4kSReOFYsMTLGkwKk8EW2up5FLxoKiW521DMZQmsXQYkqFHmnUGcPp7w
hnnmwp/U+Bs1BbWQmtjpxnn87vmKDYnILusvnvWyzdhD+M1VpKu4jKP1RF7iHQFvW+GOQCEZC+Vp
pWShT5geRIxDCEE+pAaye0SuKtRrmxLi1ccBKJgiI37uP84VdYhXsAppEyeGXhrGssZuAjmxYRud
UWN5fVKF/o58D4/1qYdjjI2iEZqynLhMzMWhidmMh4g//bN7YNKS8pe83Sd4V8f03tKVw4zdkUUS
1Pmyb0MwlYR90aOToxTi+y7KPtDBadTPWRZXaL2XFXkgh1QY5p6onsm2ca4fM0lTz1Iq8daAmwrk
ewEkgXS4/eO5hTTfWOQoKMgCFyfDeNEHQ106Vu7i87YQQYfFFX08ZMxr0ECxDx9tdG8cW2f5xKEy
vOtxMUi1EH+gJaOEP62F6EwSJqaRgEH2QNSPhV9GIFv2dSkxNFUyKE7dOVlq77IFfvcIq+njdltO
x4iqvBE4jjwRrKr5EaZBeTqFe2l/m0k/mVAFKyCKqaFvogotwS6d8clkPvr1GH4cNW33oujOGVaa
e9n9NIjpREhbyq0OQIrLzF19BRlgvLhq9J7UYDVh2tDHtOs27p9v0TzATu/TE5TpzhxGS25Po26D
sRBXltFeWXb4/T6CsTy4t4z2PK26UhYWAcuvipOgi9Xkv8+F47Xs1HshfNOYlawBnYdJzdIEwZOe
4Uel40OBJRfuZAOBJyeeLsZKvm9wiNU5UWwFBTW8wxjb08xS6aggT3cPWEQwULWMt0/fvL5pdTXb
7I77bnoMmDT1ux1GXvX3PxwG7duoGRxz1mWw08MSp+ndaLyhGIN8F23V6rS0r6fTS+J3/G9z6Vbc
3EzKIk0Yg2DjY6NRczeUJqSO8QUqr/5FPm9joQW6xqe0cqVoyfri5dgcwyzFMcfuUk3UgTK76C/o
xKKpWYfNM4quZxkcnFFxRX7cuyHb7ZPLmitAAWyE/mvxIUsnq6bQLcZBYrPaTphpnfWADJN0HUHr
AuWbi5ZCpo0LDzQ1xbo57jze9FzDnPVtzcrLel1KFnRj9xu64QfR+aDJRzyra5JpwDXuMPHrwjgF
dPr3FX48qUHyEGgTywUrzYWxH3ZXKdmlHQsZFtONvP79zLm67tzgkj6/FINpLyE7FolGviOeNJop
iDeF0QzsJUAktdxybQlluAA09niAz5tXI15BBFamszaZm38FwcOVesws+LltWgrvSJXzlyfOezg0
N+OVPWkjyf3LSysh33oFHwNnKU2AfMyWd7T/5zYNmrTM2f323jYqfsPCu39o6q0jO/l7T4p5aANy
F4+aOr/QbcqhyRCHmdvw5DgAs46PIhRjjWGAv5qsv0L//HRAGJveyRQKtZSRy5WAqPoOecsu2b5k
95gzb8WqCZ9nlPulUCRRJgWgAHfSn/s8k8Dsg9w+HXcPTmwKkSRLe4YoW31RaBaCJRN4BI1kaPM2
cH/39NQj32WAsHQohAxXJ66nPf4v22T63sw418ulYEl5Zy0pgms1GC+pw9dNoKjsbK+ssRCnrRye
RlxeYGj2Q4EjcMgciyfiY3fz5MDBOx8vpCIyEy79sMwIOc/KGOJEMXIe6gALNL8/0r+c9W6D+mEz
u1Q6CsqVDUrhC3ZVadJcwZ7IVhyUowe1WMAM1uf4Z8vAvqx4DTY/fVdmxqkNylplPBaNIEj+TCtR
Ke09+4Oi53EaWNvPrX6yWcb8+p3Cjw6OXX5xh4PulrDcifDdl9qS7NKm+Kc8INQHsB7GBKWqnOzD
wSKjWn2XCwMzWiOlL20TwIxoxXD8xqqSE9fJ/rXBVlpBmsYHUjcw4CBbCoxpcwfXw79j4qneAuRh
0cfKx8iRrdUvIfEobSzDZ6KDSODEiL260KmTWLcoKPv68Sdv2IXboQtdKYyuuw78ae6o7Z9eOjdH
4SjJJQ8m1QcPMk/dbXCOdonzTzTfwBHJ6xHrvxnAv+mZ68T1vrKdN+BEC+8A4YvEyXqaiIS9OaZD
AnaUVG+aQOiVMI5B+uJoD5dhWGYhvQ6Y1uDIo5ekq7QnhNVBEvFt02I/kKf1JDxunfqHJIRHo4od
INkAqSUK6BxJq2HwAOAOX5XnIWYejvKh07nGmLteb6dwrtwX8Md0ZyXFnP4e1cPId5/9azrYBPUV
oP+wRv0qFjfUMldVEVdtzB9iIkF8ktEBUVWjtvjBt1FR21E3JPn7CR51AOAPN2QpNwQ1sCDIXpr0
DcnZWB37xstGX4TxzkTq8x0twoX6dAdzBP2f5fYAt8Uosp2ReJVvYllgWQQ3xnKdAWAanLcd0Akn
OetoSl+5pfK1J44PPtX9sO38p29iNdw1fb+Wih/bGd9tj6F9UW70clQqIn4nxnxydB25KQvCvC4b
jD28AOEg0XXnNOo0KpTJTSDj2UqFno7A+BdcXj8WAjBfIXMrIHs37Fz56PFftDg5Jya0z1Drh4p0
CIiU01zNuUxbW1oryUOyaBqPE18/aR7qOoqK1eI974acDpA2wZuFzGxd+4A8qzYukV1OhsyzLTNN
9mqyWuA/lLvCkHK1Od2CS2Ue2ZktAp04dsHOpbXTsuLWqSCTPM2wRPJdSqhVMgOagcaCrIiCGKGg
p4roYet1ymYdhF8DMeuzUgUMwGJCZsx11W4tHxVxdjlmyIUmAtJzGF3bPE1JLwd263Y9ERxppZOD
ccqaxfWncHMYjcE18Q4OfTndzxRvWuxaeqz8BHQZsdk3JZ4RW1s7kcCtT55nqu/7rxZupNR0n9Qe
UcLzVbBBMcPoMh7OTCps9uUNJE761gk2d+pkO1h1KU91eSUzFbqatTp6tZS+IbOhmD418M2uJRcL
ePFvcVyBtYg1Hyk2GyhsbuMADRq0oOPwu4qTQDEIHjMksvZlHTjNDUH81mNMNcxSNJVdkgl9sE+J
qkHYqe3Cr++mdFZza9HAebIRTIeGmdMB74xkTuTdl4847HlZ1zE2I5rMPLtg+KLlWgwUrHJHJ9r5
F9bTVD6a8hijYABtlJ+6dL4giB5agjiHUg1+4+KYn/j84kyvvYj+oDlAgDbGpZiJPfMvhlfGPGc0
jUmJzxDbm5L0tAGXrPebFrY9f2qjgkTTKvKx2bCxtehE7S+BupanpupkwbvavnZyBwTorDiT5622
zZtl7TGbFcZlEWCsMG0budjsYnkM/eZQvBNkrnejIg3ttTkFbGoQCf6FQPvlMXJ4TK4YgVR5HIfV
JqSbWxi8ElpEgn/2qsR8m9SJWl44FtmwrQ4fBxlTlR514z8i9ZRyn/YgvPSamIhda+VLwM+GqEY9
3Ddlfzv117+bAfroiXgu/GWx3+Pk902VO6SGzkhcgHEu6f+sDrZbSv5x5WiLIbyKsu7Okuy2jSfh
82O8JOXmMGn/DUC6dgcIbswPed+HA3JMpiEcEoyTfssgvIf4IOSRbZCjuNv09/yZfXPLAxXKedOE
fYh3UX0i10cGyzjVdETuDsiYZzRrqmZ0/QFgZdTUhPg1hIBdRFRk1PoMUJwOuPubFoikcl88Apii
MgoTsNhyKqheSvYqjVmXOwUY1jdbiHCsfi3sU44QrwSqI+SIbMeBQjgkzR4ziBLSBp8QjHB5Pmi1
BH6TxpSlxizodWZgEYLQXj/27cAaLlz0P/23V+0akoTOpoZzHG5mQuJ4QaOsjMiRRmlUYuePIH7O
WsFI8Ujq+n5jt1IYfPupEl/wyIU9sPpBpDalct+w6GVygDyDc7jvi+lYCNFhK8HWo1PRS89Ndfqs
r7YLeS7wrlWI1L7duHGaVk90wQDyHszFGsjd5U8MpHB4iLcCo9FLXY3+P3ImmSnzZ3k3ZUl7laVW
N9vhG7yzeieGNDfNwDYjCy1REAqYs4lfbDtzeaR+8ey38cBckz3SmTd9HI/Go+jZmRTHqQfqQmc1
QwmcR2Bz4yeWM7h025tRhzOF8vwi361OWmt5xui/jV4/xvgMqW8viyVgANAiO/zUPhrLRsSEaXVS
H4hiSsrGD5ksehe146Q/3phK9bxdJD6gDmsuDva+U9awCdpOujzGYErpgcTfDf2stFC7iIDubgzf
rISaVsnmBANtRKMmkQazry32UEqsWCGEE14jfGFfBkd//amoPhoLDEbLf6m19ASESIDvfPMIpj0f
V+eu3m8+AW3gTT/DT4E31JjjfKs6N7t0BjpYbTCmMw8hZlG6D/XIn+B4927476pkAIcmLpBiSiJv
D393CKgQzL9aLrBDPq5KNzBVxAvM4hfEmwTe/bN1d1pWBSE6yX0BcrxDqGLjcvkZvUcSOIr5pguD
pokefN6NDVzwq5JZFJe2mC+/fCjzxljv5KPrmYgZ7b3S/+p0MNe/FWQTbFpMrv/YLPAmDEYZleA3
7WtjGzUIX5BVSa+U5SS1t/W2OyyfY+DVw341a7jYvG/gf+xwcD0RcKpLp6GmsQDt4mpBoSZiOezB
PRuEpSttwQ1QUfAQhyRbOURd9kOqr60yxIz55bXlLGfpH0sgS7wo+OCTFbGJHRd8bKb7ojVzlaPF
Ljg3WoCbknIvzjw8LsFJvgg+mptCdUBfCBU938yvkdudUCDGmrIKFqm/FM1eCiPsRDe8a7oLVQUl
osavTyIK3XShQjXncUsTHB4543JN6eZtyXDZimD19sw7wbblFop0faAjJIjVpXMG0raZRwylxw4F
Bvw5L3hSOGyk+wySOoxebzhb740fKz+bK0eoNWFxt67r3ZRUhhRZ8ss4HV2Nox4ovzQryN1Hymxe
+LKG3VK3KI8U3pybgvGV8ebbDnfu7G+adpKhX+1lEEg1RQF6VAss1d98+VthySwnmCxT3QFDvfEr
aeDm1XmnHhnnYQogXuzK3Y/1ghD7j46Ahmcg2w42LddQUFOTkVN7iWSyOA2pT7VKpXzsHC7XCSyp
c37q6bsNI1lVnW560LrnhRDyaxV9hKqTdoGsVy2XWDqTQb7JMDL3/ZLjk56MoJIFCJvgc0FZx3qt
/e9XKvCZy78eL/vYo5qTU1eUbno7s84B4tGmQP2DvH0gfhtx74Zw030IIQa/VJr1TKGfeXHnZZ+o
0oaySdo5iroqtpZ7BVW5uBT2E7CYXTntLY1RX51eiW2fxqu7YTGvkkhKLA6ubHzyjhvy/CkPXyCR
hbSHOutW07qOwFQI79BFfmBIqUiJWLPUlbYeUaDz935VsJyl6k51b21Voq5/2X++/ZtIJjZqUrA/
z5JsFJleXVzi48J4X2TpJJdd4jdBIXBDBZdWkVN6SXVTJIHdxBIiK+gOh7hTpbCJPluhKmxHv3Cp
iWmzTu9lUw35b1c6a2wqegb2eEfuKE6M6Xj7IKZHi0nRy65FRGcmJxkDgNka0TnqdwMdW4lIHPzI
A610uWTYQeVJ8DaGs/mjrn9JKn6YineWWOOoEB4/AUA53avS89Mx8dGI4qOSK6Lg2VX6pY0nc5rj
wcfewjOyYg8loxuvs9DrXqP58FhtYt/CKaR86l1MlGcGUSZH1MFEKwHQHFAc0lG+w+srJyntIrIE
Sp/K1Y87utpFWD9luFn+ehvveWoH2073CDgYowEznclofGaWKoMkbLVBPik7uVlxRnb65LqooGJv
Ylpx578/uv/Xvd+rNAEz7KeW7kZFvV4HzRySkkeRRRNKM++eXADYx6b1K17CzAn36DNqYIHWn5f4
6iwnZl1U5pHsnmC0cILwM+GDSNL0XXmlQUJcx6zRuJHKHYWzwU3jCctv0blStWFxt4axBOgJoc23
p5Mlxy74WEet4uis1tBjixvo+pGH0gNaSb7z79h5IzKE+ofUkyBVg4xP2h8NO3IUTCXuSG3RVjOg
+gH4CD/zO0zSyZArXtd8FA/oowjBrPEI+53gdIU0XTBHMhie9B80G86/OEBZwT3QHkmvJW1V2Nnj
SNpjhUF/DvOWGNikfg/L1HqQF9u9OHp4gCeoQWDNGt0gxGhTtk6reRN8xI4zJUK/qLG1dQc1Mh7K
nCgckfqRuhdyEV3XkSUr0BygfQGtC7g6v2qMz3JUHLiwXJnLAZMgkfVeCfr4Q3M0u3OsmBzwpLId
tKGmiPlVrkQHtJ/fLFSTnrtkMZuRSPMo6+78YumfoHKZN9Y3YlItvOHv0oLVIGjVzaing44rsrt1
kmmNQAJoUB/OL/h7rfcFbzBoEXpMGLD45SXFWA4Ha5PkPTuaLKNNaIEF/DG9VDOMwyB+t4fSAVX8
rzTnXAATtizai3vF48TCusHJE5DJ6amPDLz/SsgHteVMl3lK3RtctbRBG958+0YmAaAztv27MQ5v
vsH+vO/eNlsh7lxcnCoVyQ5itPEAT5OtGAAQD6sESH4hAHkFwpDo9ckYtJghrDkhOezIPqcYB6N7
MBOtB8HFnKHNVCBdjM//DZFtjVch3PTS3b5PqK+eBf+86z948tNFmgEpZW8GL82KvHlTYOhNGM7b
8R4jSVVbvZRm1NoJKowQ+LfNJ4R16ZxbEqXK7rVmsGEc6ogtp86sT+v+4XAp5Ip+BiuR6kHkvMFY
8T3S0YFrL0J6mWOo5YbF3ksWeInE+vvGYkmVm01ItcHxoYd1+y65ci4e3Ksv0hmHz2v0Ad4cmh3r
O+tawRQ2jwD2QhAWMHrRl0wQ3p+BpgZToc5bkA6oDSJp0MqsC+cG4uScck9XFbvHo9y3d9xYBlG9
70MuIt0gu3lqyrip+qUuInqSH5eV9u/9MbJ0YUbI9U4keRAxDwzXIeltl/zqciPYva5Z+HtG/JZK
4XhkBsYLgvCXEFaGvXsHOni5E9IUPHyhCN84BubDSVjRl8blk72cTQlDpL+oHNq+IhanxVDuXMBG
PdzFJaAzjIVadXTXEpiaSSww7NpyudpIsQVzjqpMArtH4RxIUmYOYn6jIPdrpnhUx4iF0FzRE4zH
xUFor28lq94gcSlYGCEmutMZMIRcoqeRtQEkUdVrcEXwc+1nHaT5PoGJaq+tO3NfltsB5n5acsRE
7wsGyGTEPX2S3WrfqlKmQglEhJFkV98nkTbuB6hyWk2hAg1Nzys+JNTRmpYfG24WNMGYFikhOiLI
cTYneoNhK9whx0Mbc8JBm5eX3WY76he2znCihcRvGSSZpwxXDQuY0yCHg45XD6gdmUyrKVdHb2Cl
lwH5u9eW7oLKkldmqFmZ+KZvUT67Dv7JmBZzYQ8m4s4f8t29q34PbEunMxrTQU9JRXQZsEITnPrr
K/40QflvoDOlB3ISJDau9wRwlrT8ZCGW9dB6IQTytqopobj5UmPNng7NklcAoT9l4z7nGYw8q7RH
1Wvp7xQF+vWNAg055/KUu1N4hstdojZEg78RwYLJEjuMY9xlTgWCubUlrZM+uHlJ6NBR9L/mWLEA
JGe1yjyJvFcrcvOTsM5A9he0HLvL79OkkzjQdXxLdSrcYnIgom7cm2JUKngjMSxYZQSC6EwB6+5p
9PVEoLZG6ahAILv2+J7x0+maAj4rAa5i9pl2v1h5QCrQD/AtswMGo9gYffHW8g8Zk0WIVTWA/O39
b8/JSd9b9DKQBggZe8Pf/f7k4Q+whpIPqfqs4lF3OEtUXMMh+9EmjX5KC6IO4tXc1QyLirP/FI+n
78CkjaHJmvGzzBj/nYg1FKPkLi6/xiugfUA5ivv2NFyK+pbkZK5izsfsH+AjwTgvbl2LllogEvAa
3RUm1lj5zU31e4PapPIr4QGemnuSzbCDua86kFjVEMqP3sV+GzjgtJyvMjYIMdRcuuPUrHUv/61I
YqcwB09220MOijk7F4VdSe1ZwlPfaPdkKvZ1FF9IInVyKHt2FWdwgXdWE0TZSTHEgQ92/iIxOXMK
GXF6aVeZBoVVZ11aCy+0DwXQdP0hkSRPB+AW8yQw1tEpYfIxcdqZ9UMWsRdzAIgh0DNRz5CAxnWn
L+X2ZzTdH7zp9erxKj313WyxsRpof0FVAOhXyvlkW1818z8oIp1LU2y//xDU3Cg73f5gDOxz2FJK
2cJpy8VGQlar5XmOPcoREW/8mvOGR0mDACy0TmPSsif3XOd4VR8xOS9NwGZqYuoUgTjjbSlkAYd2
1jNftoY7dRQw7KEKD/pmz41SjWXae5ejW68GU8aAhzL5DCn02Nn1d8ksnu0F4DIWFDGGpgWmJ77S
cwEO91jqIDAj4NszdxIto1G9Lh5bzIG8Z/IDz3wTHZEqmWdSyUVYK6i9KTky0IaDT+JBvD9Y6lYl
iPj4vDPJCu+gEVQ6+hfrTGmUPUCevzItOrz38iSx2DAdlYkf2s9fHMIZL/BMm2/BBqaucM/fkDBo
RWWN5cu7VnBahmLZ83kJeRAkE+pg+u3scV0OZ1+J0tLqYnnIKaaWF34ID6woVoz9n9KJfJCYD04i
C2oExRXzEKJgFPDzXEcs6zJxoRgAnpBgZdRIe5uNakDCK45OZVlxENnU8MVFF/kohoO6fdXA7ulu
lHZZjDm3Y36Z1jYhwgCCB78omWKm1AvV++hCZsQC9KaLeLKoBOQcuciosAa1pxa/amLdclbbJCsG
bPxCwj0xUWHrWZvY6+WqNu3pl3eoY3JlEZbRpiVuK0cKA9BnEl7IZ1YvF7DEA6KATlqJ+yDo1u3U
g4nY8IKmNc2qhr/ugdRbLe5NC1Blwul/0JV4WTf74TtJB7nPLEiMWWkKPc/Y0aBr0guX2IGQWO+r
RRWFXr9MllGN1QyhjCriEZaH6SpwPyCY6rhMMadVtJo6HO3QMLsCQ22HbUgZAoqQWRr1q2N2u2oF
ObmGUBve1yUY/+Z6F5F3hG6wTF99Kj22heeZUy4Um+Pf9Ze3OxOpcbzwQ9JHDJWPag7eO0RT74Rn
4PY+uPg4e09taMV6B2TCbN+LJPhOoTJU9+6BjM5IxlvqHVoJvBC3QudXZQJh0sXpOyJm4STFKqUK
YzspFmuB7PXh6o/31oVJz6uPTqqtXLpGCspC/osz3frzaqBwPiVyHh6R2HhgzgrmV5vD/a/g/az5
5/X4QksD3fpFsDkt6l0+svwXJcDihwpWWDbUj8CgwCDlUX/ZBn05thvE0D9oQOuJU20GWGVz/5XT
8IXoGznOGo+yTrHyGS3fFFikj35kjr9eZB23pr/VzMILVHubOT6KIbX1UnBgc1fE9RbAE2r6Xlyl
tp2aopQn+QQ+/QkIb9cdWdgGFgN9d8dLJykwSqK2CiLjhKH2E2FNvWnowSjpnbqUVqevLeQfjRb2
0K8jEeyvZZ4e/dnqWLqgwpoK+AQzVkZPKWXRd2g8dNEv/FXv4NeIQ9CdapjGu296GR20L1sII7tH
qPQQbOsoUI1xIN6VH73OOQiM5KNQ+oi9PYFv0j4Mp1kopa+v/IcvcnlX4AV6HkPD+G1/e1tMlSHB
O9V8g4CWPmDJVgoWemEuN+HaMlwxrmjYdvbBMayTQM1eY7J6YK9gBiwgaS0GyN5yzCIFqxMEl6YJ
xjvdPfQYfsNw5ewYOdVu/TuBED/wRfj7GlKNvN/1JACYoJmGYl3QtJkfYcR30Cn121S5iXlO0jLq
CfyQ9haK9sb69z8WlE3h7VxGoswm/6hNX1BeW4RPBQCMbHOdJTA388H9rrTSspF7PD94N7MVOo5z
Vh8zNm9U+TuqO5IzDOafsYI7b8AIBzQtG9BeySuGERhYriB5WOvQySWfcMWXbeOY6PH6aZzIgaPq
ub1pCh0uR1l1TpCD3JJVHHlKbSU8ceM8k4iIVk5YzfYNfhRIH4GlcByqLe1Upvn9oQBojHKw9fR1
9/XJu6Sn7klHrlbEbRGYTett0xNGwjq3dYQj38eVo+I4vayZlnUi1FnIatnXr5fmTPEgHjl5KQE1
x1BX37ZPpx76llVr47XYpH2M2UN2GDBF+DI2nyUzw0aTaKJuS18PfxUAUh3n4CpBPUi4H41JD2B3
7wDFl2cvG+oXO4XMpgcXadm/OKAziZin/YdPMi3dYoBxGe3/ENR8jOO45XH+KZap0U2kL/UW7/01
SQ6Xd/7p6WtJEfB37ZpcA1cwzZLqBoIC3pHxp+V0xVLtxbOFCqFD2GulwYubpGcvF12VfbCqGXxa
IljkVXFGZTHjto76obEQKFBrWLWHiIxtFTgNm6nrlrI2MVaS37wV2dtdEv2JyPM1FsIKFgN+3uQ0
v0NgVeHrfOcBlRQXaM90aiuK8L+qAtdTHhHmob+OR6GllELUwa3h/4x+5VxbkHWh5fzin0xcVZnv
IswQNH5QceSssgzdZ4Uv4ahJJez6aSJal+mTzJ1i1Xrr/outki0QQI+j6SdVeUJHD6OO0mWqMGSi
N8/0/VzWF4Gt2UtUJI8yyCYlYGFgd8BqWMRyvgHwYiUwIs6SLaoFB5gJOM5ip1Fa6Zy43/i/24ZD
0Yt6c2ub2R4RMvTYiXZl9aOAY44cSYue2e4ZxUi/QYMQsAGpG0VWul57fBbhrNz9/yGyNTec77j6
azIOh5F31mt1YhnQLZK8Yyfzr49RUD0NCyEc/i5h3S2m+Rn2xOsVJWjtCUHPnOv3smnqtIHC6GSq
FCJny4fDOEzgWhqWA3+oKVhInhegty3WiYv8yMF5xBSydbSjcIBeB1mm1xyN+FKVENxnIFmJCyLs
ZenSNU1FgnOEUbCHj5hK6YOfW9+IIElNNxicUqrT4e0AAknZKHHp8KXJQr25pwq1FssxG1T1wds8
PfAnBvl5SvCOzBHkePo0++Fj5O70cuQh9Pmq1bo81GbBpf5NkcNPsr5lewVc4n3tiJupoILJPwDm
swX6/+Fc7kfKxLuOiXabxrhnT1FkTguog8hwhRmJdub6J9uo2Dv2aoaKi1X9khVBuzpM3j85HBOu
Y7hPzx1g0ZcjAu32Eg9PidsKHRhXpO0ZuJ15duoFnTYrsI8j1stE/hTloTRNt0dCUnENSVuN2m/S
MGtIfV2VMcBWvMMPLCmVq/d+eCwqaAkubMt6Z43JwNl3I17SAc02+x/vnwijZZywJS5lSMDn3O8V
rwl7yHmXBFg6JI5mArwOgCcR6Pvz0WKofTbdbf8hD0vOoHhGrxxh14EGVLGTr50wU5WQ6B/DNI+H
FOwp3/IkRARDkH9ZBYD6jQkGo3sdM9hgfw/EDTbLBgrCf0nuSvdG+2hufgkPAPiS7iiR2LcgTU5j
ipke98WwfFROCusehXm9BkKixrK5Vv51wQBCOBE8FLA/dFu7FTa7Q0MV/VMALKymmTGzl3VXN/WN
wDaxS/t7ltzUNozwhiyKkrzR4LnhorhAz5mbUn8GR7IZGp8L6GzkEjJYRiWmW/JlPD640kwXigN4
0pBXV32+0Jdlx4YktBTZ1voHKTSMcM0BPKB20RA3CCmDlwcis1RFj+dlEhLgHY6h53VqA2sA8+xb
ZEPta7ZXIg64FuZj3kRVbnH4Etcwr/0Zx48DIBuPoJjByONdBrmfR2LeNuf3CfJutbng3usSnY+I
Yqq3EoLEWw63qbFSMLQtVEt6Ej7K5BhdZNg2hcOaqgFT+EwD2uQl0M93B18yXPiMzJ8iwgEVClLP
aJSxu8lEukhrsNUtnF3iLZfUU1hsmW7Im35y9NP0kiN/V0YPjT0run9KHLgm3tlTFd0ULkxYiKBJ
DwndgLWVk1txbrJqIxTEkWJaqSOmcPzfRL2w7CHwsUCYv9q1YHJnl2Q5mU8t0m1i0yBPO40DbnBj
W1VEXLFFwAKHQs6P6SO2vwtfL0at9BjVCX9kV5WWFrJad1f6ipiQ8ynCo5MNyFXXnRa0ObjV5zmt
RnJNrO6wUkPldOPg5yfvM4VJ0rSwzsTrOKJydsW3eG2FZb4EGUirEi/hNO+aYW4MF9A54k8g8ZFs
Lclu27l3vVrUefwyNlKeA4xjRU5KSW7+uYS9NO7aKL4i1V3U6eF9ondcLqDhcEm+lZ259cBWeK7B
QX51oxImLwvedSohWbndhqHz8rMZ+E87bYc4oUdnHpS27PuGdXgy43zBQnuG3zdhOs2H6xcyz77T
Z5rByimEJBnObI+sy5xuqseh6oIUO62OmQfv/N2AV8SV2NPTxpF2tunDFjdzO5snEU3kgGyRlIhI
emDMYH8/dtcePcFZ9lTIbBMriHBQS3HSBv1ugZfb21Vpe1hPwpILNFEFPwWIU6fAwAY9T5Ffg0+C
aEZdYPEZY8nlX2VaSq58heyoAADaqEva67IPSJ5h8vALEUita3RdQ4ALkQ2qvscM/+IUOFRCBQdn
/xa+r2OKY1QT95kRRupHVJXY0yZ3WSZHq60KDBSTCJFl3BNwcCep4zQMCL7yxm1YVS6Jlc8C+s4G
oHVq1xfgd+PwRb56SaVM4QXPyTyUYQsOm9KoZzKCvtUNDi0nu0+/xIaqBMPDPMyEGeXKysNHhhQp
AmHzr+LT9dKqxK6HwK6rlsa1iGnP3FSZL+uhKfvELUH9z6m7f+YVm9LOkN2Mlbo6t35NSKnx4tY7
aXyp3Q2lRrK3d3WkFAm2wsxf0ZI/1gwFptoGadT2Vrv63Kmh4s/OpTBtgRZgRyHiNvty3yGLoli8
mnsX3dEJwZaHPe/udtQvAaLHzgfYDXDrUI7HO5nLY8GR1zf59WQUrABiCvv8i0m0z/PPYIUThb1f
iA0s0efsJEkto0M4w+MXpjAHJCeQ3M2W7TFVs6cpbr+Q3mwrU2x0+Hp17HoWsMgVk07rwNs5y7PX
xLIwA+/ft79g7X/1ANnyRpBT9Ws0mq+279nulL2SLhGT+ASmXHJar2bl2pbjjplGrBYzqdFdmx+9
cK+2ue9c/EWPleuM1Z97t5iQf7weh1NpQZxkbabF4sKZf2s8pohTQu+sJzz3HkTTezK4M74AprhY
/rJ8Hb1Hv4Ogy8QOCJqP0fLoMWjHWVdhKBiOHdg+ehQNcRp8bJIV250NLHWXsBSxQP5IIhdjGZPO
/hCnoWnRONJhlAec3ZTpfxpk+wIKBCrsV+ouAvSDYcQWKGUbuJ3bC0K5bSNP1YkAdsGHTGxrNBkZ
xsSWVLFkFgURsAR0Nn2U1Xnz4/nEdUlM234NonYSjEgHauOwb6n5qbUKaOYFcMPe7uclKmlz/Xji
YUspa0AeYNhCvZ+VBKkWK0aT1R1JcKHQiCz1w0YEnIz7pLCubEHOUFmpqLUZWg/60fR2nsMFaer+
RnOsCb8BKgWRsdw5J0OPUXXycy6JTLyllMFcGbdg6YexajE8h9DeTjII9tf/s4KAYJlgg5ncMcFw
G9IqTh8t+MakDggI/B3xkSi3aAA8A8uJ7HxHR5+g4S/kFYI3XPm2WGtzncTexGcUQdEPGmFuNhyp
N7FR09/SkkCxRwRR3J+AMa16XBlveBovG/ltn06UOMHDXDyJVbLQEIRPc4FM5LJZy+F5nMS17ZmZ
FS5DHHiAFf36ahXmR7WiMxl0iBlbnErrCJmPIDrF56j5iZvSqNvwNjZHTKR0vTAQEFU5H2pswgW6
nJaQKZ/ss6nfWIbKiLXiq604Y9233uMxSTbnwKX0GoWAsHZT8dGySYTblqLzpfimf43sE935xm8J
7oa7OonHUVy95wtMFNQFPjAsRGFpBCY8BHjodBW07RA1Ac+pJt0ZeFRCWc/9FiOZ7i1ZHaDFnQfA
il7Aw8letrxko0O3VtMTbzDn2DHLpC2EN4xz/0rRUNq7L40J/SAaKuxMLKLKi2wVSYHOtw3VucmX
L5T4dCpa81r7Ors1mxJecvVibZpWqD2XAq6En1d8YOJ12S0lQLur6Lr+B8gSm7TG7Joz/p35dndv
Dtd/4b8uQn7690zZsXWiDZ72h0INa8zv7A4kulbr+WG6mgefxDNmAohE4DYW3F4oJYq48AvKrTjk
T8d4zWpzITRBVk6Hep3Hw0dWhbiSMsRmTQwZY9K2AHC7wfIzD9ZU1FfY6neAeBfR/BsWgXoGOzy3
oytdBHLRGC3o1BTUbh+ajfood843VMad3s7MEJKRhCMJC7cKytE4IDFxzsM0/jbyrNThtiA+DuGr
el5G3f41IOK0E4xFfC4M62/jNvIWKtyOOSAN+7MvtwlnrO5h0mKRUsECLj12lwxwBk3w6dm91kIW
t/7ZFhEPrKEsLKT5TmNbT3UrvG1QLQxepzYXbMbeTvcyAFDXLH3M81+5C+tom0DK+HKgx2ADteuk
pWL6aqrhGQPKem92yqg3HCyWTek8UnR+9X0QmJWLiF517fMJesn11xqmnkrqd6zw81EtbG1Bm+lg
U75dUU3gRKoXevw8xxYv3uPxukVbG+J2YkWXxBlitC7iJQ2+SVmBz6Y3XgnaMaOjV79n/kX2xMU6
by7b124tvJBHSEO2lrhG0u6SAfIUoyCncYI4CHNRZQe+MeX6b29d9EuqqA2S8b8c1lX4UdKxUymM
ElbAyEonvTCMwL6J14XOBU9LkOKwFFJ0kMvP4AO2VqeiyCGJA03wCsCrXb2VMpqCe+KTryhPhqSU
SjYc98IvhGObxeQlv3ZYH39SKWFBwuP8Qd+M6Mhte4wjG7MRkOA+rdsSnyH35ktYBcDNWMMp/aW2
BDxXBIzPDazrYtM8+IAp4wRvFJCQfZxd4cZUMYSjkEEoXwoqq81OVWEz9pbiNyvBNmNyG2Ric+tP
JcMcJXxHYKUAF8KrruxvvenV6yAVU1c7uTN39FhqXOWgaehd4F6OaGLpN7c72fPANfHjusvZGXym
kXQnYIuUjkQDk4PSoXLgLumtZi6+fyo/yMIsH1lE8LdHiz7vZxr9W+63AIumu+8zTf5x+p+RP7pT
NH+SkigpHBNP/7qKNS3A7A2Fp/OYwsdcOu0a2jTky6bp+SA34B5dKIyXsCcGNz+v4xlxr5WfSjxR
RamMKvP8AAFNMfkvsJcbjnNGiCJ5kp1we5kc6+S908fe+GuPb1s69v0xe+X6oaDZ3j9DLrLJmR3k
q+6NP3Iki5UK+rk4o93Q28z8OCcGH+Fznw3FrZdP/85KF8m6w/qHoKkOFVThpD0NsDqFF8FKwZiY
XjxkoRwTszYfsfor+cOxP9kGUv5LylTGXeMElnuhJ1FzxkszGxqZmJh7NO7m80RN+1S7Mc+7fCEe
krIlTtAX27zjPHKOkforKUcNRqrqeYk1H7mUMMcmzUt3pAYasQq4n0a2NdaNjiS9ny7yHd5CAuhp
pudooJ10PHFZNvZ5UJsLRka7VY4Dmax17H/ZXfk/nlaFqEIYzYpilJWnO7yYgCgbTnnRfsM7tK5a
q4x2zsl1028X7IxYHjmfAdWipZ2U180lXnWbQaqRSf4d0eAGC9daMF+yFE890dsSG1a+FBDfHOnp
fSo69E72h2ttSadO071sYQVIKVYRreQmTW1qoGS2MwECcv9KBFebSxcemDojc4MEZW9TVAKvUUdQ
nai14B9fg2U4ujCsChxe4miXXficnShsQVdWsZmG2bx7F4PFbf6BSTlBQxCC/A1L8Cp6neRCrr7R
hsQxrpFBYUfm5j+kKjMTKMqRiJ9I3J3ouNiJ/P2/kWBzyUHQNSE+ocrXAXTBbeWbQIXVuYAd2Qav
WNw3UnzwOJG8Gj+veY8oDuGSaITfZSjuQO9L3Rid3MrHpFgL/Y7gcuZ0IC90ejCC8A89RPHatDiq
93Y1aSKLxIBA9JGKoDgSSQOOF7JSwroWI1SdmebGKVLAwlg73gKjnruUedVDo/8URf6X/tq1YlqS
u5WH+dbUqkdSHy204vjfTXFsbF53JRxu9b7rzkrDNMJRsH1Ig5JClaHxdWaAf3MN01ZqJIOAqHC7
3eakfX4H3ZtAkmSHzBlrWC4Q51TmLg5c6A8rxfwbOqvKYZDhLD0E93IqDL3/4gaauPzTombzGy/6
SFQiSQyqDTg0eDQ11C3PZ9LxB31Fn0imec47ojhia6AUlcB77pzQj05aK3AXpEcAeNv2LkUnkU7K
+qVjrYLO2DT2s0/cJoHPI/4oJdtuFs+HLlXER3o6dXmT71LKQc1yJqr9YlwiSV4facJm5aLUCnvr
vXhrGlILOL2TYQyqmqmUTOdbo7y7muzLsR+0hZS2zB+ystR7o6IGWpV/8jXy3hIyvE51EdP4AQlJ
X3APDokHz4UGYsHiWj6jDQPt1So9uzZi+gsFPIaAnPH8VNrI5nB9mrneGxraBKyXvBrqESd0q7XG
NQ+5lcmKFaV2fncKduL5QWJm9zTbKF5OjBlcTit1Ka+7HPsZ/uSN/meOTksFNz3yeqWrcgEC4g3F
KMQDkBzLTnvj4gSnAKHPKbMNNiFu6GKJy0r/wuYUEehEiBZwWvw0HFTz6pXFE3ZF5nfWJlC1smLe
O1UE7Ubi1ktqaEBs00brgMdz5r1bBc415Sf3txYlFTdN6XJlOXeOuyvk1wmvVn9d+p5195A5k3ID
e7a8QdIY3W+pZmKZPdb90QDyFAeRyrTZGY7vKQKjSjM5oTGD9NPZO0DT/zq69NHrbtpKXJ5Yqusb
+6ThA+TGAIEFFOT7OolJmpVzm2+dhP3CR869uXvxQn4rutiK9C3NR7336oT73B2XtV9vBw2irzZE
8MAtoMwDnSQEOHbdZTSukuf3jBlIer1lFsHoeoj9OwgkRNZ0zEVPZy1mJZkeGmnkUNjtMRs1kn15
rp+612THA866eGKlmhgSlFtnpScSIHM1qP9+eTan/wiG4jdi2k0zIaMBRgS/TiRNjbu+4WZrWZYJ
6GNrIjKAMDjGgNu0gzlDIwwYGNrE8DkdXWoch7izz5fVy2vv4tFHxqxPPo709j4xzUZ4G4XKq5ho
+B/0jQrPjJKwOaaPWSSrUbj47uaqs41TwbIBc4y3P0QB2oqOp/yl1gSeTRJuvXdhZku9uLp26FL2
tWZoUsj8ZNY7XBHnwLuzRiXNARGYgmpGD3g7R4XXHRjXcShiLDR1TL+VLMF+kE8U9lb5AYvkAX4t
B8GfHPu4+El18adMcZaPN2iNYgkKPD6RUEFZ+zJnc1qV1AZh7QAbMgaaV9vbKpL/gZsxlsMRuQNT
PkUkc5ADEwB85r+0ap44ayiZ1LvrkzOp2SrDv/+DcHit2WepFGRA12Q1eZ9qbsxjL+Zd0C70cFRu
4sTrNJofUCTVFu7OG5WxbcfuRwWibqe/tb6NAhrZvtrkZ0sk0TSTU0cgH7PWcUOOUrMQH3igjeVO
YSNCWMrIMsEnkAHMwZzg00xyaAoOkZhGnLo2HW/mYDMI7Iz/RgjALGZ7fSSQj9RJt0gG3WQAhBOt
6ik370AJRMjTi5NnVfwx0MUygP6oUOVgCQ3yG8urt1f/MUDVDO9mA4LgBhkBsspf3Ur1Ze0jOwmJ
9mhdd+0xvs/BPOm6XwdvWqRPjBH629OrcxCmrGZpKhPmXT4JU4mAVBnrjcXQajvI4PximDentr79
odNJQRWuU+fcMe3MrhEYtOOei1EOqZ3G6sPbir7rUTykcw+q/7NiqgVggFRmdqXKr+L9OnSxHUrI
vG+PkqH0slFUEX/hiHOfsy3dBAjWPSq4RMqHf4BVelTFZzmYPsRdA9Y/IniUsHISxwrIxSNFwSIM
EyOjqY+vwEWbp/rRkKu0H4SD/CvO0ChPDdh2XUvJZllC5Vsc/2vEM3gEcopfr5QHdzIqsu5HmGjo
33UZREiCMHxE9gdQVDQDhjkinVPiYVst+oNb8MOhmoyt9L7Aj1wgKREDeAHXyTgfcPjQY8xWm7gt
1ZoRhKLaGNOKIA5zKkwCAFTmAHkoYeYDz1No70WwHzMzDXf/Na7X6RfCcg7WB62pC7VBUjL3C/No
fCslchaNEGO7YkxI6B3qNieT51VnpgAY9s2UdIbHpp+1HJS//eVvOexhawcrM/vJtBdS7mZO2JI4
NuI553BnnCHRvUSfTz6qAVX9nxTzqOAcoTFej+rwdTcZV2ASwgffiGynkVGA9y1TrCDiDRFPZvVq
J5tA7JtzpVzvYj5XsQZ4XR0q4bmlo/dVhBFgXA3rK0EFTyaEIMva/ElemTfaUyzIlvCH67MY3J4X
Yww1kfKJjf5hkj16Qkp+SDbLTxZuSfoDevDQnH3Y3GNiFoNwKmmvZIv9eVSTIxyiAGlnBun/DxGV
S4MH/DmNwnmViJRvaILiSQ9OaT0BYpI+jpLoLTo3f8UFwSupPVS7P+Q1M0jkIZ2oceMz6szFPsVv
qAKVT5u+Zi/ajKTi/87H9J9KRKzBr/11OFKlyVHR3mozSdNg/lRVunrjMqdOt7bGA27q2GN3j1xE
tB+WCxaliNGkmHfndhe8P4moc/WAvXB71vlTQgnOAqFr9Czx/2mMMSCby2TRI7avwWnskfi7VnWK
eaG5xQW5xk+esP2zG7oT30DaUgnkvmGtZ/FwADTUm6v44Z2RXmJJpit+jVoULILuD4pRcQ5s79+C
0v6xJ+rNZlTV1rrgLVeCqB87Ozh2QGowGw/Yxq/GT59pzwY7PLOr9V7zXLkk14PzlclNlwkIUELw
8E+w6CRMsb7w0MEphYW31q1UBHb3AMiBYii5m2Rt0/uO0pqo52zQbOtiwXdP1jkW7mbYC5fHSSvm
CeWWP5fPzjqirM2beaTeOiZ/oDiLBADb+XDYwXkn5TN6Jz6DV6cUf5laoQjp+fSkFaSLnePZgW9w
O6QQFHMiQg7/osapcmi9RuZhcuQilRRjTqIthY6qzi+tQTsp/wiwhsZ0r9IX5Rj8bT87yDEVdy21
6vOZStn0gRf+54WHttKPqb/tph6wXUhLx+frCULPjg/qb/XsHQRJRgfSoGnvUoqFOy+qWvmOiyHV
kdCPKYEM8XLpU1buk46dLZHYCa6ca7Y3ZuE+ahPKzjffEAUGMsmVkLi0fziM2dqNLG7qWAWbKAUU
yNaGw1xQMsavYtobV8UJlKluR0fQp/G/K3+jYdJNcbQ1REiRdVwM1ARftkqbY1uY5kssY+5Auoq3
8ZwCp14uGnrkx0QwYMtWRliXq+2AgDQuS+iBb1AoZQlO4sEZ61TYEGo2K+ZS+0gvWKC2NWO0WLGV
2BSdvXPzzcxXs/a/HsYV4gutV0fdckiWYHLFrEZXfqvT3fIiKbeD2dKOrFXAWKYCJRY52MBe0iVs
jYo3gAP4zm9/qrCDH/FN4nVDJv+NM4l4JbE8XABHJ/XIobfkLSSiCERqKVQB53d2ItD7fJfJXX21
KDX7SZs1wUPFshLW3QsVswTn7D3GQtygiimhHqMk6RHEYZsY30orTmb2R1FpN4DbnQesrSl/HD4q
zyOBnKgZ3lK9i3Uo6rVYM/IY9WZcwK8LwSTvMQUuP5U+67l+rHDDiwmCFavdZJh8mUx6FGjTHDTc
YA1csfNtEBjqZV7v3tzkdwCxCEFjU5PmuY5rbV6G9wfZQpMk52nJdKZVmAzwftGvjXExTekdwPfO
odQ6SuoLW+Tpd+l0I2Sw7xDRgK8ip1EieLBmMtXjwrILmJ4jdCYSpGWSJFCWWn3ndqM2TLd1RXCG
yXSbk3ypbHtkezi8OHEBUvJPJ9jCzqjLUxWo5OWId/edeBeulTuqNJs20eWfrU9kcRwFrItpcSvF
UO9x3aBbbr7xEGGXbxOYJF6Bb9kcbcnQ1/7sn33XE+uDfErW+Jr80AjIg/o+en6q/8FBBUTcp5ei
7Q5brbDYb/MuzTtuiSXzNcM2kWf/H6P1ZKWEGEqf4IqS24kODHN2pn4iLaKrzP3ypEaPlkDrhChu
qUr8QZZ352aWlhxfL97smRbvMmpUz+amhR9eBgC5gcEOLJSu+75Cd7854L2I9/9qEZtlTnaY+FSt
Jbl/++6adimckzY6Z9q2+Hxb/l/74yGVOyxrZ5r9GPdEnMdKDm/OhsaiLGt6JhdcXlcZ/sbBS9v7
K7ze91s6izpUToXSQSESio+gqwNy+fqwMiGlPH4g7B+cLaFm/Y5VmdR8k3fyj1QoDSkNQzbU9rJE
Hf62/4k2fuOW4NG+LtTQI0rd33OQL9AGBoOU8ya0D2j9SEVEqgZZ1bGmbhUzGaiUWzvvftL5abXB
eMB9ggKDkN0m5Tg8sry2IYUMiLNnga5zjD+jj0FI9WozVHk3gvNrsyo+xkAbpiYQgYi9awyfpZFf
0ndNDw4cqlha1p+1/ia/VfiWB54w0zYUtZwiMod/IO5kY0+aAiSgTSKtEJ/ydzVXoZHtmikOoUi9
PoUWUMXteaHOWht65WbmxaoBdrt2x+jnkDWY/zxXsQNo/XRaxaACcml782KdxEu9/k82BHynd1hC
KAFoEhN44D7LHiwhaSV0AKZO/KcYvwvYSzvVIy7lzopknhFjaJiJxxR47pDmWUMC4ULThhMPXVT2
f2ETdLnyOPPntzsaPXY1ey+M3KYjeGU8onyOwPJ+ilqim4R5E0j4O4FiXuwGg0eJHPCMxdCWva+a
BwMu2PmNzyUM+ZjjrnjtBvGMNDTWEVE3NiJLDTSGSwdgLBFo7oS77AqhDzeMLJuot/Jng04maafj
ZgtSgPtvap0AtPKR2Md2kU6PcIOOTSA3MQsWLzrh0LD6eHlEySvK8BensFP+lVn+EG5PmBA6PsEM
jwakk/AvXPPQkqnW3kbscd0GkXDdlEBpzy1RhQB9j8RiaP39lA80IBeNmzVp7HFPI9S6k8B533gi
do2L6fMJ1D5DUXTS2Hsm19UofyxsiMGoOhwuIpkzz4gKu3S+HIgTv/3X0lCMTd0vAO3LZZWyC14d
FXLjHDC1OeytXAwelTvpUTE+nIFmRphTKdreCqO8fqnvL/hajlzPmYA+2iCRvimURvl1YZkslBIm
TFZ5RKcyUr+WFHGtoUOP68gulrh6uBMkLeLVNqn3JiVBdBnP2x4DnzaPocArU2pUXBVSyuxOrJTJ
ZhWrrhGWtyZMU/j+DAu9UL0Im1jqU0zS+RIU2ShcetNSEj2Nu7uvrB1QCEl7tY1Q5XHRm77Wte2R
RlGoy06acs1/gMvZTxFSyR84bY/baMF72DSJ81SgEx1D86SU1b8aPFw4BJyF60HSfwSF5++38wJv
E3F9ThN7t+e6Eu2Y98rlMjB7WTK8uMhgoVvfn69MfFm3tYWkjsWizfYeh8WNQ3ysHZiM0PWAJTND
q2JNE0QiJVRuGlu6T1XryDh9J5Jx8DLFgSFGMUb+T52SIsbmPk5n6KOnREiHDIU6XGQWODNxMw+P
MlXRp2nuo7TnkbjZoLhj4AV4tjxeX/Dkl28slyHF7LoPjQjRW4Byi6JH0yIPxtyZKhi2L7YPFPBO
j8uKTDKDffVe0XdWH85YumHk/JrClIGVewRc6BmihEU9LBFw6YWk1kJou5y6N+QfIltDHPIqXg2v
XAWJ8VyCbze/zxpEyu/0Jg4CHD4zte+8z9PKDnl/hSDapqhaSniLHV5kPtWM/liWoLGxOLSvZoML
YN7MKA2u/TzzZT4rectgCpOX9QaCG0Fnur0ywwicLmyZgBUHA6rIhgesaqYQML/B2EOiUUOS5xQX
/O9U/Fy2flE5CwY0xkVbqikE+IpayN2DSATMt1cL/7zSZ6Zi4pXn4cTdJBHjRSfiUqukI1PcqmUf
ophwcjxo5BKCXfHyw/GYYpIHFBcxzT9f5UnqTB98dmhulujQ87qIRKFxqs/ZeOjgVobdUNe4gBgb
+v1SJZ45AxqjWQsjczkxn66wswWHnx3BZrDW/BTMjUnc/vj58x7BlejZ1BIGArNDLIR7thhfWOeC
WItKRXotgMOk/PKHBalQpIQ2fEXubNqiIqN2CaZhzWFftxRHTWwc2J6fRf/k9ooERNfNp9AfToQb
0ioQ4vNxjYSauurqCTYBbz+1e8pR9LfLTrYRe518rZIkr6PKVRqPsN500i8sCZLvabNFYAztJMrW
JMfyYn4JMpjUbldRlW4+UNAO8nIi4SY+yQ0Nm46VQk551CatRelY9J0lysvKm1sesrNFvklDoOce
9l5ALkzyPgmqidhYJTydn+51/LK/j0OPwHaHeqOZxowrTOO1YTpvXc3q3SK4dftznLDBF4+U7bGO
k6Bpe5RzVkSV6DU3AbJ6+G1FlNbDGzVcgi8yr/1PGX3qnNhy482peXoIP5CpVoxaSovTOJUUFtq7
O9i8N3kuPw3ebs6AX/ACOJV9Nx/SyyqS5ty3UmX+mbqx8iOrZUSpr91VBVHybgwjx3fQRI55RmV/
lwkNSVqEG+jOP/0HS3oF0aKZZZBLaqeXsRaVtOTA91Yv2QcKO0sLF468THFR20h5lkKMyjLPsoB3
SnnmF+DQ31SWPV1LGvPVgRAwLpvd5/056KqElf3NRMvbHnVPncA3Mxth+WbaQ/Ys2jqNSKxbXLn/
QZknWE2ACeXzil2VchsV+/5zPlfzf5NC/NaCKBIAV/xbwXZFcdcNykQSfH4Lb8l0cwgD9RHjcS83
HHHPe77JqIxORUxXP97j5YDfbqQtNutn0j+rsJxG5IA1vpQQLIX8Dk8HhSMnbdqsnAeA9ZGRqgDb
dSQy0AQXj1T9wXCgiHbkMB7j5nnHGY9scxAAiDjP9rUh8BTN+kFk3AVHIp5w9t43hqb7f8gUjGo8
PVQBakyOxpZ8ZZLkNaF+iWTGj0Wly9HWOfwh5k4AkaV9sLoqvaduyHIz6QhrsKqrorYoqBoliWP4
AX8MU1wtIvFfnxj353SeaTYS+yt4ebYiZ4RGBlwQqiABDuvWGwHPpK2la/PLa0y6WgfJ/uxMSwu7
dIR5Sb1Hf8K/Fx628+e8VQJ2I/f8GNldfvgUfEVqhf40rOcZvMORBkzrGqycEGeeRpq6GpEdCyf1
hudbywMPt4S/tkzzOWTS0yX12Vp0IIlXau0TPABastCf0/T6a748Msemr8/xXH7SwsnDYW7kPvh6
glWMNo/B/eP+Kr5v+Ceo5hEAooX9zco2MNzPAil334LQhzw0csZAFqQx8glfR4GH6RlD1BDqIQog
6oHVuSEw6f+51Ftsk4JhjlH4rtA+wPBcegQFZ6HnnlJEuZMwAtj1s5CKqartgifvHQqca0Z1TSRx
KrvXey9imuH8wbu2rJNL4DTJ3yOtFjukIrII77uHM28ovtREFevtId4bsmuZm6dPXI45bbnnCaqo
m/TilcsL3raVuA0WI2DFKHb5umayV9Bcl0U2GpJxk+6bzvnatwImEvHZ5M0EyYaKBaRcQ5ayTYab
KxQ5SZ2pdglgV/+/rOuaYjfohhQViwCLJLqq6U53o7VVjI9oTrrx7rmtM+g+s/Cghc7R2xcCWfwx
fSXnSrNxQt8TxkXBw9KkvYgvKGeZpOzsfM0twVMaBKxP2qx802cdF0iMlZk8e0nGPdzMbrO/OhUr
P7r5zKolsasTBFMLf7zduC1MZKnEqH2mEQnouepU5SpC578zqMM9HMfh3l+tydkl09L/vS+0ccqo
bpV+Hlg5buM27nibZD18vhlIhl47KOqdkbSUKLrmU4yQNEDEwB7+dkrN55VAHg+DhN8JbeL1I50I
szyK7mEjro7OAM19D4MBd+Fh+UOydfraqfEXQhsDJpCoceH+qRxKdnlRCCmDtgWDCgsjDc6GL++g
gBhqqPzfT8FtjQsLK4EbcaxuoO9UVv7jSItiZTltPwcuenTyrTKF0+jdewnWas2e1ZWyUsxmaCg5
ChJdBQmUfPmbfp+HWgc3N90bnecnUXpCdnDBncEtE3Y1VWbkDb0vRHjJnz3SQdILmIrAJolPlLJU
JTTBZfkwkNBJpx6R7ZNrjHxP8pAi/ycq/BtoZB/ujlJ/B9LtzKlpYzXji7XP0JSPPPi+i/59/ASv
MDonGHPTg9Ym+oZcTl+Mdk8SnHccN9zi54Q7YZu5w4C3c1Bk4ZzFQiPxmwUJEEtdy6BkjLvVc70S
88uKA2jW9iDTFhpImnoLcqCZuBN7ht9lJ4lEMlSScICJtGeSayq8+FfZVcmKMtPbbsMh2T43oYom
1oYpBg5kxBmDIRcad9Jjdv7wt037a7r+Q9eXqTpMZKDt72F7MhJFB/jmIit8PZnkKeVGmZgWSrsB
USKd+/ETu+MMQCP51v6hS/BFZ43/xS1saa4nfBszpEgIh2uSFo5bWbttHiII79jPUJ2/FNADGX9f
8TP3ovUz2ut+8QLAzAVWykRcasih89yKLl2qQUf7F/Rxf4fUoP1B3vUC+8iJDcSfhxYvaGLiAIRR
/hU7Z4qOSzQKVVNJ5NFKKcIQZHeShP3XFU4f2iOrYePTpBQXyrY/z6SdZgrW2UKWWxRP7dY0XmID
d8r/ZjPE+QLr21g6S+TjhSLQguKAmYCsUJ0uLAbug9McyxZNX1XxwDZTAR1Q3EMfQDRN7EZJoTfN
NbhDPSd9PAKx50RQtFoKpkETGWKTxvC+gaoWNo4mJUerNTK+iI8rAvWiB3Pm388KG45rfsJTtC8Z
YfRGn3ZldImpL06ZoRYzA2RbLiKyAb/Bb5E5RvhLyUvhx36z+Tb7lablrVk+sILpQegTnZePTPWq
yTUxtYWQ4ZxoRELHHIU1Ba/Nl22Nt893tkO4dTVMv+MiDn/7biZsCiP+RjlyMtXuw0sOnkFO/j0X
aykBiL11Rlxs0GI74wX7QoCKLh1h9Fsox1DImI9xhuQXJnY3CgnweBjsNs6RxLU80HevDM4j3oVi
bsXfz1mC8Ovqp/8daSbBA7voLnM3xQF/DB+OpyXIGXyd8iXBMYss1AF7Kh4A5ZlgKAE8I/tymc79
7ZQq8Gb9Bv1DABlKLODpcdbMJhPQ0OW6C3gxfokkMo2U/lJokKSgaUDEQ3Vt1DeE0Swlz1YB6G6o
TgFGPEXpj9awdb0EdFeQTx0kOGlbOa+ycqzb1lvzDM6uNd6t5YtgdvKKMPaMNIfg3aj584kBolfj
xSEwTkWtmTp4MEQAw4Adcg/dFsuE7beO+30NK793SLxlRBYIf3DT4NVqpPPVUXkbrJDwx0F4kQvW
0ZxFYVPVHQZWX0fCZ/j9pNxy0sbqsx4E2P0smGkZq/DCusiQtYxWLQ7zKYmK3b5QqA7434XPTHMH
KTvRsgeI/mg0EHA2+8wNX1GJiihx8tNPQ0kM2xKvTu56xg4pIVINUPemNrcGdIBGwTLqu2C6m+nT
A+z66+h+bNH5WfKhwuVnL7zHajhKlOxOI7hmWk+GxlE6e8TTdHXg10rZOy+bMM+o5dO0Vv6MpMII
r7CZ1i1uBzSVc6D3h99iobl8/N9l5SPxPPkUiWFa4OF+TmRlmfFmE42tYNLiStq3H+XXCANMs/zY
ChsbqjcLe9EqYZ/uF9NuTHScA8FRbHf0og0jXDzXFwbZg7KzTgOv5kU014oQAZRHIBM57jzW2X6Q
uiZPHrq8J5qKU7aiI2RYJgB/Y1+O1TpeBO8FIiB9DfC78YyAYKSqSvJC++8yHvUnDxrXaOLa8A8P
UzlmwL86PFf+NLTo2e4x/sHoM9EQIQE6cJA7uH2Oe3p9Ck1bzEpyzF/Bt/ahThbeCIKD0Xp1gPxd
FQ6ss6o1iUYcF/ohZ6DgXVvKKvizA+4jdkSGIvFL9xixsDYBwj3tJr/D00AuxrRKmTyYcwyFOjqT
wFF5F/aPZvxPxLloOoXrKzKf3CULdMFDogq+7rTYJpN7sCIQt0FYKVPELENWBK/TEFSvllllaPD8
8oeUMDwohd3viNNqPXLx5aid7uf3s1xGX9jUqJrcEHpX3U/HV5UMSBpRCwun+7ArqqPIuOfcw4sY
EpSy88EGkus4/3dAHPvkGY7U2wKaYIz4uL4ma0zDooHRTqZ2tFtkhuOBE6l7LjF496NgoRwlpt9j
BNdxSHbQ/nIvaNOv6Bk33fFFNb+jEmjMMRaqKIW6B+q7P08PQT/HZAvTfWD36nKxofdhWxhAWxnk
XWZK6WQK7H3MNvQQfgzI7yJ5M3Q2Ra2cI5GWQSGTOYHOo7nk7MlGlrEnAbnf4GamDpxy72bmFiXP
yaIiaxS2mzgCrentT7q14G4Tez408mT2rqA43cqIWl3WjnlBY+JlHQaltvnkxq0O7bTOQ4Kcmaba
bWST2pGpb15xL71YNX/ePDRxNIF+DRq6RLZmZNQNHZ+SI7gYjwfMHJLpxsKd6k/uC2SPmcx5xw9B
+ylPqnUuJyNTCRW6APaseoAMD9CcXc/j9wI2xV4cE6f9d5kVolYTp8M/azqudAdxKtUFAKhHeT6O
kAUVQeoB713O5xJGdFWwZYxZoFIsqlHlODnatlX4oExnecr0NCE4rCjjelXgzviasz4Hw4snoixP
TYcnoMBfVLDkTS4ICUujehanPBnIdBXvQVgoLiQ/h9UF/d2hP+BfWrir1qmvj35JXoaQXmWmjhTx
8JEXBoJfW9PKARDfXEeoRCSNdR78cZeeciuVZmdcAeQb6tNkthcXu15fDvvJmFLwnIj3lUb6+KUe
/qu7Ht6LgYXHY4JMOehN1NzjGcZr9gR/ZLgSdIDLplrlCsK04X7zRmjYuUtqjvlvXxXRnJV3mURY
WpkYcZdagPy77jk6zAoCtOTzXCELVaJT9/1UOAXRxcFIdGHqyTn9Ru6GF5B43F8R9sMDGzgCfZVf
eUd46mIEfJ47VxS5DRVIoT9W4AECH1J/fcWHUYjw+LwqeSSWEbgHjdc+RLd+amVaBxJj9IkF9nx/
P7jmKe44HhMh0+N51sNCTYMEHnPPqwIzguT2VOOektxbYk+4HIahR+Rle5hJdGGZEiRKJpt5eVBD
V6nrCm6j3w95Fgo/SkXk1dEwiWGBTR+Re+01qIhgwcMcDbYdxMYJPcnxxWDJPJGkn4i6YiKNvrlI
F6/9uPWbfIm9JMODsIyjPLL6IfjTb0Df9gv8gC8/oDWmawjdxeJmLMJLiShYvwEkj1gbCb2J4OXe
jOh2vbNE4PVonLum6nMsi3edCt5QZ9CFvgw0y7JiRoKDChySthU7E/LH+CadS6bF7ecNmkRC9lRs
G4yhF9OSDSXa/ryke9TIuDvyKKRPMQWH783HRb7hrxR8sVAlnN8G0cjJcL4Q5JnxB9wG5oWEPTKO
O4sqXWAXXJ6RY0vvOR7IcV5mpbZTsCCUHdzyX5AjYZwT20SpE25wMArhmDQfHgl/H+CPhnMkVnCS
6U4srEnDfvCxhfSYGyQnpNIr9SOr21bleidwcETz/NbuGnAHYKRHJbrW3mkIjhXERtCpvujvczZI
zx/CHshOuHvAvq0CVtj0j9OpwDii4K5sgza2GwEZ2ZOthCbYCfwQ61iD6capCrgcREOoEDJuNXKM
u8Dac3t7+owRf5Fh6zSuUhIevUfKGV6UXb9gqBhTn5DZzZA0DtGom1HgDKGMf4afLSwyLvSrJuCi
h1xNmGdM6ssLjHNPb9fNdrYnGfvk7IYDoaoQndV1ghK6L2KluxZD89/xky62VbWbXjpz6RzHe/Kx
kybhxTCL2PueTLo6u62D2BdEhEsWkRyX85MzqwitG43qD42pVLBCIAseNogiXeZcAOdaYtnw3Ogk
IWSIPtEq2oCVOw8mBsuwzdOoDQJHMhcyxR0HELaG26Eq8M/Tc88I9WXr44V9/tar0sjaLPl6TUFj
WqcUiMqS6pwBu03GDs+TTXiuihDaVA/ZYYjK8+KDdE+dMP+etdkI6qpVcTdheUGxq52C6J0FwHK9
JU60NexekhRyxMK7WdRbA98Y3Fmn6mgMbQY9kLznjbLPddUwa19IFhzYIoQXzu2vUj2Tu21VZjDV
+LU5iQ2RB2Rxr7dY8odM08nO/SAtC8+Cn2aVFxqJnyXJ7RcvytVs14Z1mgK1rtMtjE09OqeJQID8
DWy1ZPDUCfrMJZjQ7AXvXlMcV5ZJyvLdZUZ83K4+HVpNEuM+k39mz4sb+Cguo3GnYZqfAUO/Rsd1
UvfLNh6MM1Ul1Rm+KuCjEGZieSvKAktPfCPD+ncN5e4JOKqFOSL0iu/xEpjaGaYX0IhvvYnlD+dW
0gkfaQnGdlH/i9IgkObObKI59OnF5jax6+q8+653kbhTkoV0vQaQxtuZdeTq9vtOHP9ORyAD2+hS
1egtNEG1fs7xoZic6GwgP1Qq6f+GUu7/MVGQi7I3EGo/Q8uzN8YxCIL7mx1cVa7lwK/GqOxqX17c
0Q2wHxc43UtLjjBqdagESumIZP8Dda2NE99MzhPsFaRkkMx04E9I8kvb1T2shivwfgrfohEyXcLy
4+oedmvuQ3wnrGFbzMq/VbA+ET/5dF5DjLCbhRIGaMyUjSV96IF/ckzU6gl1qnTHVrxlurKvS+Gb
0lwPt2HejMW54/1PEJagrSF0bnhbpGvx9yq3JImato6SIj4PwRV1P88MG/SaL5TAu6tUs6gWJWOi
6AnvTcIcBMYna4rnFv1e5t1ap7DxMbNsOfkd23R+HhxctmPUz02lKB1G2GjFl9QZk6nwVeez0+wi
ke/Q2hA6IZFNc6IuWd31+nebcPh1cyov0It0lOg/InHmaon+psGbA+Y3HJWq1YdwAmatHa0tG9GN
qdM9i1eY1HUgnTlvJhxeGr5Mu2wDIiWAMtH9XeE7bIa4Jh5iWS886/sIHdUAPpAClj9fgT/qPXdC
a65+VDEB1NC+oTDTcgpuNIyTA3Up4iC2jD4BEOKmZxTmh3iohOFAmbhAnh75VhFJCa4a3AfE3duL
YEVrN/mf+3SnvQbzoRgv3qyuNCoTDfBRVzvrqDnk78JaMh2OuzWMetbEEN9QYczgg2kH4MQy15iS
OY8Ds9A5aBdoakN31oF7wYpjeWckitGz0nTzignps5BzKe2W2T8Mvo0ObTiPpbsVRXMei7erax6z
ZDMAEJKjpdL1ejdcEP224udJeP1/PXjBd/vWlD7QWr5FryPFcyaR+Bm2OwPjxTZVlYfYFfWkQwD1
XQfS63CyXGDrENuK9JDUp9V5d6ULjZTGk7X6csiggXik9oR14fvy/5UCri5nnpqGanfhrytgoS8C
iV5zRCA0WC9u6zf5CAhurRsMq/sxKMwzx7w8a5zVqhCAFeXCgH3Re0M3d1LBtHd37L8SLETIsxFz
lKtLBDXEX8Vph8N00WHY/zNSmOjyzyNNAxoDVuJhrwqnu0wPkmpEuHNBPwYpaJ/PmKQtQ9j9+fHz
TZQgDQLUo9cTs0D6hJ094dKAF1BkcbOHV6/WkVH3HDSAXsfDc9WPCnm8SUrmN0RTgNLOde3+CJEz
f6LYjqkRylHjajNfrcq81zKfUgXW1Jtnuy6ZZKacAs+pvJQBvb/BvJlrCd5zr/MUhBWsj7xBW8SO
bbDLHTPCitQRfyKJX3dEDA4nczv7OabMW/1mJPAKbw+wix6RyIEpUObUjyata1ofzN20O6arh2mQ
we9NMGR4/RQx3o/7k3VXG0c1ODE2eewNA5Z7JRmCjMJsqdfEy79Qz0f2OQ+geof+2DqP89oeJlb9
Uam8zz+NvvFk8+zgZwlUYl3N6PQNEmFBAQ5z5ta70sVBN+cspkDE6PiP5lQNo9toBqEuQGUqxH1n
Ijl8f6+7LcjXGLvs4Vdykl9iyjV6MA+SQprbqXND/7MTscdE0hbjFWGNx9fb88cmehbX5LnOaAIe
Pn+55/OfcNIYEE8ZLGgPI7mKLiulDOR2W+qyJLoj/o1UHP0Cp9DMcGJP9E0HTZUEayXFAAZB9g/e
0ZNjgRVbrxoPYlZikixg4B1NLU7EQ8IwH2p1AeTywknp0xEMyeRmnPcTC9qL3ke/ra2YNc/6Nbj0
RTU1kGOvrip+yG/+9c39Wi3jT9Bsw4r5H0qjQmRGhYnbmhAoA3MYPSqJFs73LkTr2lTzmeAli/8/
EK8h1GDTvdDdAhilRiA24wohPYvvFXAyH+oH88Lhsee9jxjyJBYixypXBgZvBH+CPpYP7bdNCS3E
siItngAU8qWuC6RFoVvoqfOflNWLX/z7iJB08vdp1yAYOKrd6ggvYFn+ZEqnBBXNWxovLdvnyHL/
+qGv56PPt79wG4emt5gOKsAH0pzx13iuD1YjvsKePkDLiwFfEavPI+HjsukCW8Q8QaLhLk5M8Dgs
bP8sxaFu6uK1xDqLWD5i25CPbiBcONxYh4TyNL4SjCdlz28YZ1CChvoZdFuGHjTzJGNu7599cCjp
sFDOP+M51tFzBQOnNdFEiiJI9VGEyMUE0KtmaQ4N/OKZUTOW3AorDOCS+yfx6rv8R4x3d8Jjt79T
bLibNk6SSs6U5W/oscH6sSPNC88HE89MMwW8qiGVkvWM6RogQoe8tXm4hoX2V+shoI/Wklslz5FK
elOThDOlYuqekely6Q6FLf0FmVyoy3v5YooWFbabW9O5O97/EYbFb9UB7IboF5rPdopoZUgMBori
p0MEM8TfGPk6y+YiL2u/6s/v1WEp82psIvcjE6voWJHl01jIH3jVWO1nqgtYQcUHb9UlRPTd98Ls
YqDsZ0V6CQqgTIvM62dqVbe7l9jX2JaW5lWzorWUBvWqgkBHl1NOjDFHDzZthsKXWGvPdskfjtbK
QrcjMSI4RU265Nv4MREjopmrZwmCMPS/ea1Msu6NVQeNh6ALLSFY1EkOhvIcx6L1PMnANGbb/nVm
EzlDV6Hde1zT93IZc5m3wlV0agTE7Mth6UUuOlIkIllgl0q7GJ0XzWOQ7ELx99lKkMd6f5Xkc/1C
+4jJrfkCEjTBwALTP2ygI8gSbwcbFF8bBvITpK0I8c/bwAgufCOhVMytIr2q9DgTEz9SnFPjcAEu
nm8ITB30Pxzkf/cxtGZQli6ck+bjejPJe6b/uFvfYVuPR21WPtd9ndBqMtYNnNlDm7K9WqPQYaUG
twKUX/ng6Vsp4VHTP96xlJGz2PPwN9Pvvfo//Td1ltpzey4DGTSskfSe8ET5a7i/ap+8SPNN8fEm
wy4BB664IRDYKcYbC2Lmo1yfXZ47ALE2uLuu4vmlP27h5pqD9aOGX1qjBsI9jfeA2EkhwNWZlSAP
WIp219Ouzg0T+yucF/w9BBMAxnZKBwRxCY0mIeyzs5Rc4FENCIZRiq6/40cI4uKYIbl4/RaWCaFh
t/2Gk+4tEKo02FuJ5YR6sV8ab7+NR43ndRhzC+yVTEsabKJ54GT/fkPM3jsPQLWkiEJHqq8/e1Ul
lgcd78HJ30HzD9kXX4ViHcOALk9gvzKaKMPuLISKWiT7HEZvZ31uASIM6pbgl52DLGbZRkMf0Wi+
fTT1cI7W+IaOmqjmi4/syVRpexwIiFcsqkXdoSRhRn7P/djRZAmSNmaJkjHybCEeF11gQpJghnCt
Utl2DoSZA/Z/CkkKGAqoHxGLBDfDcIMbU+G4tvM6lZjIOj7rLlLal2HvopNsnhKYPTah6DKk2WAQ
FQ497vR4d2b9HsmJBo5O/PWbps6OVX/5EeKXvuZRQKaInPTRo3i2ululSPIakCPVJg5FTH+fCxhz
TALqM5eAZK02cWLM3eRODj02xPYFxGPZwFrahxSjMUdKDf5GG/Gw42Fgxy2er1v+LgvXkmPMUUPs
CCfOyRfL7SiQ5QsxrZJ2el7oB9XxSCovwPJLtemoY8G8TWzQOI2cmUd0H3ILObXGIZSZvAepmyYk
E1koqG9T+Am2+6SjUh4YXzyhKDYtZlD0rQqEv+ZVBG/f7IS639rCkYGPWG3kHEirZG+nBItf6WAo
UUiinuNaPnd4j3p1SZtTeVIsWyH+UReDoFgyMtp9vezgOLOioHwFwY5fKLXFbgLoSDl46Uymz6hD
O3d9FF7GtdvstmGwHd+TOrrTH6ct7N6RauhwVEXZnxjToKsAs5wtao/UnK8KXlYK3sTsgsHa9Oea
yzSF0e01iQVNNSTud6umw09R5mvHIIGpL97mYncRLd28eoWBm3+JgiDpzl84zMIzixeWNR76qT85
WJHKLUTrdVq3Q/V4ucRxyrnsOB4hUWLM0TTYHxcPmzNRZEGfbvs9GGcWM7DoBSvKVKZk4OOgEjXm
Us8z4E2ZOyEY6CMeSkmlkRKIMujQLMibHE1YljZlw02FJpYVkbvl/Oswt+MlWPOWaw4uzBaaIZzV
oWNf79ONQap1NySkywZdLiv+zqwfm/7Gsqe0HOuWxJULo6Z6LRFiYp5nmxrfuOhsFCdeunk6l/5G
3ICe9K6lxNoqihYYaOxh4r+5h28Tlb4p4C/ki6f/SX6rB4GpdkYkHkkkJBWtnB47o2l6/eMNi4P7
JsC/hJDf+/s7iMWHuE4wl0mQJDQLZLC+CO+fis83MKTcznHmiOIstMUzWtcj1fdI9g58zKC2P5XB
UhujXwmdQY7Zre7u9THT+zYVNRyJksUB3tmVyq+tx1Cvdk/Kcqf+bTTEEar7umJ91wVm5jIsjWkw
EhotNLQl8vxvOACL4hSBZNUz2OLUn9uyZz0CvQy5UzCr7VD4X/wcVeJDGZZOjw+Iy6Ord68ZSylQ
I1Soztubw2VMbHmjMS0Dr0PK1CDo3xSYZ7i+6I/9Dxk8mPLtd9Vj23JORGxfVkJ71pKA0WN2GPLT
8Zl3tboDbPgabpEBWv+hH6lS/gAkULdGbh07FgAmYMZ97x4zPOCRisdV0rNaID1vgVeFEf2HWw4H
RQroxFrrlJFq+CLHekxYpq85DDT78jZl0WxA1z+hshhd2ROWjCvqB1b78a+XLMMNRu/CWhQtxRM8
+IuF8tsiae8W0g0Vi4Xn8ocQQXl0iFTALIWnUTO2FTfAkTJHvUdKIc/4pU9Mc0XHeErQOBMyqhwf
HPx4tZd7YvOOH1skItwq1wgC9bA4PBgScExH0LQMg6BNnjvkosHhF/o7/5Fvd3c5K4NPyK4lNlD/
8KDgniG7BvMkcPyrqfGmo5kqsyeuOorWsiGrp7b+DTJGuGLY0Ffs7L2tMnLPT16NP7ozmxWuZ4Y3
KtibYrG9bEXEiIrqdTaIFbyhs+OMAkDH38YpPUuF9kz2E+SfUioxsWHFqTwVz7MnWXaaeC8M1oEC
gyjAwwcVXnng0ypwDeWWpgV4LExX6LVquJymzX6UghKZtNY9AyMVU5e24ikkvgy5ZWNITJsmn+qv
ak2jT5Z9oFWwh8DdpjMolEe9J0hTrGTeVVLN8F4+ujFgLS4B/iohVBD4RqFHKuJT7QDqi3hc1oJF
WKwuW/+xsN1dLAKZZl6a3rAXRKhNm5StiO7wf7ewlJ8c/86ARbipDlL4yGNS1XYDIvMpDqKdasDY
pWjT5YRWPhm4tVw+Qxk7glnrt2d9Z8tqYmsG3GUeHKvrKFwCd0ctgClVH6szg7OYEOZAkudaaSmk
FHWf2ijLOlFD7/5dsJtTpvFqKERyHZT1E8g7MR6f8mXV4xjYAW2oxDfQsUEqGKJ0dZhd+lvlninm
xlEU4DkJNegQVrZmEqQxbFgxxmJEL4LxJltwSx4KNo/DDYPve0Jpe5jbLBJ4VA0iYZ6+2BJRiX2B
O65x71FK9sEe0EtkSmMAG3/rNqoaO5clvvXZIpEyFFXBE9qpcKqimtFmSCWsycKLJ0/uIGnzIPBZ
il80EZXVvm/akQ1zjVNayABG9iZtnlnTIoUgHGTku2hpLUHHcjgZnDoqcPGw9mvTfFGJNju+QvwZ
IcZowMhhCwn4cxL1U02/fwvPG58or2ENgZ6BIOHdo2XNqRlcEArPcY2ndqjiJquZ8jYiP4TJm/ZR
e8N/yiBncvHUhOuw13TFnu1pcPsdHTqE8Rl3Q+A+UvCkjSE+NqDAFDR1wxFVR6sDNJVfFh0PfEQn
sR9HYpg7ZWYE88zxFMRXltK4jlqVAgXK4hzoy5rfJWNl5Ds35NTpYkug1/OCHVX9xS691Pu323V1
euC26zxFuB4OY2pl/rL6OIlqb53+GKFsGa0fUw69MgUW1xH/F5DiMXvKVwIyI6AR1qkWgR6dDS5O
yMh0KRBsyjmEui3FfFZjShXRdmqdRwPaRfE2wbXp5cMTerFWJl5wPcEPYLOoSd19rjKmKKBBRtsw
wYlfu/YuD2xk6ncoM0I5GKXFIDfbGKdPmRtYxFSXNHCR+fmti/plhCdy6bFmKKfZugV5SMrNaH+w
zgipCV6YYmZBFSNFaqfTJ3YQwdh/ZZWH9F4A8fnBI7Wus5DxVkjBPicbOHK5xlx5PMLB0JWtFp9i
1qU0Y6FyTOL83CMg6jlLo16hUNzJk1T6UI/wP7pAAo1di0QThOONm0S90Re5Du57SvFdyON3yJNr
h3jmU5gP47gVL+y9Lm/rbC0Q9lkte8q8bQUOauM934liJU5eLMWDU1qBQdRgbkOk3Iw2GTJpiPO6
vEBWNRzyutik7F7V/BAXQ4W3VKXq+jB9m/zzmy/kMZMjmISeHUzSBr+3kblSHbR+k6cD8xmgnvZy
+Cnixby/rTuQC1Y9YwKNICCElKtqBT9NBdZ2p/imt00WEJXiEAwO73aFqy2hpNOnVRkw5advbqm3
YixaNgScwmmsCgpwYPfif57YWD4W/M92uXf8nHe74hcmfVX9HusMnqxXEXCl+qjl6G/5sjCEToHs
DqUgcpeuet7Ge81AfaB6SNnfqSYzsY8KjsIvZUK47tIGZMInODlbAPXdHH6jVwkrpRG/dYsGRsLa
5dmYWBeJFnFsCTcv+NcBvs2Pu1BjBi/HmtaYNcQQ++lX/tQwG7EUHOEVdgIX/JvpCTjHK6q/uoKC
AtzD6Q5DyhLh6kBFUNb9+Dg9hAoDgULEuSxJ4lb9QIhuZ4qm5ANykYCqyeY0/zqorFcTA/QMmimA
xXkPqTv3cbxU0lzPwakmPBCVzHFVYoqwjhO/ZXUiDHVRN9ptabTnfJ3j8vpjpYz/2LRnArJhRqtF
IknnPJOrMeAfm1pJrFEOhPZEKYGfdIXdGSSgi+8qpw4mLc5L8J/rQTIZigXcqSCm+mTtgA4y3UjD
cWgbdvGptUPsFybrp8FnWmsXiBaggmIMRIjeXerOMdusm1RJKtqIZ76YUnUi+q0pX4naqyXYKnFG
ujOEzFhOGH4tbl+EHOq+iqCS5YovMvHE4MyUFYMh7T8ApFhXOIueMDKQ1MPDgiEVyUrn4Q13Rync
QjIIplyyGF9wLrhwTfybNvwrNfz+4H78zieNXdX/ufsyqZqN6WbhEdJf7oC96l1sgrHfAtrsfM6q
X+VUGD8qstBGI5BG6dBQVfflvZQtDlSJkzwF/UbqtcJocFrBa98Xs81jE95xcEKDyDrINYfrMhOQ
QgbbiQiEB9ZrzpK/CE5AqycYg/YRg5N4SJ9TN1wsXmq3axASz+s9jM1FtDxV23zYk/+hYaTCxBxk
8hstJMk9uX6B+SsuBQsRYNV6UYwNCSE2IkQ60CXo4iCRgSGc76CD5pThJxEtK0POdjRac0K5CscI
Tozj3IVWR1U/sT8bP8u4XaIhU1ESB9kkzUf7s4Zglhdr05nwiL3qtbA44EptlGuHpJwW0msLFJUE
iSjLwOyANv66h7yDjyrvLAZzXji9OtIBXBRwyJgm1dQ2i+6yMZ44/jU7qRRY5FRS/sCHFcJMrAPN
vtaiJnx1WAPr941pk5tn61tSB6NNvWpAgDWfdDSZR5v3aArAcHtO0ZYq25isoLP+gCPMBaiVvBpS
pfDm5LWPGWI1Z2u4qX98wvOj1507ScF1Pz7wqGR8CI05VRYI3uT80wwTVT9fdgeAIGpf62mr8fty
8tahzymnSzzXxLWiid1PhY1dFVnooUKNqdaCg9AEROV66rmkxh7VsSnFhlWoQVbqT42+ORc0QkuS
lF/7Vi+MyRDPEqzjERqovyP/lZPcSIZ2EbAWBYcmQhQDQYULP4TjTp5coed5KC5GatPabz1PIIs4
Un/8qi9BYIgX14DX8PRL278sZRMYNyPt7v1oh7+8ezBDdYSy9T1HcAkuw22cZbeZ3bKEqp5xzXis
e5FNbY4PakM+1CjAd9TnF5lQA/8tI97l7yiCZ7FDC8JC5dRajXm/hA5DCSACeplvmfgQuZRB6NWx
qpuN+5LLC7+SrcRiGt17LYFmiIa4ZYqI5C0TKRLY7x2z3MFD58xZIAilQRQ/vAwlTTt8hjvsXBta
EUsg9OxLvN/sbt2GpC8Y5BQV5uZntrgFnUPAxR9IZnGON0WnN+yoLaA2yR8sGAf0FyFHwyRXFCVd
3U7TXJSWgQ1PCFPR3YihN5vdHXK44xO4QtKt74hBPWLIHdB6nU8Lz976Fn/Ev+3BlIVmZ3dvjARG
rJxhTQyey1wVlMnULjVgEkvTIJ61KsyVNL693QJwFYxaQQamg1bZCyA9kCdUWkDl8KMTECoWYoys
FNCSHelKyKFAEZ8Co8oiqcf9bo5uK2E7ypMJExSUcCJOlrY29O21fEOxAF6hnhVoEjP/ATjcRPst
Z8eS2M/5BDEHP3S99y5B2npjFvUTn2gbX9O1by3i8QtfeEx2ex6ZumgYqt7IBbG+TFZU3BXwlnwV
2qCnkxP+ePhglIX9RhcBOJF2xK7sV/msHf30jn1armYwoPVaMoc4Zeh0AU3fDbtPUc93+nMeCPRY
N2ikrhRp3YhEos9AIJIjh2sPRz/or8yhGAn8L6G9qtctKgOoX/3AzqwCW470XcM3nM6phbY3t+3n
COiNJzk4WKOi5FgguGrnfSvv45VOWSFJSafzVeItF0EAzhDljN2h18yy9kMdxcsqZTCPq8+oa0wV
yNh7HvURq/7lnwBSpOkTiV1NlsIwcxSmo0KAjqNL2KyTXDV9C2+WTTD2KMkS2ZdqryR/1Eb1u7en
3L0tqR7y4pJjGooAM2VGAfXD/8Sl9RF+k2DPuWP33yzjdTzO/G3zOGP7wyYZ7UGG/lnRmo+TNm0l
/6wXrE4JlWnlZQ+QFNQ9ZAXzpVMCK04/o0Z0S5rvcZdKW4SQX363Z+TQiGo6aB1jfoIvP9ZBufvB
Dvj0osAfvkr7pXgfKK79paE8bD6i9/XOBcSrhxzg32h6HuqEnXq0m6dzTUOZrglN1G2vdbvrRM5B
cnNsPnfvuOFRRAP4CeHnVZoQTxr9Bq+CuSerrGzGbWFHaXByRG/WoxOcuQiOP/eVJVYSw+MWObAS
PI5dTkbtiDCS9M3wtGASKgV8cjeIgOF7nj0uElOfamAilWNcMe/F7D3B7KnsLi9vbCc4xhg5JP/b
lQ50DXyE3zLV9Ps+ALuf82LvcQFz7Enreq1/QvzWYRUFp72Ar27SeYgdkSShWeeinQG0AoMNC/1T
+IExGSsC3tRJi8/uAU6e9LzTqmVpT6QOK+2JiLD/05hM+cNjhs0/E2aAJmqdsnJCjY4NOJrHMNeV
VH6JpBrZdUIT1bR9/7HS/3Fm52HBxbURWTBEa3V7y/Ez9E3IpsaI25wR0pdJEOVvyKzZnDkUguTH
05i8v0br2TTU3lG+LflU/wcKTGSttBKs9KQkaxFJOuWN6r8y4BY2twMEow7vu+kOj438DQz+4Py7
iEOvipkp2drfvuwiyLNtHwlcDHNtgJ5raqsXXz4rYf+uhUGHFXsu44b/CPH5ar8KNYEl0L4Torw3
GNftWWkA8n9O9eEkHHHHn94KqW+hku2Tmu1J0Z66eKDU32hYA2LCoiotcQhAG2fbMpn+KJmRVUQz
/I82qvd436Q1KgfTVVVyEfZvj4D7yJoIda7KBVJurQDYDmN43HCaKnKkh09QTTeZ/3I0ot1HI2Ic
0nXUJeAs5Zlynr5nJIQTuX7Oo8GJmxrrgkyWumvSBy+gI82ept6qgjzoQ9IttnL0vTQcjeyuYhI3
isrFws46XGMcj5vMC6WXDtp9STukujSakh+pDj+KsURxkDjbx24nTAx7YX1BnZ8znSrBiPhnZisz
pervUyhMF1DkqB114ZHR+xrnXKp6cUwS1iDpAkB4xdn0UzUeX1DUeLX+tcEtyRfF9xr3j3Fs064E
L1Gwomqe7MRqEZB6/8VOpnb/3hvgUAEsQyI3JqrJ8LRWY71jH2MhFC6QKMC8dwsvOjiO0iW7vOpq
DMYZnNPjd0L3r6sP53g3qrzRMCgc/Nnbj/eiGCW9qlpW0wu2TQeSYRRkOQDNGolsutaBu1fq8GbU
OGZSxvSBJnGvGqXkAOBh1xBadoh7Hoz2XBicrBJL+dpKJrsVPALGXJ7eDQahk3+nHhTThi7R0uuQ
McxneUZkDZp6OzEYyJH1an7nDiUT3s0eC++z53FKBEXwIq5yVJ6RhmXu8/mtUVmftX0TeQfbUZFm
1ybTRym10F7VjGCwNmToJ/5fmNMOwbhDNo2JxlD+uCp920biYnAiQ2LTOesbVVzNV1t8v1GD9gS9
29Z4Np1Wa21oCnktMkRUtc/mC1Issqf/OA835ba3BDcQoMfgRhqksbmeB+Nht5eliWgxnoD4ZDfM
paNtc98QVlOcyjwto52EJhvhW3rjJsM7K9nzq8PzA0/We5miCH8QdVb4k62j7NduAkRfFwpNCnUp
2sJL3LHyFQybDBb6SmmQyUcIZn9P7P9U+G6bcWgpLiOWp+W/I59nJpLOAbMVRLzaSD3xEl8um/PO
V8F9H5mAX0CE5EuIGn4XqzsZrZ+zQhPKQZbtvMSN3nuUrxvYdeQg1r0ttOVh6XqlZq0oHZNQH/25
nC5+kOk85bhYLlmoXXmOlEk23WvxzTqPcGLUT1tUXfXpuxltb9C8eTbT+EdO1cKVO4NfKIXRmeTN
ty3Vy0y0wYH9rVO3U2TV36WEgwP4KhwqX7OP4KqEH/G9AQgncSogt+yl7wOvlR2I7iOrkuQBFfSY
kyNb9P/Xj0K1C2tkL+Gvxrao+rLsyMn+iUI3ARgoWlMusje5hurX3AO51XItTDGXVUex8rqSNlMe
V7nZc9JnxUkhCRliIV4B2oyXi9M6OqQcGpyd6cFpY/JsrWz4JPK4oCPTtlk8ZxznT4mt5rWGOlHx
Ve3a2n9bm9+czWH8fPLiHrGyAl3FGjWQHQjj2iuu/FdJisq2ae3j47eJ4RbgsDuz3tmh5qOduCwW
CQd6cl7R7UIZfY3TQWhzp6JlI98eBn936/rH/oNAGeAzn168j9a8INYObadzgad3mfrWZsHkNe+a
1PDltCP2YV0HYs8d6fHobVu63pjMYV3+R9gOKZ9nBRc9xb4Q1a4WeZGcdwlJteHC1WtjlEscCUX3
uoF3obrHi/BvmUVHBg6gZreXTaA9N1py38xywKbr8y9hHCNLSc6ZdgvpiodzfWCB2scOKDOrvVZP
IwQS6M1d2Z88mR17bj3UFgxBLsv5PHy6mNKDw+ZWvD6wCpe7Ia5TsBO8zb531e6LQgGq4CdMwf7X
gpV4bqvKGz1mZ/gKCgiki/xPYVy8VPVwaSKQM2ubzsBMO/Vlczph/gd1OxfwBl1dJ9F+GU12Yyjh
2uGvDs8waVoCkKF7Inwsnyrz7GtdnH1Lou/4Z9HZ9nb5L8ioI3SvyCu/XEy7bkRhUykYzpUusAiR
lxKCDQS/2SmGbc72ndmaemSz5cBHE9xwMGclN0JoJ9aJlyg//FH6E+mZNHUVLreDsjSJvta+CST7
/+82Q7MSdwkuypqGYM3U4cOgm/KfjYSn85FQQEjhq6ghtL4AcU9QB744xx9Qfkd2PZUS8cY3OWVq
WE5rdklHNV+JJFVbGkbxDoIwJRfRza3q49QEhYpJ4BydEdNtbKbq7PRZQn/4pT6O0CEv62wC0n7j
QhCxcrek5QexPb5Fm46PPRjXFhcXLQ9bhJcS4CpaCUT34ykgHfO4RE/tLhCo18+Xh0HJJAP5XYPB
fJnmrp3To4z/ZzaNQArvtXN6NdWfnxtX9S0kPw6+9ubo+wwruDQ5hHYtHR/zTGGnUTxPrApq6tAu
BwlvlZ1PuhsoXo2nA5T7+ILeWJ7YCUI3BiSHtDu5uCwRMPx2hSFyUnAFgNgQqdNvpHAxS9odBrQc
Q63rL8UvxOPMb0wwGG+cxsohPe4rH4aKfCU9tSWiqvsyuUpzT2GuGI3P0+BXVz1kajZy39gmzHFr
Kr76V7yh/yCuOz3bhtM8bKJStMISG0zGLAtuhz2KQ+bcP3X0gpZnm/0AGmr/XFkJSvvh/B4hqz6w
/A03aTqborZ5PsE32v0j1ZcVH3MNpc3+F6fYIHWFUx7Aoq7FjmzwTF/870WXCbf1DccPtH3ZgUt/
7Tq/vKe8ARntRP5mg+eP9qhZ1TzvofVC/4/pZdk2eWxqHm8iopMok15fjuu4vfb8LKqFq3Q/bPQe
tHRyoCoQN+dzjro5jDgqHLeIrmLYMZjGadiSFttegRtqI8MMXevjyzRKmqKd85NBqufrghbvKfXK
cy/BDmjjPCb8yACNilc3xBON9aG8HpezDH6lU1jt19RtbUIgq6FxsHm5u0KrAkUqDAkpoHJs9P5/
3rqQWZ7Q3p8E90fD8inbFiFsYXlityQlcrQ0SQB1KGdTKOE20BGpWmeohmyiRaiy/zERthcSFaeY
41weXoJxYlsR2g0CCetZH5A+jS2ijwIiiGJ8B+JSwShvFR4zu3bSpuhupI7xNahzLIIexAvn21H0
jUK4GGgSbQsxqeAan+gK5D3KyP9C7Ue1dfY+q7vnm8KnHW/3LWsugqsvTWQ4VXNer3qBmQvTSlT4
fmSPYd+C9PS1SHyVvDLaEP7AUktVclhjKL7NE5nZ6gJqHHcmCVAMC81yK3dsG3SxRy66l5M/yGee
ik073h6y7LzMb9qNC/zL661joVbMEgt6CPXHh/QrZ7o2q1v1WaxmTlbqJIpdxVXC8rTko71zG7/u
jRkQCDOvEJTj23kpETiLs8t9dG4ToPkjI5BuhnJzpseR+nPiXuP1SuE7UJ3/+7Ll2pVD2ADQBfRh
HDn5THAv+zv0L6N16a/69ec5w5dPEkr8Z4+8U0VwbbfW/TTOFOzugDQl3xwRujNIDdpPCmPBKa9Z
3EtbXDVHvmlmYAhfvEo9asUfKM2ymKEdx2SOxq12qKmUTUHg74ERAUYNo0O1zlxTjnYKNOGYjpLK
ENe45IA50EcR0wEYlmJxRgZkaKTOnqI9jeO9qYBRvKZFtVS7+NZPXU4tiFxN4GZfhEoFnIOzhuL2
gv+vx11U9FG5DRGYOwpNZyaN82y0n0gDaqyp7P0BHOavj5I58kQa2pkvCtZtxdlgkMiyVDKsf0Sg
4Q7GSPUOllSEFo8paS6+bLKTFjQFegamEMsaparOWRfjd9ERzq+zFwneISPffjTAvC+8hAPg/ftc
2dnrFiaWeVDWvpcTWRLQuYUmA2Cz/7+aLHr6u7pSX75WEvSSpEsF6/v+pOTf15z+GAGLBnrOV7nI
mDm23UzTo3lNW8TVJP/Nwaiv+EteDrHi2NIsh2m2bwfHa3IVkzk8ppaGzQW+geBtRndWGc+XXuTU
YmVw2XiHRUQiA4ktMmTZKDVmxWEn4kSGznRyTXl/zhRAKSdix86lYhCtt/ofD6ZJDMHdZViDwjRz
X4HTHS8LfLx1cdG+y0NhflC4/dIhcmnV+jFAzwDP8D4Zebsz7JQhcQsb19g8dOH4ui18s2qaba01
ID4WKOfotu2XGIyiBWbBFD/KNNfsq3NISbVsonQOy5jQjioKuberegm2DRaPatM5YlZOEFPK/j3R
xfh17FuRKoVarcBdTzRilCBcdjoXI9Ykoi2tcXNPhcTU6xqP/a4gnlcVp72rlTqeDf134BfO0Tz9
locZWnShT7dc1MK4lGWqrEBlMciEwkhaSSx6pwptvjTu1KmxoFQ+rZNrYpE9isQWne37/yFKb5I4
DiX9pF9vAJVkJGT0fh+u31IOSY4iFsc73w9ok9MApez+ErXdwBOwpCp1VptKTEnRchC+J6t6ps8H
Lxy6rY61jxgxhcOpKSJ7hCPd1BrVh0ThRl5ndOYhFDCkCabQQZxznnQRNfZEsx0IT/WejGKsFcIL
OPdrRTbqkY0pMThPoUGJrmmZC3V8uk06hpjbuSqMjFyHOgxDNovtXWiO2NiLzV6LkGAqOJKxMNBb
Gfxtau5iG1FYZF8SJ/sB3da2fDtrX9JBD0yvpIIZ82NHBO3nhUgrz0vjT8UGQIX2DpJR8qian1Cy
ZJiu9sX+2QWgEUc56g4UhKAQ4u0zLIIgc/8ICv9JWX16J6kM/gZhuB4lBAwF0yz+m7dgZ3C7mSRF
z8A3PkR1lvQUIVNrVQJvidjwfm1XLX4xVvdRGGJHHoRN19nUAGP2H/1dndAmxgC8f/0KQJCZ4YGb
5KPuaguBVm9pYxYNaFeJ7IWrKbbBxHZcrR8DwcbLAH1Q/SZmcwL3RT5Mwn90sWHIJPNLqGfdjVAI
M73s0ewJqGOtEmXIKHcylinUWIhHOmtD+FUq7/rYWhlbpno+P1wtI45lnkHGIBsUoD7KllxftnMl
UgKu6lbN6uOQDqEJUcDf7iRJZCUq3/OZ8O5AGfogVvQ0KRLWNjhOBwd1GiFpca5LSBr735w1HznI
BhMjNSUuZoMFqlqVQ+L2vVUnRXcG2PYwsHd4P0bkavsI8ay1Rk0wq0seViX185E39luZENyf0tBY
pAvjGWWzKxGYlZu0d7qSfPKYel5klI/rJm/4SfZuf4GhX3WT32J02Qx5jX8xhXTiW6LRQcCvZjgS
AeT2WQYdL+CreNYm9hIRr5joRX7oLp+Ytjl07KGPr0Q82Ie25M6po5TimBV26YBt/voaQih+LDu2
cDBjC2K3LqEAZvL8yiuDc5z9FHLnJJg/A/jNPBdaqNQrrf8yClEQLzCv0l4eihud+iK3cUdg58bH
2cdtEDg9sh3zT1IbF0p0PxYKglaYC+x+OWph8v986VGWdk8GSytDUYH+W7LQ2X3+LiPjNJyPHKrw
LjcVhgzRCOmmObf186QIBvroOEASpRVZONmXFWDAgJZsrRErxwNgkb08AJeYlkSJCAoNdaecLlX3
CqrZgDeH2H7nFvBKOQkd4djZfI1as/HA9iQOysjR7WJWsQMn9Pg7oRXyR7Z8LR7LjIN/bDKehji6
TSiD/GP1rsLoDWQEFaK3yrwDPm0DHX/Rm8RMlXwKAG8EEFH6Jf/kv5nE/F24pux7bJzHJc3y2i+Q
Vc+QK82u8sdIc9Gkn2OZA7eJaExlgtfb2905XKfqr6MFe0VlIuWIwABNAQ7XDjKv7+1YU0Lb6cpN
VjdbI6Q6HkiFYBtOQo7uXHzpY69dAWty8k6Ar1j43fb0Dxw7CTWe5qXf6nrmIm8dxhFSc4Eut0V6
kaQth7uVPAUeZo/wHnVtTCCuRrzl31sF8TY4PxF86eWLUMpS6N0H2Rtxp71HAzr5ljOMjcR+KvsO
OAAxraD4xY/KviD1WrUC4z7Yb5tB+YXxRauVI+GJM+HEBQ/K/HCg4of9wO1r2LxIh5St8WmeP3On
U9l3uFgeJ3ju5VTSqU4pffaw2Cf+wA2b1hPVOw0BP0BsLKwUucE4269WNfl2kVkAK95aVacsL0cU
x6cXQU+dzgvGXdFv4nlpeLhxq0ZkKyu8W292m6tDe6BT6jG/5yf3OBiWfHY63QNPHjFXhdULnz0O
l/o/Uhe2fYE/SE260rdNqe2FKEI9JzhJnXDriCntARLGg1oLB7sPDz+4vBsjBcGRPGFX3xNhZRKe
RuyEEeFa0rZVYR/NRFsCvbGObYx00Hoi4yn2Shv4oIPbWHDBxh5Qa+B8IgJ9j+sGkmRHZMExlnQ+
kd5WatS/AUXgpfeecZz2zziTtZ/H7QajXCAqMgWfxPTRAh5y3i0r/4rxp25qjKzUZF6JCFQ3PhQz
Pow1OfLKL/iqD+BAl2kthMOYZCGZSrDnu1BXMD3qzfeiMNuVg8xOw39LfXCufT3VBnyUU/z+Vk5b
8JstAIVu3vp5TfTiPhe2ZzADD2/Z2mTsx8e5Xd/37uUS51b+KGb63tynlmlSON7kAjR0PmxpJeUL
+eDw3YEaj39fpsBX/YTv33XE+L+W7a/xto2+eER9mfI13lw/ZqCi6uX3/2+h+Hz9lFyKqHFbVK81
KPMAIVQ3gNyy0nu9mACTr6rHC8sQ+rKUZv8RGaHzGF67K6SAhsVCWzLqiNQvpisAgQZYCdOaeohK
EP/dAx0kHm0jdpag3x6LbxE42hbcBAKXGy6VYyYaMxICYnaQAzZ6bfQrg6fSwK0KsGnZa7rl/VPU
Txk5upfMZtrom3NA/GKoNpB5gt5bpb9sc5wpeTBzPn6FY7eHauU6DOCS0mS5VhohSvDXp6FI7H2q
rGkkWpz1IEOPv4xJs7+yHwyg1d5iHTczbWmPPkuEdV/TDpbfS3W0vcEdd5pRADlY3le6HHSl9622
3IHmu6nTuQSFIuLBWL0nDRnToyATARzU+jppZNQwLpI6VoH9AFtuqToCPBogZRC+z3hVqvP/EUuH
tqLO0BIk0b5DB1t2hgyTmprqbl2d9KjmYEUA+Hqmjd6KbPqDyrC7kuHna0VRSB+cbpRM2Dzmeq5B
qTDhAroJNaG0GAxLFwELxxUmdZFYVtkyY90brRBxZqd1PHSxOHu8+yX9phk+r7Fg7B3L25PAEc68
yrqQI+kGAUuJWRxm0BmHnIPjPQVoitiUt1jsUr9GU3pCXXWSu7wOQ4nb57+3IvRFNFnaR4S8+mrD
Sdcu4tUoWLYgJfN+DAlf7StCMHHk40iFLs9rPQ99SzE+LjyJZpDRG8HBjhxBm/29aXsr2udCmepe
z2mjsH1OYo3x8+/M0EMwLNr7XttXDErEsLBIHqdo64L/1wLhVvxGzVwet3M1rclfTYaDJthXXuJG
O4L82QrQ4v77Y1+cxYYGpzra0mYlWzGheaWUhFqcPD2uMsBA1mKXs74FCL+f4b/vOODjJ6u6YdYE
h1u0NxI3iBlYkm4dg/Ad5XokK064BCD94r7ek/Gy8arnGiDBNHpXn/K80qKSIobXSlsuLTnXJeDy
kKJnwSEENfAW1CG5Wm/W9jgRgFwzscn0f37Z1CPTk0RxveSQiO5NCaoxs1Y0mmLD7JVFvKwSsDPP
wmDdJk4oQtYfTtubAc6sZgaVey1XT9jb/taOE4jUSqcarEiPj+Xu+Fhh40HKGE9gJltAVZZEhSdX
5XS3eejSvOOzvPrtRfT/qQKm+aRybSswoLn6UDAnAjIPEv9CdnWjXvh16fqt3sFYz3d+BkepcB1o
DC+CoPl3bce9pmwnjGpsp0l3dlX770Uz15wm01JXaf8ELbTWKjEGdmUXZ1a6Iaz5seWgipMOeQSd
Gq1oWlG8VfIdl+msVCIIxAi36zkSd3S9mBhtjflHstyvoakqTX+j2X1ZW9BmN6Spsv6xkrxzk6r8
bSyoYA5GSRS/Yi9ue5Y1wP2J8YHcLyH/h2Xxl+x+IkTrB+qElk7fQGACtO1H6tB7yw2TUrMUYdPl
z+0P3hFPSO6Tp0ofl1zd/+SVzW7uyoDBZv9CsdC+dbuWmlGEqQnfbiuJ3S5ACIAX2AMjGSH4EZMS
6tcq+b0vItKZFZR/LqBqQEEYovDAfgiDGl69k6p6F/USvLSLesNfbUNvhtY5WhFHgdUmlxo1i/82
fVvCq0pXhkNv/HSzsZop0wejYHDxnDMxbLH5a49JzAhk8JJqCfvhGiLwoHc+GUyTVYiCYVbdV/SW
sLZ4jKirNtMIl+T0ka9fDNk36zWYxTN5ggUr1SLnID54YXejN/8C8SX9r6i+oKhVI8XIa9y65ZT0
gh2/iWDKqjoKHecwFq9JEgitg3HMKGzBXrFiUzGF7olrl5+mcZJqBho4OXJzZG7/ot+bSxB+eX67
i3mVtn4CsACKZ/biIB9sCUgWTjqfucjPLvXx9wHCuu5axou/imkSjIMQW8duCe+2gLoNLqflkuCy
TzaoaRtDrQwbhf2Rlxxnx08shWeH0R925cYNS4v9YxX8Q/k+AJLm3fdJp+4WL2CS0pIdhX5mfwbC
ooXaO+H77NHVr7NZPAmL1d4+1NlEheY3PDsc+672OsYim82/Y6D084cHpTH4+PF4hNjYhC18YUNj
vOELJY9LRnDhVMXw8AXQCW/TFEXUiLe1HzadpNBRlw7UdO90W1zI5/kB5T8BtebQOaVgLKUBsCEE
H/HdtCggl+p4eVYi91BCTX+vBvstLDyuJmyt4DqqU4RVD/zRA5CFIy3nblSecwsbpvTvFDGFpLS4
aX+PyGSZ9JRenaMdGOs7dOrWxORooMgpRXHV+yJw14swbTORqIRjKa4gnc3mm3SKAo7Ee6whb38i
XZVYG2xyiaH/eT8KY0ONEd5CrHhFnzKy1DvBekOrUiVzXpFsCsWz2sTV3xdrvjWMjuWCZYO7TDBW
fW5ZXBCy5gcvgAwtHvlKDknA3rnbH6SiTSO96EYGD7cqUd7s9XHXA1BVwz3yweAZaSyJB7Bby/Ff
6Bdc+IVHVym0KB0Obj7d06N6UndFCDRydp5RSFI/JmzN+vYiG497rch+wxjoeExkxuPn7MDxZKMJ
NWuE9NKZniWJWzLIcVkWMqMsL5KbUrgi6J5hjwYZsMdPB9fkYfmXFrFHrzREXhau3stLY6KiFu+V
HX4gpsUh7dIXsg7y7ed+e8zJVMS21mskgoBrBnHRAPh7bPdlMxImkXRM76+BtZTQAMljVq9MZMdK
6mrynC3jz15oIoi4vU+o1SFePBlxQnTdDlJz8QFLoYL+zztBtOnGHWXwriVL1YyxfVNjUKZja9+G
XpVGmZPmme4A54X+9nQuqCHa0IBMKAHh29v0CezBXkkJh4ra30Rg/upjmHQfjdT6YRy7q1p6lAdD
NZqRk8vLSX5NHNiFAUxa7dVeVBhe9qawYP4btHVRf469kmNNpbrjPxnJhgJT1488+5c2uOwdS3wQ
hpF/wpl4FUWkWskIoYlca3Kyo37b65Y+G4ovHqZE6y9kykKoMew+5JBCyNScQ2o7lFM2UZ9qCW4X
v+mpqcdGmCm5q5IRWKuxeoyYWozNhvYZiiHe7la1SXoVQAYNVCazZzFQweCZZbfHuxN4tWp/ICgh
SRSZX/107IX3ADSnqfI7KdDCZnu/2Hrd5Lvn8evaP4bcyUagwpC60hcdDBLgBS6RJQvrz2N13j29
saXkYqVECba71lypuMQnpo+GLjb2BcEHGCUv3HJF10Zuk5Yo2YaokkCLXHyiksl/iXDYM4omj6kP
BMAPeJxBhbSgcniL8+bcno5jLtgp/VuOhmF+vor5KTY3yX3RKQDNpaJBAxaL3X8szyOdFXhGvaWI
f8G2fd/+ZUX+1aXV1jYKNeBBcdXQjDNJxWtlEvjIUt0PCHpxVrvbZg0je+T0XdoAbixTQvtYBoQe
zXq01QjfXbTbjt9QdqAB2EYfOuVWNOM2oawkVM54l4DqrKEqgJGUMOCU5WxX/g8s3PiDzIJJQJT8
F4Ly0lvMxOHuDlzNoW0C3voLPpKQHZN426Jg0r15wn8coIE39k/VUf8d/ZPTQBchUPJdeqQj84qQ
/pf04fnFqyLBzyKefPxZFHxqbjscANsdCoRJoaZatcGVhmfviG/tOCbO5VwmlG8F7P7OSaYTCwGl
ZBZER76uU7ankkOXxOegww3j/YhSwRsJox5P+iJbk4EAjoIUbgvZcA8eREtUI3wmCB0+24Vp4oEw
8gMp2OUulvYbQgeP0hHDEuhCmfi1N9M6FQ8tq6urnBtY4yPIz7zcn01Fp+I6g9Cp3KR29SEP6tbu
CKJ5tJLw4tv66CRHAt/UPE+rpJuegxaBwBWMnNCvJsDje2SKKZJR5pbGhBqARbNWrTx5/ey03FBl
kLQUNrpc90IBtJN7bSlB6/CV/wquyxM4i9APysLmBxGQ9yF3Yrq8TW+qiqNlkMvMPzf+JMoxPTq3
zCgi60lHORKXSrrJw0ZLXrVvbPrJhKJ/ysJsWBlgiCYcw/RHxCu+jPPdFdtRinVcGRgKqbf+ujmy
0kcfxwkQDIIywrlrwZ/h6c20QcN/uRX/km6D+uRe0qe+zPup0pyCpBo+MQPTl6FthBEV/8H9HAVL
4eg9Um7KOC0zS2Kx0pVuSXKqm6JoOTPlY08pN2VqfwrVgwt7r8FwiIqRbpxM983WrMiqmu8n6u+C
qH2GqzdqNEPZdY1q/jla2PakbOO5FQJ9pwEvIJiUiJcePUaEUriV0tXkGUR8HNtZoWwsNCR6WK43
mVUnr0WtZa1jgGc8ngOCWyrzxzNfYDiQ3/3EATfvuBiqpp2C4b4BeLvC8/MYOpsMT8vk/2ZF8P7F
wHazmOSL3cZ/AbWdPIribnm1VAfbnYlDMJB0c3b0hmiqkkuIlTet+gZFKJoh5TAndzYP5VCy64SH
dmfp8GZ0Bdd+R9CaTpdl/dbdJ8WQ+bzEQDgaCQI+xDTqzPKFPtlY0CD/IPyj4sPxkDKxJmbRciC4
974zcpsXCPrgbGSLRTPz4grzgEsR79+QgL8p3gnM0NC4weZcMrB9PM9bUVcr3kNeOFiJwOBBkArh
DbU4WDi/9hz5XVdJrxcISojxMcSLSxCc4L1EXZdyL6DWDaL1bCcEsFrEP1lGCyyFEn2bm8ku9jhc
t+Ji7BEtO4NTWJKEYol8tOhsW0Vzhdo/gJCHao6XBLXjwTgjy1OYZIQo1Lu2wvfnQghcBJCpm7Sa
bDxM2Ftb5sMIA1ro9GQ0dXr9XBOr2FZretXVWtc7vsvqinJtrehm1QiKCzv8o7KmWIr2Q2XiUGKT
Ssxw9/Fg4dnvEiYo6DDiJ7+A63/7R9a18kUsO4KP/NCKQTYAAGprivJFWvySKkYvOy/coZVSFwXR
70rX8lmWVBklWYWHswj0JUIgNvfhNDCVbpz2wa/6mlKIu2sysmv8Q16Y+vdOAs9bqDU4Pypte5SH
n/Mr+ZuSl5Nsi92NA5iSeQ2R/9DC48k4x2T+5iKGIOW8dEFmUFZjF7SbGBLvALUQkInuhrlAa372
jKEiGkxtQF+ERyL1Ro8u0NWd2PvFBm1HUZhTLyhiMVIovXdxtCxah2alN8XJ/ZM5IdbHlWrb9hxY
v1xk1EyHhiQxj1nB4+qWPJjwtBsBF1dwibxLg34BP5SDCMZQKWDhwKxK00pFEgWpPivSeH5CXI4L
0s7mGwmh4B13cS2U4aKdkXaaYdZx6ShERKX8md2CqN0LRDGliXQQhq/biiJGY/YpTsFoCu4YT4NP
Uw0hBRGcfYjJJyDokc+NKSGPMg6Z+Xcqz/EEXO9LswKJANG4h6NJo7sU7fdqpyRtNKZtb0e3Oyvt
63Z0/2vVhSXBUNuhvt0QVHVpqP3VyzLV0kSG0lpn6j7QaN16aIPd9f2Iqtdye8s0oYdYPPA15Kq6
e0auLM65m6Ol8zuYf+ZylPvagSyCy8snz8L+hFyAhiqTdt68GfxeM+F6JuSzbXYsDFz0rZzgE9aS
/pllfR4jBFKftbEnMHqBIFQvJzZjSNBYoeF9hJvufgnjrVh20/hT/ehutTniBgGLaQFgju+XqFc4
rc8zIL1BM6l3WSpqqtkIiaSXPU23NFiv0DLqFGhYQK/P2qn3QY9tQSZlxHgSz0FWDSJtca0LJd1+
37AHpoedTtcgVMJlt83zncTi8aydfKui/1fgwBMhrIb+ygnK55G0Pv5nM7cGI4/AVA7uJF1NF4jR
RPwgtE+wAyp1KzqdIY7aIJKgYXlEiRA3OreY+9FIaUW3w2VRVmuy5cpnIaQXCmmAwkLKlB2kY1/z
/I4eL3DNLnL9wdkbEhtSQnZFIBuayKYn6T0eI6Dt6i3R+lamm+ANYghKODzb3rRRCYGJdkWmvUxi
sB/6h9nJARYzwgsZAX1fVrC4AsO+uDGJk0tOCIqpvy916DHJnVcHKZ1ie2DftHDIDVdNJju6eqhY
B2UjIn+YeyLwV4rsX4xFHSuBctachG5fcUGpg+60m55LKYDvjSVpLRcjpre8sgaVxxXOYI3/ROgR
lnSjx8JTeCQuaiVrEVCKwXWJPK831ep198Bj767rmFgZ6nUwTWWgEOYW2FzEFJpmb0rXvyMm9FU9
ZRWRuPOIlheafKarsZ+/A6HifVSkkOsIMQTqcQrjETSVoYyZtGuWyix0+fjm3BbgjewfuX2rhfDC
WVwhbF53kbDRz2Ayc3X65l0jr2yyNSWef3v0frdWcH/3UK4bfbG1KniJ7mVNsLmHS4h0RQvjPJc5
kNem2KRbKM9gpcMsYN6iWa4YB4+W9yCTS0DdChwSRo8oKlrJXoDUYc4JnxmeqD2Xz93ZeC2K0k1n
61udfT48cI8GSrppugafh0Ioeq5j6kVqu41h7P+dQHGoyIyPfUu3spuVpQ6FGlC5iI4m2IjKruYJ
XDrhZxnfqnUS74Blfdy9hdbpr2P7zs4lcCDOz+CBon4ccMVnw6MEPPc1IF0rzyK7aZMp1DfQyFXO
cryh8pAFWkMS0jFziqEdW/qtQpPai7KcpmeGHkQNwzZYBruP6UDj52VUV5nudkziAH4S8yHNPj+Q
t3kvAlWpAng/8l4uVEvNefIVv3YYgu/eMAbkycrh1Iv8fqXYKAiz+MVjka1lNUR2PSFo39kp0sPW
ZzuwJkoIyyLOYyorZisKvP7Wws40QiKd2h4v6leBEvBtT1sNQz8p0IvXZ/wRuPFNZany4qSWwyxA
990Z++bODxYin5trdfHWaxFptpjz4cdsJ/wyQh1yHG08l2LJhylpM9dl3ITXVVGaCiMTgRl7e+Sz
UmXtpmhv4DJaQGcNAThGXlxWDHxgqQs826fiTMmyv7EbKFtcMvDxtlUcvpdrsun6hpwUuxEFLgDS
tOMIs2p4/x1XSE3rZE8iw9ps4hAMeXkyJl044+L/OMwumnkf0TmpGOazku26i+ub9mzIwnPjC4p5
UyU5qp1QbEJxvwyQtU3/wf6yp8tZ5qf5vPrXgXw+uxf3QGP5yvuKZjxVD1GN6aZj49NlA/EIMJTr
9QFlZIB83kSlEjg/xY4RGuBrpBX1TZ/MiG3qolxn4JGc6h6ISnWWZqq/HgWeMoq/MVkC93zmXxVI
AM0pzfP14K85RoukBY4ikJH6NCDeIVnv3N2eab2i2Bsor+sA02lhBYrIzXV0YBhynvpR3EPrS3VT
qUWJsscRSiK4XXeQpEuwvJtFPE820rFQwq2TokK1eUX7kytMNN8YPCr4IZGgbuzsiXyNcsqkrkFx
Pi4nZbtd406h/8LfjMZG8fGzjNy02MoWnSyrH1x7fSnu1Ku7t8VZdFl7MTYYtRIyQG592Ck5MNdF
x66Oc2hsp0haOt0cvLWEQ8Kry96TGCZsCtxmRWmqwtRdbEsguPX9bBmhgM54Pn4TppajQvJeZYkx
Iiia+OnVYPyI62QX4hYdYVoSKhrIvU7DP3p7eVQMdw05CUsripuLtiBKTjKBwEgVI12NLilCZSVs
98l0jBFghFkXzdzzWys7uT2fQhC0sRo5q9PEm7yDjnCaLCTg/3y/SpiG/tN2dCCG5MHRobQ7VD7p
SS/1IfHLsxJzGjEDW+lwsJcjIqDoKjGWmiYDe9HB2yRo3N3x8Gmrl8WPDMh+w4sjY5T5j6++DI2b
vJXejEMmoAxUHv0JLh0DN4CHF9N5xsshMG/VZK8dUPJoqq6xqlhmDkHoHHyrJcqvZJkKLIqsQuWi
VBzeAw5tqxL2yD+7CCfhOSwJTLIsWlk9z3A4SmdvDHYaPi8nAAqim/MD14uy/QphXP0tRg7UYWFU
sIo0349b/FGt3tZgMw7GZh0gDJtljuTUyM7kfYg0a6jSXujNKde6D16FIvaAmhAhkoIdkPD/afek
h4638auzVoe1wOpVQIXd25eUWAW59BLcmOaR4z1uMo76JF45DcUnyektvfwmxTQYWymr/GaKkHLn
b3+ATp+hKkXzM1huaeQJpsPPcS69luOjS4LgW3iIZ82ZrzF8PcwTJEndoOYbEcu2gZL0h3/+brLZ
9fXy9s/8hHPKJGChrnBEyLT8UtzNQ3eodsLwBnlkeJKOe4gnnuvZ9VpLqEHLxs/+SDSxjvgNtete
EA0Ibqq5TWEk3x12HBT3Z16fiXKPzP6guyPqH481YtVkF22NyJdaKF9IswITK9I462pk97i4GLen
fJu3+MuBpU4Cc7EBbtpnSM3QTtfxrb6niGu2gEAJ2vge2MqUf4TJvAhREEcxGb3EoK7ZlI4sliQP
vZFP1c9N50sKlaVOSdrb0fr/AXDjY0uTbKQOfXdraOC7KV+ApMzbseELRWtRRHWsmcpGwm00o1db
A6vVCPgtoLVJxo2/gWAewmlERB6amjMEM7YKEaYgAt7PmjzOwOO5DXnqd6Qn5CXby/26rMeeyXfE
GyDR9dTpAzdiVO3YpV1CDiBLkMNYR3cpUNV/9qYnFT9bbsBtkLRd20xsgBrWhgnfHT/Tbw77RUfh
bgQalScArFyF6rCtYT5N1VR7btEz4vwpOwYdpenFtK84rTV6cfND2C5IBxan5bAKSxv8ipcu88DF
u2wa9njrPNtKruvL4cfLNEZwWCevZ7Dks79GQNtjkpf/1TPZmhGzuU6CH4JWgUXGsGyGcEKAIi9k
o1Q3xti81pGjyQlm50IQm7VcEPZxkm+WQxiFJG25pVS79lQj8LC4D8mhXH7rOSregu2AHIrLDtpl
aiBAKPZhszsPYyoWe86R+vt5i3u3XNUBZz2OlxguRGuztAr6D7MmxUvwf4c69lyE/41ihDENabtZ
PU1SCJmY7QIsMCsQRHOJy7nXaiiESpZi+xA2Qwo3wt/NML4uRC1qhu+L0ZsDlWWsQabotZpC8Ngy
W+hCIUzRKtRqYjLgYVVe80aWteiwtds5usRXC6rZnAp4hdi20P7x6hobYuvwTq8cNyuBJ1ivnvae
yQT0owRU/qDB0P3GrJMh2UsrWF2uDYZzfID9j6S8AXnmPUDxzfR3ZvKpk6JpiPO1ZfHHIdVOUUol
E0Ow5h3vgfWRw9sxlKYhbXgcRFA2duaSeNJ2QtNolUiA3uWpnSiki98zeWbTeYC4xsKQ0xC/XyuJ
+n1YWAUOAZ6Q+YWxa6yU0Ggu8eORmLs2aS6zR2c0yWVOCe2b1EHPMyixUcVzfeAE4TPoBJzWSD7r
Oy6i9qDOueT56NAHKPTvj0aI1K5mZqhsqCPWP9aO8xN2ByymFLshL0otHdgP4Nx5DxZS+ffgRiJP
4f8R6KoiJlXiHTBSJkMBHEY+IUjhnCK+MRpC2LFZqGyCgoIPZEJ1Ow7I35CUlv2TM95GphXeinxt
bA1D4T7lisltbaPgHXJrgdAPayzr0xloaHUECdc57JJpG7AfGgYKQjTmcOTT6qannZFBJX0/XiRd
emIhywr7KHRVmiCizM3FRF0r8ErXPV74dNKXIUEZtuoMj3PyVdobyD4AKDx9hj9UAdGXZf0MkVVk
9ZddrYGOYUUY6pUOPAFW9pXbi9f5YQlbtinWgW3yQWCDnA6q5eufiZ406Hd5LWhSixAQmzwM+cWT
6pCapQSfUTKJev0odhW6H/XWkskilFWZHKxx8ELT0lYjJSplAwgzbO+EZ5rq+IVbUpBaQfu7OPzE
cIg/Of454UXedS95G28JU5QgT5BQbEcM3UcqLr/WyRJaTbElXjwOJV8/F9K2RR60gS7Glp1qhEK1
jzJSZQSBw55FfEge22SrhYCr1+aVUrMZjN2hseIy6cNPQDdT9Yz/zYHplYfNg9IkB9GLr4Yz9LTe
zqS1holF7lnUJrBpng6mkasbZmxTGRvoTI8oovk29SeQjBpQYNC+rwE/WkCSbOtoqiF3SuD920Ep
mZAMdnrb5RuLy8wZQZey5Ws0VUptEEdcRQsvHkC4YEVOIjpY9IfIxZjwataVwgaG4DWp3+8uhPrr
H3/Pth+rU2BUuB1wlXhj7b/Rk+EpAJp20B9U8U2j+PMUM1NqWuCAw7SpXoKFg9cLfmanMwo0BHPA
yqZr8tylm5Ui91petaYq9l2pj26QP9Z7Nr5CG/n/YHQMa8lkV/rt5IKq2lnyq/JsKRHLsNkeuJYr
CoAy4Pj79ve716RmFRgy1qvVFjPKxwM9cUjlv/Vt4cQ3dbgu2XP+p7qwFdF54zQe6yePC/cxzBhw
YUqlncH5orhU+T9LbIfsNpDqhtNtH3K3y5Aa0KS/QjcP8ays3R2Knx45Ygsd+px1hIvRvwULiCC8
OWRxUSsrLZ3aJg4DpfzPfej5uN3lxUVBiXQ0lajcI74SfQGFzvZlsHXfwilur+dy0hEy4QxAEHU6
DTDyuQlIhrrugTyo4mZ2Svdh4HorDprUU1rVgAvnuZpi7IGMb9m/8oQH7C+jSG++bIyJAsZYm6KS
37aiT8IFDrkzcEpJ/aLFplu1VDDXA3cWrNjbhTkQcwh57bm216+8Oi/7QSuPfYpdiCod3UuJ3ykQ
aYFkA267FKZdM/UDTbGoosaMvfsvGSV/dJ+TZmKl4RtHT7/Mp0cXKjZFH3Os4o1O5zor0QTGe/dN
UmiTXW0FsYvG6UhbBrTmnkBbu9gpBi8CgrKz6hZO2DywfhVTwdzN8es7wA5IcPYQ01o9x0xe++Es
Y0PVtfhV3YdZvravDAGplshJrXNCvYjieU8zckldqRVi+3of1SXhX7N88uWSPo1OnIvEDU7JfZbS
PzD2kRZy7eP/uorIbaWktCDxQE3b9Qxc5AyqprkqY/IKL/5ZV7i+p6sS9Xg4SivJS4en5xIgsW7P
2T8cfqepAAKGj58bM4bIUGzA3JrAdquvJcOBV+WeHFiu0Q1G1q2M9KgyXs7kkhxrjSxJ50XRKjfC
00rPLv3fd0D9tcUf/EBpQBem+II8mPTMY6dBClZmkOHlVyygwRzEb04AX5oYWF80cCfx6RAFaPqh
wCPqX19b5W+fJdPSzqhJ8+MKLZlwvciCGxKUTcmuhNmHDjwjEcf1ntg5hBnlLAvSuF+kw8kF4cYa
kivyz2pj7zOtMfZv0VCf/i4mdbOtolC2uTST/3hqbz3bHvMMeDSOLa40lwIwgovuEvssYmSXqBgW
IfzvGM8HCRPv9c8iGnynlA8IJc2LlAZn+yX5aK03VlGpUdbWhIEH7A4NQfGrXjNWktLoCL/lod3G
7GduGXpLYAVBEw54eLqQgFlNqxtNxbhvu7Sj5w9zOVYVQsZWWKPv8M5EZmO/ecODHreNET2lpwso
Opr6j4AGiJbrHqg7Oz2qUHwn54ix1F2feajFu1CQBQ5huv8Tf3Lc/HT6xjTMxD95asFZ0/zK9YGk
7IFWj1ivO6eI11fKB/IXlQPSUGTxnt9hb8mRPV2u206sp9qzm497mp9Yov39+8axI65S+CCeNE1D
Y9p1rxCnLIH1aeUAhgXw4fOX/97w3EgA6tH8zDnZ/7UgtLLGc2WBvL/wLsEITy61CGRWD/CXos2r
HNPtWGPmnZMh9wljKYBwi81rS14KJNrG8ZqDd0BmgzaM9ukxLQxPy0vpWd4JC50cWNGQ0Gc4KuAP
yPGKZPc8COY4lO4yw6ewBGPVkFFznzfr1404uu2CpQPI7i1qLJNmyAawcRGnWohI2C0q6TjO88jM
mUlkSYTv21kCvYGKLVF7VQ06PqpfXN5ZEgGYDt9MXj6COQ6+bjzXh6rmdj4qlZwfWmyw7Ur12ELX
bM2DMFxNm8Q1a03b1O5IUOg6dQ8PUTGIg7pnVvDSMIBiNQeUIPA/nBqKswVL+OSrY5axMpEZq4ec
TZewdCUGF1YTnx8cKhy9yyW1yqMM7D/f41OfzuPVmEVqV+JbgwFZID83ykTBGM7jSB/VtGd+2DZE
Vv0pGWefFfU3p/IwVOXeow2hN/x83yPm96G+Ai3PoXRUZn+wE4MET3+LNjISy0UHrKT+jU8ptZmw
RE5qxetoteixsik3W2CisrZEiAT0dPfPFCUcyJpAuZ0l+PO9jAHz4ZRQGqLqRRqWkYoAxEsprnGq
1P2oF+nwSMmSTuNK6dVs42mcu36YvCQAxexaWH6fdvXKp9t88adCUmN+7F/QCA92HrF4lpB4cZZ2
PFx8flt94cpX+A1pl3EmDvT7PriCgkiL7W0o+Mv/GaBE8MQbGBSuFKj33Z1D0mhy6L9jRjJaWFw4
kjcqxL4fxgJ2LBeHGyysLlBUdi0JaXep1yT7k3kaflBQHFMrCKAqp+wwzcsimRo95opN8Xs27+3Q
05R0rR56ygapM4bGPp+x/s6Ve79xFFBvuHYoYuzqr7NL8yMeoSjxUz463rJZtsGyLY+RoJ9YHWeG
1ONARCgn9oa7N/CaxaVSQiaqjCElJayh+U6M+7VQFg4+dC52iVZF/xnvXVlXY1ldkzd+05uX073u
YV8kVddVPhRNlfb0/GDGDIfSyE6fQenJcFvlritog8c+Xl12V/kDmSq2gN6yYd9oaxBm7LTpacK1
h5lCxaqWNgPAblAAOcTFeFsy4MSaqiM+xN9mjxZza6uFEvIuFdhC6GxJJIawYtnQCQkliDHSSQJH
niT5kJHNCfNbz+MiGKWcqzn5wizs+WqMCAbDpihLptJ9ADL48QfUL23CzxEFFbTrh/0C8OreITrk
CNrKdVtmY+HjUtyxTFraO2WGiveHGZl+HAFgGwItg9HAduTBf07VdMR3jZQhWmHOvBFBX85iOEyO
0zHh5YCyiCO58jL0Pt1tmkrKA3zUfFasgct8E72n8D0fiR3yGBcwj98UYUnPCekISI6HDB5u9iTV
7zBkdazKJwoRub37QbYCSu13Jj7L9vJqnH4oygvwxmd1lGVO9q6r62BVgUucaKCMDL7AFo36SxfH
QNiMpWjfgs3gG+lXDUogSpsFkk3W1MgyVl6cvYZMoBlfqR+v5U4iqqQBiIo4whgwiH925Sp9TcEm
OZeYhGPWc1nut7pY+FKx2vlABep1usFEH8fvsHtft+qaEOhLV5BeOWbi/fiKcKtu6g0KCjZbOrVE
YuBpMztKA5zbzsMXqRsVj0KSqVZAS+zLrXdmaTR32M1Vq7tZWCFJAHjdJ50Lcr+8wqtIZ2cGpBaZ
CwG/HcRRRCtU231dfMW7kjQDhHubZ5Ueq5/Nhgt4Mn5piyu2iVsYfc0feGvei1lSHam9V43rVgEr
67sDZjEtwCDL5YhXDJqgmZfHJhu+Np+r1ceB1At/VgpIfz6ntkXda5RT3EjatoFkdtD1HV2C9IHV
ts8lAKokvl7K0GSj9YH8MJaiHuGjCcr4zTOQ3Cz9fijDCHKt4eKSj/3LAYs7HtKSwpUfNnVzsgOI
hVtkwUKYJF2sSehipWlkm4+epPaDFAd+qX+S2IL16MSSPIehPi/LRwfdtB2CDXXbYuyQJbe1p+/S
5PVggnuvAzpKzNNOviiN1fBKo6LQDxbUr7GTJcQUsOVkZtCxK4Y0bQU86WuzyTqE/gr8mYgbziLd
4cD+1XsJgXU2/WjRFeqehGrsAYiolAhhkxDsx7gdg5heXDV99DdrWhZEgrHOzxiCv+5H2imBhBwi
vqucYXgLpKcLXhhExBeAA+ValVyaLGBeaw8YEmq7V54oG3a+Y3I/qibJgf+Ba4gefT5mRbT/7bZK
Qe6d4ZPiFVinz/b0OfS9FBQ7p9zx55rTIl+PQkgs/vug8yFPG2NEWJlZOL5w7d3X5XmSoI0gBcui
bEtDF0t2PiEu5TBrhwITSy9qvg9fUQZCmECwvFSm7iEELV3G2if2YOicI18ibF0tM/xFLi463Des
DvVUv45LmC3edNGpwEcKKbPUPcpT7fDPReWluYIAd3cIFb/qneDa8CfVzl+MNCQ/hncaguwSWsdE
cdX7TqXEHZmeXOPOdfhozK8yP5tyhTFje6SIXFEqygM8PRDkwggJCtTNxE3shuvt+LgcE87jQnNw
EtUAfxi3uHim+6/HCwmaQD982NPjLpZdazXMBMmp02Ybg2CHcoP0XpQ5jz++9uJlDU1uy9D7fnvt
bbjfpx018FCloPeGVHldyo2apBs5o81AlV65X2qxora+y5BFHayiMZnq6Q8pPZYDaKpq9mnGL0fk
lTe7h0trZCAKQ1/idJdrqpTvA30x2uK60sqHTUylY/LXx8x/BD8bJ+P5LHUKGm8aTQ9/eXbnR0mf
Tt+IeoTJgnEBourP8LZeXzaRF2LYiaK7p0A0YYpuYaIxDFCznmxPNpvb19tthODKfxOREQ+gu4hN
lHoVG/AjjvoQ1wTaw5y8hlfE3Uy3Sx1h29WtH9Gq5Xt9T3VnI4i39ZoLcEcX9cP6L5N0kyNKrWB+
jg+vbOK620eTZHeoi00Ztazo7nyToDTlMkifhrVMuLRhrLgToi0OIzL/wvAD0sogQD/vFdBr6VGs
He7a5sbFYRHZOzm6+qaPkBbn+WW8T5EbTKsc0jyD/lERL+00EkTI3uJKZ5w9bWkZXfurK0TNhPhp
7+6ybzxf6LHs8vv2+eyDPu6TmFdU5I4uXglIYpdw5g5FLxiJsFy57m3utq6xMjExwDb692UvOcUe
t2d7+3YaE5kwhywQGJEtS7XkNtp83n7/a0ijDYGgO+Zps/yJ67eeEbbIGO8TccpnqNVz3T1k+zbJ
MypDLYLcVlO0CPCsyJus5qEXS7fDnMitEKnS7dDtN9cwNVx+DqJB50lM1HVK2g31T/t7GW3/j0hN
bTAWNrRn8KrM37+nbYEEmayi0iiaxJX03AQrNmYTR9n9igjpmVvmhPBzFobWL5I68jMAYIOZhQIo
WMrXQmsWKcg9n2FJXRzX+xP/6CU7uvz6sadWqlYRAi9avPl163HSPFfvXLOUSSphaBORVySCWedg
Qap+Z88x9oKxI4QAqVYmEMS6YEmvctaTcMEG8q2+yevyhdV7OgnqRmHpx1fVbtMul33i2028uduq
UzXvcpDufwk43RPmA1YT7MoFs+MDQ3BbH0rxKmWOk/h9RTXbSLNZcL0Q4y7K+MOS4npuNSBOHVFC
GYZLoowWivjNbNnj7z+0kqDgOSK4xTKbhpKYckLfirxznT5GCyMZ5pkDrYrOlPL1bdt+5Lwzk6op
KT211JPlTwVvfjNZo2w5Vl171A4s4OQMzb7WL7tGWWF6LDTT7GuJ8/MttvxHrAv194md1cBO70f5
lJW6ArSn6MCZl3CB2RBAPN7yROuVjNr21NonFaloA3RjB4h03bOO4+LPGVe3cnPM/6KHitfVXJBS
xqhW/Pb/5MgSnvHAYdLzXMLLGPP/V18PdGJ2952DYO6/Poc6D8nsgL4GKZzHsRiJc52ikdmp8Oie
v99x4RuvLfhSOALAXvoG+5+YQxubNkwE+EhyK8amWriANZz0zqKziFTUSXKBMpHJ8NTTWDoKyyZy
8crp4UWtnjk2EJCTHgOL9UfsVuXawqvSvEmH3ePLjZ4Ec7NanMjyal/nRJu/11Zb/0Mc/ap5KryY
4/JhW8PWsaoFEHi006hp+wKkmjkYoBtovZEXZLysRSKES5n4kGSEwWyUfmbR3TrrLz+RFZtvaAX2
W8RFsyIPRCZNemAvANBCFL2w6vbwBG4dG5gAVeJcyJRUWN4H7l6kb+n1QsMlT3u7ThyczTMcmiJs
u4htx8E4LAdudwkrOr5ZjP4MRdDg4IeWG25CWwd4abQGzZI//0puqHj54GuI7+NSpjjZsOl0AMdK
or6/Mj9JmMkKSK4p3YpZSc5t4MHd3WiX4nEixd/8CNE0owG5SB9N6SFI+7yEtmIfRS0BqTR6AnZm
2HSP1laICB0fLnaA3qeU9kY/bnjTl0OSafJqZaN4uLZRuf/p1/3mP6GoAz14qsJKfWD8vYtvRXWR
CGQ2V1JfgOWmmsFva4hoYV7cFqd3BakQ+oX4InR+5Ox4BlwbJj1zCOPVeY/owoONym6O4VENkxQ3
eFpiaX8LhTtuoIx0zk2WD3gRpYaeo+NHph7ZFN+k9Jz0KsOB/3i8ASHF68kgwJyY0Ssax5cfP4d1
dndC2rFUFqcB+lVc9UB01VN7P9Q/aRZy9LyXGBombh1yCklC70cnQk1UN9BBKrN61S7X4zzKP48T
oQt/aZg5LymlhlRmpuPvJLG2Ehj0aZYnY5Eqhl/0ky271II2FZPsUIt3k79Rv0Wnsrh3BnhSq/dZ
IeJNYIh+G1hb8ud+/T0fVnRB0M4UVIBsIZLlvgKZ/xozYGfEZMggZM42g9d8/fIpbAxKqxN1/+23
4cLUQVr39DVLJJGr7VNXWT2/wJLilod7SJp8D2/loUoziLguWPwQ4yFFzN7mynClqssbMq2u/N73
st5nHMHH+wKRrqGgJ9EJJLD/IvRuibkiqAJAfy02pelq0nDr6tlhuzcn0ZM7HRYiXvqHE+uPKLpB
BT1T29dqwudvV9/dToQ6zQBoo/ZQdnhwwQh0W9IU3cUDsyJW7RQRbcIDYwhFgWJ2QSNP8/PX2c+X
mI0zNhLAe0ir0Qlmsde9UnEn5iE4hdEML0d16JAEHAJLJaBBvwHsi06bGbUST50KMMMg+pZSBeng
lW1pRg9fBsN3rMpGKoK/QU5Ig1FlWj4VWVpG3Ey2HhTmXMQH6Q6gAALY0kXtfZR4hv//nwhv37JA
m5GDJFgOXJChSBiyHWoTG9a4UPBlHew1c/fQLkQf7RdITcUaxwCDxy6wxiewxDr8eRXgAPf7VyM6
bX4TwLd4/PF1pPZBtV6f4HO/f6uypWj/Dn5vfeozV9nKbT8JBg3H0jx0m2q57bnSme5zM8+00v9D
QPQUlMr2LbgOu10wobyGvqq/9gXZBXGbVSbVfI8k8MJoecm9LEaDi7Kgjb5tGRoR0vJqm7qUfKmX
40TDx7YmNO8m4Z88TJ8TaFDvxU6uWzn6dVmiw3HIiqS0K3iDlqj2VQqIbFRX/EL6OkVnYO+DKDxa
mujbHcUqkcNwULNg+W10eN1BpNSVUgnjwLOdRWG66KI+TBPI/yW2QEgVEeBIO3iH2QnsXxFNI01C
pxk4mcWN2e/H4f4sMYLUNCW9zOwd69LBmuKIYKZNg++ppJluh/rbuRzPdFw1QWO+yd1sfDCJ8Bkp
WCUxKvZaLP9aaGI1thb/fqpPH/C3KOofnNJpNdDT25Huf4U3ujoGy4OkDTyPgOcj3GY2QNn+C4q7
2LBNDPi6OOJ9oucmsAOWY6jI2DvZCLifFrkGIa4gbnTAzNDVN5qPDNE0noONlHCrJbL9bJJmmeOu
1Kiq5dph2CQglocfxnzPd9GTwC2zBpzGYxcOyYbOp0MJvcyaFyrlLjXwmVUP5ReDyjoO99ra0D7d
qVqGqH0PVFZhz0QumXnrpejiDIMAcJ+2fnza6p8nyJyr2Cgtn9MHwJ8dpc7PyKQG1WSTJco+7cu0
64I/Bd90HZSughi7bkCCegNOQT9/uwTE/LWcaIJ4GyumCiHHaW4XTY/IAItb8BwWzZfCss7QQvcy
XW+JC3vBwB7hc83kur9kkzvEKHRq0F5TywgT78hE5JOjOyHbWNbYPbfo4yc/L1uJm4eSUWCcWkUv
i93aye1Wl5GFy1CvNF98PnabYx/5LLejlp+CUxxaw+TS3o/P0sRKn+ykbiYG/XvaDWJPOLD/ysmn
kGms3UYUq7IgyzFUMrWmpaXyBUsWUcKzk4HQXLWBM4+P1HX4CfJaECK7jdH/zUkVerxZDjD2ey8G
rDqsEmL/vTjhxZHWT+01NXAclhtp9WDq0j7YgbU1MI7aEG+Beh9kgRABV4PXdEj2FaVlYT7pIxGN
OK6NF64RMDNfOafWx2B0W+vfddL/i4XHAL28YWA8RBVKWYtMi7iBKOKa5Zf5SjGgX8RAkvZ+81Xe
3gAQsZVcQtY1A+vQUvBfyIG5SyaOE8l/Hcub5pb09ePHsMgvaxGqSVD3wvCMs3eLswCFBA3gpZDt
yVy0h/ke/zqgGGQC6KsIJkjEHgaPlefPPOlPWcwjCT0d3MCmO5Bjxy9jYdwbs/SaiBA8yrc995Xi
BzP2bPJue1mY28FR2Xee4Jn3E9/mxLuLreQHZ9WepvZX6jJWbPqYx2GoCCAZhXGjJmftgU3xwYP2
SFZeuERKQAnwfNZM1WL39Ps96o4wEbffjLVtNNRGG9wZ5mp6CnYWNKiPDJ5wwtmHT7eSfUxqmF53
q26f38rmqKKKL8lPQUiGp4TDbYZabq+pDCJiZ4MEU1rw0rzbRNiDQW5kbAFXKukQNy7WuP3u1RsA
AJoYsWiQFUx58pTQbUjDZX2C4UWisP7hUvJ8l7gZc8WtmpO+vnErZcFZzv0HhN2rZG8MmCAy3Q3V
aQCGwWiDzoeoB2QafHl4n96GF1QwX76FmDEzVYdP3qlw4PkohIcP7PnZxATjYTu1QuxSZmMr07eT
s5cuajQ+S1tMahG2Qfox2MS693J+qiTc0zZWMwk+RfO0Cc+O9MTW5AdwqtaN+JNyDtjCeyIGjfdP
UzWif7GuzlDgUgJ8AlbWxQvrtLdPh0gEYv0vH2PkGbDSo4YtEYIssle47yi88ino/YOQnvLuPrq3
BNhB4uc43ZVpPgIMX7Xlqtm4xEo7i4+QrNU0y5JA7ygqdSnPj98ZeS3ebc0EU26ZlCOZmM5FTphP
v4pXOapg+Vj8dB6bteOH+/b2KkSuOoFPg3I1+StibCtdpHic/eLlOuT8Sajt7Iu1TUu6OO3+kxXO
+LPlY3ORjdcZuscHo1X6hgKfWVCDtFbF20lYa3Akt/7kLIFAiDlc+bCmuZyAl+00DTGDmIBvTr/b
+4MD+46ApSYv0q3mhefqaU1qnKaWCXUDeiRqsvFBDkFrySpZ5MgPbMz+HjRLCswXgbP7/b5TAbA/
tjh0J/uwRVNeL3QbPP3MR/+k+DPiQoC7ii51F7myZmSAURwpQq3dtd8I8x0aXwj2NWD0wrCsb38X
/Yhg+xrkabub0h9cmtWigwGrqNVJWMZq4J2Op+9vDYT4Ww6kmc3moRCtWqabpWOsoH+golWmA1J9
kztAJoLCIjpyTRKm/Cn95ZWgu/pCsN4WtdBLC2A2dpNWTEyM/t0jDG3FBMK4pSCk6WNO9hbNcqwG
mSetVIaCS5mOtHLqBA9WW/mZ+Po1bnrQwYkRJfWvbp9QWhgnTDGxaBU36Xp20x2gJgWcXLbWsc0b
IKgnd8w0Ti8P6bNkMMCvOoPmyqp1fmcO60AvxzHNltlmhidHM1d+KPsBabxJPw4j+RG24AeA1JsC
ngF0ngciaXBnqozBg2W7N5LihbQ6JJ7BrCC2565Lq9TvrwCHHx/QO1buuxLrVzAj59QKT7VNr9UE
i+EFJoQGW55vU64wF/OaR3pfMMeNlSNJAP2Br2pvR8VykLiTs1Sg2dD2M4zK+m7MeifDL56OYsJM
StDM4LlFO3EjMrJBslj5Sd2UEWZ568iU9kFt799A8etGiNPpXl8NoOED6c7wi2ZF8itvnqC/c/GW
RT767AEY03EyyuNMwlrvmMIZU+b2EyQxo3FnH3XqxhwmYgnYq83uRLVJNXBWp7yPv+4/et0PzJCi
8+1zlVejpm9FMExC9IuJMPrWIhjPBJeCVX1nMPjEyggiCrL+4wfe0sG+/b1ylDeLhD796VdYLXrN
kQmbwii11Qpnz/lAbxR2gJ4C7LuyWQ8sH4nnmEaFOxZf0tsIjL1oWm3ier4T5xOY9ng9vW1e+uN2
IcoViVFOW+7Wyff4oNYYgHAWy6F2UFB/hXuAWxD9IaPohlXorWZ+K4aUUoDzevyi2fMWbkgWAsO0
6PZciwptxQ4O0cjzgpaF65FvRW+kxbN6qlWhY527NTPTire/GoEGjFZO3lX7iKUy5JWm87ZXP0l1
SVRQJHtvGBpsVQRsdSaXJGU1tJ3atCWqadS/CJl92rAKTwI+Efgmj3w+pCt+uphRBv/YMVpZDV58
G99ZgklOaZaZI65xT7n7BxsafubaM42SNww9FxXrzAQKa9vJUEM0QStz0JLszFzyYcIPs0ohoPW0
dw6K+p6mqUWAOuFa+xGLLawoS+22WcB7zS/btaEodGTH0q3sLXUi2JyqWOKv+nghU2TZWyOIHvt7
pNF+mPxYwgZj2/cJjD9hJBiYxwUsb5JU/F6CLd4CDb/lmJX1UcJhtmM7xUROCKw4PBxeSdJDAczC
N4ldx41ZbrxjqJfc8NeWJbkcnFaTbSgxLZZfy2odtrSnVV3E4H3a3/R1vYlp50br5fJG7ilSuDzm
PiFMy32qxZqJYDcvn84fOAcmkjEjV30CACh4G4PVlsrYzycgBr/uQuQdak/7bRNI54pR004DjFPh
LaqIpIg+gPaeHy+h1gHugOlOQNMQ4XqoRjHAmRMIUPV62oJxBgrlchcwpCYXrPSMo8GnaM7MAafO
zHYLXrZnOdTxfDosryhOA/oPEPtq1fp3ixkW1tGmo6pqKLCkUzJC6xWhzHG6qJ/EowtmZU5+DiSr
sstUV4TR//WF7G8eJJwhauxz1FnnCsrHYx+yDUd7NkUwYYCMrAJPhojS68UjXEeFCjMqddKR2RIr
IP8dwiEpZ6EXcwdK9UDwKcS8vzuDHCG6IamZAHLiGB3W0V4oH8cvSOBGc3FKNLbiqBvbBiIihx6z
7Mzce025BRAvORQKhF8K4bUmLs7gFlP0AV7d6tN1OJErpN+ctURp8oxJlXgF4QGi7t6VnpTEJx56
JvLhIDdmdMzU8M+7VaVVGXcPoyaG09EunYMnOxtX600j7THh9HR1XHOZZtK12zcopYahjUtW/RTU
OJcE6QVTFfHjILcCPVL/4q+Y7e6j7OMb1t7xsLbc43yAcwYA2juIC9gn9dfL0WIUp3p8Juuu0NzW
SiiY9FK5eNiEZj/1F9/L2q8HnRqOeyOP8fSS5ZsZsAAMyXlc05kxaADniuIciY8m6PVXkpKXxo74
KNExavqCV+C0FwMQpkhTkD7uEmoX7b2971Gead/shLwQsbOAHiVWMf6XxiBRSw9rzKLxb/Rhgrxe
OWKvbfwJUx7thWAsodaYjnfpoUb7KshG+t1/DpcEOyxp/71ToDXNi4mEGGhWnX8aT0l5OKvNW6f7
xwdNYhsXw3Emhzz9m7x8+ml0ohmswd7wp5/Sin5T4xhCbz7mpcHIojfWjjB5OTJYXvUuSYaDPRLw
88LrGydgvEmwi/UGQMrYVXnrENENYwqkIz9STxmj8xZX7AIYZRoIFTVHuiUacuLpb8HM4zq0vgtG
Xocvdo6rnW9IDaobxC198RnJlRTVNGrBYSd4Yp5hQAjT2BflzU5OPxLNkmb1Vj+MwnobxTpMT2QF
lUquOIWPx3EvS+slm1uQh1B0LbyBzHB+96a+rAVoCE7BOi3fJQk9uMQUk+NDviFOE4SNbieXdS4u
VCgWW0kKYLJwPAgRtwsEffWrkf7l9/eyCFxUN+pbKeQ8wl7GYRniJ1Gng21Jn+4KYw2NCHdEZZlX
444mTsY+si+EHKUWxGft9TDh+pDdvJHRhuK486F9ubtadas88nkq9xsGkq2mIbu+6Kdh1w+p7Abf
5LIVafYBlHEyUmQkbMOsYyKK0f7ngWJtBqUQHhKLnxMmnbgpdN4v3kr5uwB016FKV6K5ksUqLVgz
ZInC3xXmnOAXlNcGUV1VqUcrAjqWEn5EtqSADboYOZjfhmA91Gdn0QT6CQYt47XYowqb6j/hH5gH
C9ljdYkAjCksomHW3gNomgF9EUumhSDQLSfddxkxY1Bh6aBdkK+7cLqcPkdgf96nGW2HwV0DSrrs
LYxp8B1wPE52ctwv5ehoErAD1wuG1e9GoalaRq4nkhbk9FYcZuA6Jplinuua5bsYP/KoenvEpMsF
oi/jPty9PYV2CmNuapegoOs0cLpp0QtFrK9fxAyf3duB0Rchk2DXrnvk5vLmH756o9rGHPmJHzQt
QBR5lNuHDa0PHb+0HKvfb432wFkq39o3FRqtwx8+QcaK7iyIrwBQduqxsbLLc6OeDj1hum1MalNH
HZzG5LDvn9GHdEMNUYxAySLZz8uBA+ctcKNB/tpT0HE7v4ECnCJDOOoK/MPp8r4Qpj5GY41bL1z5
2804txW9jCrwmrFWBHeTgy9+8Ct0y2oKxcSa+hqdOswbhTnHhw/ZN07z72UIyS4533LdvA8ssoV/
jvc6kvHCf65ljLJIjbING6O0JTPDYdMv//p8zKffOCr0DGL3LLNLJ5NQkf33+Kq3RcvprM2uMV8t
USJU9E4+QuzqC9xkeg7FSlpHYtgIDKpZitrsaieNfmVwZYErbVJrccSNno5jT+2WLN5jxXpSc+vP
DvNIncF5gxcEQr6EDpByTuts4ICSuDaXZHjnwZx4Lcqaxc+4qj4ihDDcwD2DH7jvnYHAPkOfUWNi
dfZDZ5Lep+VOjQcKFtv/L8VqiI2yCxVTPzI9VXYcamSIkPKdxF+3oUTsXySx8Yg8Q1f0JtT4wfom
3N0MCEmd9cA3LF1yhtNY2bbJWu9jJrfE5pDhuI99kAuFSICu9NxtZGb+Ih0Qq4nXF6hPvsgj+Iv9
EHlnD1H9DdCx5mkqUQj6epPGGXVmx7aAcHSfZScOSJ4DT9SqVtZKx3hyfLrqlmIkePwvmAmds0+c
XeDoQCNeUyloireCMAJ15hQFz9dM/0r0NNo0gT7EnJXHAAxZ2N7wMyoAgoQ/TFexCsQc6OPlQaW1
Fp6aWZf9N1ESZoTh9ATw4RdXD5AdTBvwiTl3i5648UFC3+r22FlzjYpAzWRxKfRaOe3bnwa5gVhT
jYXr4E3K+7NUkPoA0mja89z1pD/usrS8d9aQhLUUXDa6+szLx8BCN5GWmaFlP68CGSeNOVJGPneT
cAg04NlLtu6WANdhNZ1vce8FndgU+AuKU05W3kjuU6UN0Z3tq44efcFlhx+63ixwEBNBhQjgurIC
h29DduxVNle9zD9oqYrIb85+Ipb/TJtQBiLZo3mEgFZg3Qsn2uDUDwe12BtAEJgBFBnXuZ/GiGgp
QvlvxBJbegXdkfy6okjJbvsFjCVgqvWK8/R/7N4FmkHqiQcXlBx3/UDi/PuHX8wfchx3ChNsOt9i
O+OAygVbEMKiuinmi3EwK9pOiBeiG/fV1wLtnQQl0OV9GaoilMnL99zR8ffUNRH+bwdmcv0oMoTL
GA8HD7wnkD7HsV8Ddg8i+90v7b09wyJicgIgMLJJ6CqBJBsNIRX3pcEgWcnfeEIy1kyqsO+yNzOo
RamjjrWIusFfv6Ct5fJffRA7EYIHcFF0oXxGQ7c+BYt3UaL8sf94KuOCZwa8+QXl7/mbYKU0lq21
6ghIB+jDGy4w9pKlpn9x7pdbXoFLWVDnFQQejff4gbIXS8mUvGhTjuyAyWh1EhuGZQAWPjLsuKyN
9zqhr1XF9r5JslSiB4qOTVR736ChkE+XCPelu9C0BUuKOzlgmwUaCJNXLzRRZBrYVZRj5A9NBy0f
CqI7gXobc/6GHeIj3HYJJ53Oq1DngYosn6xiZhBQAhMQHFiR03SLO8xUWztS38FZNAJ71g1UIRkH
42K9KU7lWV7EqynSmL/jb+41J1NmS6qaJbHusUTWheR9mFPzNz1m/yOdohlWQFfJSnjTDd+/oH+w
64aV3/GwuFYMcl+rCC9YhlfqYTUePcueXhDQi9ACdT9HgeUrMRLhiIXu4/+3XiUyefUJH7Io/Q8i
XqbfHvC94ZjWmI5otsAkt736VtQdXddaM6NJfAC/SCkexjLHsiZehp/N4zRNmQZ8JYDmNSU6gbFg
BgqvU+t3EpXMPAafzbE2bbFPTw5k9fPd7o4XO0M9UUmtsiq+TmaanRQ0pyeERwgyq4jzEaCflcvR
gsf/ibk+zTt/QaUrCRaTO3NWuZ7hgmyem//L1VldSpv8vDK9c0/SEFGf9UGMFXZOs4cXBJTfV40s
kurARGfdoBFH9HtiXADdC1c9geET22KMN+Kd+1Vk+aGwXwDC6/dfICaSyJP/F3kjjP+93xbAdBSE
UhDr89tMnB+PKSkzl9OSMJPra286+Eo0MiyRNKV2c5Xu1vekK4k80UagS7m941hObwlwSCBlftH5
k4o+ZWziinmmKLP1GIbmM/HyZGbhTIRlXfYlgfXskZ6FJ6ypuxog9Rp0PXwCMKSz+6yZx49iwsJA
JDo5vIfGDJ3G1gyl+h+wKhhPQ3BaxVavfcrTkwbR4CHMUwZSZrvMi96SXWRQDuhh0Ux28pp7ppwq
X8mSG6qRcQHZprD9grfNDJ4B5mC43tUiOMceAfbJnTCUVTZizV+BjrXsJTMxKP1SriZfH9FJpJcR
MyvAESMvpRRx+ef98BWZGMRMTStp3dejHII7qq0v556ye1OQYZOq3ALr1eT9H/EGOEKLEmTAkQ2N
DGBTQef4Q6lTdz8noS4I4f7c+GDNixnI6l3y4rYgFCGNNZX2MZWE6mxw9dtI+kTjRasycaE8bk32
0sZj0s1VdJb1d++GW8p2QqUul4PZyf08VZgYu0wjl9hBk094kkMc5E7YadwR3N6oF1PkpEd77EXo
FKnnc+hhGCw+cjeMcKEX7hvbCsTYdcSHAZyJ+pTNgfF/p/icuLYP1oWrGT8Is0h3y8Yk9xjA6G2O
uUF40tV6BgSPNeUwVxeRNf5FrTxHNuw84Hc74EIqcdhYdZrmL2oAp0PB4vlaHkrhOsXGX+BbEgGn
Qp1iqcH5V/YYvjJCikzH42X8ynhEQ9IVI1mqTQeVedTHBFZ10FGbb9uXrOnpEQ/PxFE4BP0QSTN0
GZqTSEjbdTgOVyn6TI9asSygNlN3blzaSXKUIP+QNRwpaH/DNofT15mcxEWOPetUFrV6Q+TjLUzi
7LjQYc4bu+vmw9dggQW2k65UYLAn9eKNMiZj6PKjGpy410ECMffOA+PIK4UmuLquUf3pZXJcOG/h
Xm1KB3bq//xE9g4eR/dZB03yUr5hlImddKt/IpxeDnl9ylcZvfmm75IrWAAgFx/h428GfNMpLyUj
nAyQaGBrdx6U7+kWlV/ignix9UhuRF4PlIaua1qkKnqKx8i6y30qBZgSS+70KRau1n58paN4NoSG
3U1eSaV5ewaB09XNtGvS2hN/4jDSYLhz1AwNkeiP51eh2UTi01I4gCCh9ChRG0HQz6fKii+WesXo
utVYa/09mJy//z7yv6HsMNvmB4svarszaN5YoBiBTQdrls4aUi/N5Ljp+OygnRqWJc9RsNegEWkA
h4EvjU0zZTdumNAVtKEmWyrN01vL/rdtxNEOhu15iV9Oi/YPHwc+W8/m15wnTTZ/b3pkdaPTdw5a
2HaQ+MEyeW2mqqR3RhevrK/i0gY/7SAXa4pEIxhuETpdnINnUeMpJESbp2kwS+xweTOXPIbzg/5o
uCRzK8AX0KahpW0wAjtfOdSgvKytjTMkYNMoySCyB1pN9gL1ECiBiAAaehv7W2afbDAhs6FVu6Mh
qWa9Me+/c1JS54VYWeZR4eNeTbf4QtCw7l5sy4wzTTmu3k/Pe3/zKppkjwL82gzAJf8lGl7nwcN2
rrgYdjS67dhrsiYOj2ah0vilIbANK1RvtI/4DIsUUFJDAiNnVFDyc0JMS7PWpt3NrS79CHoxWRb3
jRo8rW87S6r/6F51mEBeD/7vaGlNROTIAExxkc922HpbonyXplME4U54g0xVtg4yaFzwq727jk7p
EJxg0E42LbkvTuNt2eTy3KySKswT0JYPZZcgN78Tv9xZL6VqQzqjZQxb2WKEPQYqCLr7uEsk63Hw
7dxE2pQHWp+MeytH9aKgQAhXhU9xchrK7F67/aLvqRbkOgEKVR4dZmb0UalqkZUc0Uw6sPjpqtfj
3nfLGCjgcxuY1lj7KTgebQ5mR/TQOf5AjqnfvGqWBuWGlbRtFwc3yqNjQS4atAAZ5k6kBbWuSL5a
+lhoLMHY+smqmQU8u5fZEQec/gXk8xgrYIMiuaBERauit6vDAp1eX2zEYwCYBi3TgkU1wLs2R2OU
U4ShV7jTB6qsBdMU5oMfJJTqanHdWb7a+a0vmL2ifar01pt7qmUey/DAUS5k56u4UARBq3SeE2xL
4TsWybkGY3a5qFXHbVseo86x6A8Ocd/86nXUm6SoHcyK/UuDB6owEpsFl6VUqps4smT7q8s01Qmc
PItlaBNefIrXVHDVNqKiZhfy4Ragkf7gKGKA+KpqD0YG5kKaJeN665pOLpNSvqKwJnvhX/4h9bJ4
mZfLC3KevnnI2+0bvbKVTQ8VWYAbbIi2qGRFDYPE+UGvyiTuKHY1rPimGxEqxFEAEmTH4A9Vgge4
ctgDmkwr+lL0JpkTu6RyH+wyzzzeq6LuwLTBMf3yGslgoJmg/WXpIe1YVykDUHKrUFnWPCO/Vo3o
s5znrfisdsSvZVGbwNYqJwvZmk45gK4DzI11W56mKTR/TqrlvujzpxuI761apbNBHSqLhqoJFf27
bK01QmOrS13ASMnOablwuHwB3O6wDQ6TwXHE7GvndxtUFPBRVPpQDqSh00RV7nMVY3X/178NfBv7
PBjqOtYFI7of8H3kF9/ROZQywDuVjfioxUnwTwHiyS9+XDE2/RKT4L4mMQ+ODsuANk2vdFvZHyua
p/ySmO5d6AkzLOAFeiLkSLa9hR5hhAqCRxhOW3ls8mTu2s00v+2uw7n6rC3AOwZv3ymXe8C7zSOl
TZxJ2FldjUn2yibY8mOwTnKbYFAJlCXk4dz70kkWtEDNcFelV/izLvYOFQ97ZoXt7X/KyxlSD/Tl
LvtSOHTXgvDT027mkyL3VJrYTmSA5qCjoWAv944vc7dhgdYHFMmp4DvHqavfzTnQr6SH5o9E9MXC
+s3vGwNFxzWkXcSfUeV8d/djC+Hf9HVnlikS5gfYT/EwJnkXkoZ80hZr/tb/BMsuihJ2VSGIeKyM
uJ6/EbXbFfWvxarXkr9nUm0BUKnR35p2HZC9JAuSlHuzggTfHuVoSNXFs+k3D7q2bJFW7YnZmbdl
9IXFc4S/y9RJXXFKeU5OkZ1gx6Nu6Xo4G4GHgAwO+JjAl8GWaG6QSWFvodD/yXtTcMfbEe2/srp5
HgFCcj605/LSVDzu7/+Cfp7H8RgDUBCYxVNqWUHKH/7nMEqsre7zn1vDedk/6UBTf8Z1QNiYkYJs
DYSJKgB64droY9M+4NiGGzxPw8zqaRpxobO5fzaQwxzMVjq4anuYFLLwEbzyH6uCuxkzoQf86eAR
AD+0X3MTnVoUmlpqToiIKsWZK84ecZIbcM4ewq+ac1KQ4r3JJUSj3bCWXeUsK3gBnudr76556rv8
XzWrj6FtnvG+zvbncqYFiBWJnqZvMy7L3ZHol4bWv3W/or4BXgjxs7j0VvsxlDjr2SHq1uPclNMk
5py9ULy+ciBE5FP4tmtxOBHud1TYkxzXUPcd7bU1/YARg3I0Qdts/8uH/S7hGfnD7+Itoej7dQH+
CDRG3WfoBaYVx/lYoMrwnVFJk3iLjeJhmdY0KlvacVbcLWM32bfB4Ji2KKL7H6ai+aPRsiwbWqiL
L+rHjuiEPQQXV8vcXZBuhjBvDlyeARQliipCQmo0KW5sdKCSpLou4X1D1FxmDKBPezbuKunixxHA
wB3cgnx7Q5HU1tB8hF2oy+Q2HTeCLZyZ5+UmGSVik3zsSdwDy9b3zpFue074U+/nO9HkA9RgYKYi
xwYjrKnURbPJFn+HV/x6UYXFQQC1cj3C4mM1OXlKcYlwDiLIgNwGDSgPcIraOYTDG2ubGm3oT6SW
ZllkvWd63pQ3yih1cYWSl8DlsRTDsTpYtgY0maCEriaZ5Hn/7nhYhMPuYzLFh/gllZeCtFpM2iMj
Crd564ESQ9YvYBq5J8SQpiq/w6u7Wrq7u3dBEn4bjOjelF8A20K0IRxjqD30jX2mGj/evKkNdKU9
P2G2SGrDKw6xZBddKeKfh6nvIdRaP+0AYRckIofU9I8Zytk5U6em77rbAhm6C8nJG7LjcRRjq85Y
gFPUwOxfMXksRtHbBNbJ7mEpRymRcLm0iGQacBJyoutNDaXfxPVVh9wBOchV3CQbGX6WecHHo5Bz
nWx/2GMNv3uhGGIYz4S00fGnBUyQjEcBv7OiYyzLvhTFn0sfQ2+O5mrc9zcPafV863A/Rodd803T
f0YAv6jLm88vqZB6MrVuOef7Cb6JTKOYSTU1/dSgD548bJ0xeWxtpmdlLFlBxRgLEnZYX/xQKfH5
D0WTWal6bvUyYxOiNrkqLjoNwZpz8Vd0hl+6GZkiRL82B5z9shFngIoRbLAn/+ra6hU7HiSgpCzJ
960QmcPucBFUvv7k40R22+XXRO4WFfQCi1UKZPqNiMj5AYrzjmE1WSqZ4Tk4wKeM50vz0m/m9xyz
bHxJUcTs3v1lSK7WiPcOZ0ykPAA+/7jZLcc6gVy5Li/zX6NFDSYhK1RhvxyuR5slHbuIC9GE6H48
io/r/7Rqv5Bjs4n5eP6tGiQqkgh5N2RrVDVj5mVNMQR5KlKmzSUDLRMVV4hVndBN8z9iSop0Getx
BH+wy1TQD40AWf9N9TEDxbH+obxPRsPJr379vERuND+ffCe0KFTrt2aANRnfiqUm2XRUf3WHkdmv
RwzYufqiiqOK3IXrG6XvV47Fb6TcJueNk8lTxrG1/6Tvz+X8xIw9KdIG6Jl9ZC/TuOkpWB3bNLOS
CXrvdtQWMom2g6i2cK2DfHme5/jwhWcvcvkY1Y57ledYS9mewvp2Q92JWYNvT73tqC/Ce4TR75qU
wWXhebv28p9VxlN8gJJIDxOPK95YXGDXGw7wbCwtHa86eMu42HqECC0dz/t+GqV3W/YOneutL8c/
722YTIWIh68NLZ7SJ0coytNjpJX1egOFDqHrXs7YGLk50mvKQccSbV1iq6A8jDnicK61vv7vRApd
1NK93XcP2aAJyLYMW/7Kk/K7gbmLzOFAKwUfNylwPzIb3y0ikX3QtyJkqOyKqLdgwiriP/z/eaU0
sRfv0oZiJZbmJqyxO7FEeBfMAfBDmpBtwbwv9XRmInW/3Tb7sehY66nTeCU3OXGmvmWxkmsYrXN/
5FxQjobLVsAaHi4+DnCFXM0pJ+N3aSNUaVQsmuEzWPkrEj4AsAosVDtZHCGlMpp0RQHeKnJUqhxm
xOEY7TO488Vcxay/2nRqnmJS+Cuk52QxjxYBbNnp8XMw+5iX44ifLgDLfh/o99NrCz/WoAtn7sdg
V83fm5Yl00/WziNmvYOTyCXpXDUbWwRj5vxpLqcx4dH8zRG76cuMYJya7kqWYfc7AS9poBpl+lYq
YE19UoA9ZqGWL7qX2wgNwsmoaWXLuNUXu9evm8/BiUnB2x5ahCENapl3d/BmKjZHNwFvEkbtGtIR
YCwJS+ya08gBVqOdw/Dw7BS+uV4ypl8R3Gzqx1TNpzYmSJ1iVcPavb1I6+wiLv97tX0hTsaZDYCm
n/CWE9C/18w5A4j/o1lNgJpmfTkwduqlhv/384hx1TOSsNacJCcGOafy62DV+sl8t45FO2HCR3Hq
MzlazKWQKhaM7iwSY0D0VtWMoT+61v72mfwB2Jr2fXNFAdX3AMgBHr6RfcaRXcyKwy5yIEwZj+1k
EdNoxQPCTVSjsPWP91F5shlhXA+Pj5bdfR3JJxB4/BZU1quxL+VVRpVAkQPoVvieSDEZ+iPVgZii
v90stHSDqGtrE4ZcZx06665JBj6C8p3XUipPjb4pG+v4E/zyiSljCn5ZIkqhV/+LiIS37t7NoRn/
OFe8YQxFg4IN6CH5sBmw9B0gVvqYIgCoVScHGVzb4jZzPdKOCamqw+Ns3teflsnbcviz5EWNDWv5
ziW4Jj6ff5BA8g8eih83tEZlvMI6mIrT+dkvoHucTZv4QBRffKPgPvNq5vDaLl7tux2LzYVKNUno
ULhWp6bTmJGP+KmdJgKMpUD1OSFOQCQtVKHUA5rsSzNdPES3oA1Mv5HvY388s9kR8WUmEzt3/quN
bXzaWqCHrHgn7fTQTngnBrFyWIXicnQdsbytskLUMTTYgLur/gZD7hzKo2uJXSpuqPmjQeKDLlcB
s9sjj88SaRvEKoUYwx//yrc2jit13Gxq3xhiLR2EVGWTuK1+HGibGPnBaibwZG/YfJMtYfEZ8++l
KQ7digKhXy+ldS6vE4osmbbVk7i23jDDticVyBT5rwM0QMcS2+yRJ3FU0U7BdCbPffXM9uCfLe3j
itukqSIIvxdIalE9uNUPTD247dd8L3xM0YcEdmbqe66V6DE5oVg0NaqPU8o7yvTnNPH4bUkNvY98
7eTkh2Uazjo0CTrcw0DKxKsBE23E7eagv14sz446il0OwKaG0AYehlSDQ9pa10wqGlsEZSFOiTnr
K7cxJy2PYhXeg0TUtieOvhpstCtjRJd/O3kIU/thoaaDYNCpPJQaNAGnvy82OJVRENBXlvEphTiU
lU8tHIB/39z9YZhgthS7bcGj6kPna7lEILDR348483h1nO7Kpek4qU2HwKT0IJo6mML8l7JnQYk1
MVZ/wCvaRYSUQI6Y7+tot9OH+oRjDORY3M9F8Aeq+LRXAW6/+BBzlYrM2ZMwzqtQaloT3QLYbSzb
fyC7NCMUt+n5FGxTGpESELU1hBkC2vtZLG66MH0ZqwQxGchF+DujdqWdfLRoW8rZ81lgDpLd7XEu
b7jK74/SvQ1cdnwmjLW0VzDCBTutqUza46pzq3WCnKI5HtbSJ+OOjoTJGnchurguNsFsIagOa2RD
W0cbzRoWfTV21edRarKrC8CijN3t4svDSZsdNeQj3m/OhdkJDDrbGs20Jr9kMvadYAj7FUhk67eV
KK9UhEimkMAbCGkTzUMM9ECPp/liQimZ6QMbrec3rwEEQVZrIMQ5BHRjriuWxV8XVbqTdl6UTMia
hfHBa+JnHzT6c/xdcYXRyZ5Ve4bsSXW1YWnXiZvxoiRPVwGxnO6MA5RySEvHAgIw231Yjdtrws2N
v+wfUPU86Cpm02+MkcyOy40I7p+3KO0M/qwMLVvQCHjcsZarFaVvk0ViTtqDlP7D1IQrRcvP5V2B
CxWaKNj+aMtPLqtzXJVwaGCI4d2OwhP3ewAl4UjkfoV7zdAuSTbTLEZhvrKArjv/rjHx/JbOygLJ
0g9K8LNXvSsefHxnNCDRPJf8x3Pf/yBFnihye9NUbgPrL3xwKjJ9u5JWiH9TiqCY627/g0xLkCrm
xLZHZQsZi1LXAKwZvH0LNj3Aq/Xeu6koa7qiYNE2E1i+w9myNR1kEAMr++AZg8EvlhMkoz21ro2P
B5XixyooZKjfzhpJZ6ZSFCMRfXVlwSMNLi3ZBbCMd0YMBjonAG7Jf/PkIvITepevdLk01mQvrhUO
I6DB3s9A2btek8vT3ZMrEwfSrN9ImXfrDbw3eu4VmtGYlD5sWHKaM1Wa69sBIG+127rGq3OvutSh
Nz643mwmsVP0vnBBhZ8vpe1J7j2+4xhD66dauAG0theknooI9bSb677OFTJu8EHKpYGgqFi34SwG
GI5w0pp4/xqIkcFHNAn24q6JLAWwfY78mfwt8Yx8bRJrH523UnlC6krbHvr+TkHuKqRRDt4hmKw4
KjP463QVtNNdNwYGG8PR9m5LghbAM9g0gQS3sgcIp1QLDfuVY0WaXjF78c4ujEEDON2x3RtAjon3
uHp7QBcqhEeigkqM80KD9qrU1DZXqBK1T3BvgSn4n9wZVTT8L4bQ7oQhEzPibeZ0KAufbDFFI0VO
CWzDODgS2JWWMEmNnV+ROkXuCMYFyc9uTFPMpMyEwVtcSvQQBJSZTpwykQI8YTFzHPt+jSNP15zu
L1g+0DzlH72DOE0GFuWepsixTV/K3MspCZnsJ4bIlCngY/CE27YfBTQn2mLUvGDVScCJV+xRgBjE
RCYBeCPyv8trX4eBxs1dbb3kEPfFEPmdiu/oUb69VrHb+Dfyv+vXn/S3EqgMiTOaj06OFk+dF7n2
lRTOKJCbq7yqZUkOG8+U3byIDJz4botgsTfTpmvmMSsrksdgoWbf+HO0Pi2cpXZ/uDA1H3CCybl5
SJKCyqSgGv5StBuM2Y3HnW0mo5hIootv6gsOVYWfFYuvXa6hlQQVh4tFG34h1lVJB3W6I/nEVLcb
GJdHIvtfYt2aUUCpZtimDhIEndMz1WyjBQznAqGGe0dWmnC1eJoRU8vclGanLYMkTgfRXNHNqfXR
PFMlNiXcRxhdwzx8dhgC7rA9F/z0t+gHc29f3w+5sDZTxha2AW7dUkguovPzI3GqKCMNyCg4UVh5
5olNYwll3yLvhPoBj9AXx0d/SDpdnxaQw8xcB7WFFFW2oSNbhAfL9mCAm/kifMz3ld9P5ojPOyFA
cMCIdh0DFAU+qNWKtr8oBrctJGWhWGMcX0OBrAsna45D0IED58brkvixpg70x/+UzUZryFrWQx9v
JnYZ1gA3QJfLebU0kIcRQIi48E8dynVXBaIuOBOGNdVE807shVlCGeXbuWKN1mysLHQr2sA4Le/t
TwqufGsTMv47s8CiWLV9L+1kJvpXDVS1ykvyV0AMcE1DZEewR3K86PuK8VaXkBckIfubm419tsUj
/okEZBASLW9E1E2AAhMOkPwNKjdKefYpwSJg4Er1h6Nc5QCXVXmmPH7m8BZYj9ZzUnyH5MOzl4OC
U7qxeR3YB/1mfnmhmPgMgEZjljh5dHn2SIY7ZHZ5ymT5/PKx4E+EysoR+pCgytpHjgZVRgErFiBB
kcaUHhRkVYw6hFafsR0W9R4sFczbNMNTpgNEZhoJAODYM4i4GP/r5e9nIFAR7KEw3cLEm7n3O9Xo
7kSwiSSagkMid0KmjuFBCRxLCTH1JKBHV8FGADiPQZsoF7IHOhIX/Jc1qwVHyp8IwS9j4sqorsbk
I2N+MyX3KO8UuKIYN99zOxPAprETZ1GGYAFm6V6yb3kM9TSMol03QeIofX+4ZUGOY7BJrW1BX+7Y
JNYLeTNH/3SotIcludnLx5bm+n6Xyu3JQ0ZtlH5y3uTVgqO1AKmeLxrBZRiCnhBNjv+cNlrVBMqQ
g1hkoP35c1hDziHLzYbSl/ltgIy/YkyLvmh++eJKemAhPakn00hsXdPNnVWJQBg51QIUf7HMNLvf
kpKjrMykX6CkqU+pDK8Xvfb8bJHos3YYgy+lRNZ35TKrawqXq+mfAEAzQX3SunVEvTCr/5ASTXM0
jAeV0bVbGh3NSlwwEUKaaHLSJq7FicKr34vZqbhJv88gNX+QuVNoPQHq4V7PfGII4IQ0AFYOF46J
qNxAPCac5RTBfK0WsWzVM7+RDGnfPETNas80dZ2Ln8qDZKo2Bh8wob5o62Cw7Q3CsyXECh8G4dhK
ngCH5CrxUtth8FZEulaisw7UBKtjXTMj9D0YTc9TlMddiJ2r0n/FcId+MMpzvify3WzZUfJQ8F7e
vxdqMecVXCO+60gUa2ZxqOlGtjaAc1NK4qjNjL4DrXkK3Pd3Gkjy8IgSeTH8GSNhBYc2tMT0lz9/
wjI9hk10UdNg/HVNJfbjZs488Nx3LoS9O0PV4dVqgS8arQcdFjmF2xVQp0Eb3c2Fv9ZCOrHpkmRa
ZJvEYtjV6T+gik123Fo7pQQ6xRz7LWrD/Z/5IquS0ljmrysRCHAqyDsgj8iXlQNh4J4htUpv1NMi
IEkngK8569mWd52YYR6fqNp1CSeFgSUwev9gMZqpOlW/Eezft5K0ffvQnovqrFYoS/8o4m3HTAp9
vk9EpF9CWzoRj7shnHkaZ0Z9NcZBCBtGqQ+FfGqxCfKoHu7b2DbXsyq71BDFm4ZJACot5f6tXToW
HgJW4baXkQqodAjeeqlmhwg+57RrOhectXCQJb4QFnvvi0QUx/jli6k3kJFqKP/PCbsbX6ckb3cs
xCfgSfjYaBQAVbbm5B8WYlLckUADKhncdJLLAiRBpJA8F0/TlM0al6BBWAM7N/eq1NpbPR9ffbNJ
mZ+SAE5S7V0ubXkKcGaytKrMmQFInT27PerTNHy9zZhNEMVx58HH1sLe5nNWXvh4TMgSNZ7Zg0WG
XGeZNmX+WTVRbDi5vNTS+a4BxPgTY2i5WNIYbRHBcB+z+hL8EHPULS6sABxOXXEfDAOo9cMgwR3P
ECLAJDIS1c0uEKQm324UZZYzJtzX3i1Bgf+6YB0ba/MUIV1fYw/mMuSdoYFOzl0wyC7t8zb5gf00
IK3RNVHcTWGxgTbTlg9wSFuVb64qGQVliS8EG4fX4z74SixQCN3wIH2u+s6zj7MZluiBHFFN+Scf
Czqq50XiO9a6d9s+dBQQROOl1nvekS5H8/TvVyhQ0aUhzw8OJqp8zMmRIYGVVfkt6PQhkPD038Rw
Kt86JQyQuftm5NJfZ9nAOc92mxPCqAMpP0KrMZjX1pds4zaEb+5Y6dFd1kVzKusah/w4sgRawMmo
WAyYGhhPQHJ/Nz2Z2van5En4UkccS4MikbQ7CuCGuAhsWYviImIgKDraukzy6tyP+0r0bfP/+D1q
VG9tOGas3Lu8mpgmkrhDOhUCWRi1t/0bugcWfCbAMDnoOZ23N1oR10Z0lyh4vnTpBCijztRoTx8Y
0PCUG7dlKQUFIhyR72btMa51cp+iNS9Tiv6nJVXUsmsMVrXeoWlcf20aSxqvAdStuczT+vPob+LX
i+4eDJaawy9XrOygnWPdwWxDTfNQEWCaByav8/VBXEHJwrhjNg7XaHlApej9+JQ3nL3aPKmzyEVi
YGrHkyvykAELQzgNQ3HrFFs2v8EhkP+HLiMtb9PdZ62ruyPVsHTYoZPkGTcgh55Lr36WDrMH9FBm
V7/yZk3IJQbE0zWRKNmkODbigNIa9dUIwPPsYxtuVwNjRVbnOCIh27hCaQDOBY5iKZ2pnLw8kzhF
XeVQ/VEDCJTY6zfOMR0aPeSlz0Yg53Xzxh8a5CMUsGq3NGUI2cQ6wQwRTfXrN8F76DP+xTN5bDFb
nOyj3Z9Q8OUnvG+zzYVkFw72fIQfvv3sKA+d7PV8EDmsDekCT66OL3RM9w7g/MmxZC6y45XO/++s
9El26cTvkQa1R+yDOuRi5fPCA/30CRDH8XBE0pNTDSxyLw97WfKrwI32hcayr/ed5dTsU2GtwMj3
gKKbbupJIm3Z1pdJAHMuUPgAu0gX6M80DTZzoklQiLsITzZzp0+OrDWk8l52g2Hty9v/Q+skYIF6
mmkx8dbtqi9OmgSdH0lv38KiNg81vHYVXAbkwJa7oWXvkDcGlbHYhg99S91N7otdinwx3eXNVD5m
sdW343HVD0hUia/U8/r0ZppUwXgzY8PpoAhE52JBHO6jUT7sxxvukesqPlTu2N2e3emIXrqezxNN
8ESc+9/5fqNktS5XU0yuQnRlGCszu3ag3wwsxt6QFuW8GZzHeaVvMhgPGRRD2h699qRdNhc424wG
bGEcpJ3jA+Ar43yLZxjT6VQvAi4ccISTMcJfBy3tJkDNG7SZ5h/OczA/Ly654tSYC/09xyrEIOkV
YK4svnLkS+FnkzYMDyMsBLqrE55olPxIHPh6Lri5ApSzeuDauUCtEqU6bJk1YEn/rrrE9bqBSh+5
/0L2kVtSz81zCyTfcyC2P85FqDxT1M/81ieSeLzc5dMnha6TL2F0v+iwHcCYrnIL4jSQ22mdrvPT
uoAwwvlIKmZArFgSc+WY1OAn3VOfiIFPe1mO3tHA2h926mS1ljwhCr0sznez8BWJuHHLrSSnIk1k
ijvUdbWZmjGHTeaE2k/aUs9uE677FCv20+GMA8HM5CyIbHW6qLuCZ2uZoKY4D4IrjyvdEaj0I8ig
MO8fEjwHOXTuMg9tK+yEIm6hNK9sUZCL28xzCfx83wwYoQ3IZeZuvmz17Hikipc3T2Lc+xBHzI2p
r9a6uZIGol0yswvNi5ice0Tu34DBiu7V5UgQV+tMcn0KxZsESfi5slVKkYaKec9pScf185qL/etS
w+s7Vc4mChq4Otr+PH0nWD+R7ZKJ7D8xOWj80odSv4D3tgYe/XD5W5I26htEy+THUaSCqeF7vDDd
LBMjxZ/LDElXhoXhFgyKsaB83hLJTYXnYKOppFkfEEMWMIFo5Qovma4HYOufa+VNPB0Zn04V/lSb
DK85jWxHvgNkl7WrxfuPD5CsZKKY8v1btsCpytF9c5g6hxHWXV7XaPLWr1ZzD7NOOBELRNqkWM0U
7zxIKoOpHvAh+o8Yq5AWhIX+PL6GoEKFWVKEAoPV+HkL+Xlw+qkQz+6SqytaJIDilpr1qyhyMd/D
3h+k1jqr7ASVqCwsNgqVay87Dq1hwHvblhzI1nqIeYWZ/lXHJdmOQDymF6m9U9capn9HfVY3aUlT
0UofPQ1P/RLsrfye6MyeB1FTBYwl9NgiiraYjPNRVuq+0rXZo0hfaRL3FdAcys/RWmzeVgP6nJEO
Rju3XE+Wea2SsCwyTnO83MEwHZETOcFVxKkMy/cbOrN05uXXUxLAWHzfAcb3zh4RWgWNHSUsKoai
y+qEDQH4vq7LsOhGmuH6/raNtQ9MFzlzaX9pf9Cdj0FAju593KAHUOayfHw+oVDqSVq5/+ySIOhU
3e/t0ZLaFlykGzgGrMg9B2O5Ww05hXhXDLmluIJ7Mbj/VzT9vdnw/oaOQITRWNXYpeGTa83SASqK
yxzhOrXuE67zTYkIgAQhLv92bRmwLXaZWYEV+67xi+L1NRbNLAVTZqZLNJp3sfK1FgISIUBLyW1Q
HG/f2n5TS+TT2ZwPFES14Kskf4z+l8/PeWGlUsnLcaNd/bTLkuCK2zZZzRfZPS9M8UQhL1B4T1UG
5BNceAwnrG2Hbf9tNgod47Giqy6eHBpgi5x0lq73cBWEr0QjuZ/9bG/xQgKyXvFU6k99+zsTNhbD
rGTuQcvwVyDhy96rn12V+0TrOBP76cl1Y7ZhQD5uYMakrBCFqAYMD2UOEGOOV76lbYfu34nZfN/W
rCAmsPpZqNXfoDyHF95LLvL4f5658ICMDOf04Xj5aR49rXdOWPcNYVd3mbdvVNRRBkz2e70GTY1S
314fTRYUNooRN1EsXi9umg8hsv2kO84wT2yYW3Nc+WG+XXFPTreQi8mJKHVRbl9OD0lOuI+abdlp
h6qCigxijGWuaXK9wIoA0cf9n0K/gir19JxR4fLUqLERmgH3C2Qa5SOsXjV9VCmbk56GwJecgLw9
lJmldY3/qGXJ9gkt6ZomyxJ+So7lvH6NGKsqrSF1gG1szGvfXjm6fvs2Rw13r62kKDbDldF/rDeG
rUcRH7iXZK86lTrnfM1SVaUVvDgx1Y4W3ZcZZUmOSsNju6IWuvnfsnZriJMKkKf56fAnmLhS7oDA
Hndl5wRqq4K78lyIx44Nxg0syCBBTHp4IkVVzH576Hfn35FljqAwZ1U7N/Of23Mw0BKnyWXsdfOe
GdyT6SiAn3rBbp3Bu8wrz5mcGCw+aaECcCeF85rkYf3NiBWZmVs3nt0pmfci1aOE95YiO/qhwy5t
ZuN9dHw5wCijVbO+2/O8htm5nwryUnv518JWjSDiV23UhA3auap9u0fGbMySAxvAw5c0gaTSBcJq
5HY23xTJEwEC++ZNL5vNOB1ezd+wNBfjpzfbr0rnLB1qW09bLzi05G3wKPn7mzaXMF7Ehy5ReIs7
XHp7Vvtg9kTCugo7JQ/o8uRhOTv+IxiVYBze66yI1ybAVRiqjc9UuWILxlVeS8FruVThoXId1j4j
qMkd/rD+zjml5K1kVDkJs8ELzFKJRcUKX5dZwCPogVeoaVLezpvqHGWrvk2tg54OkDHz3gitXUBr
ICXxtgTQBvk+wQp8mNzr7woMOrEsOielhmIBaAMSQVGA+6szfizKljXjZdmWzEnFGkO2kXc5GDMV
c6sax4r+rpZQypfHxN4Vq+WIb0zO+OBOH64Dj3JYajYHhR4agrZK9LOfOdSILNgPAy5Fc6qb/RLX
/erU/gm6T7/gMxOsIlRTWnkAmFxvb3PzYqZ4KQ6seq4UKfycaGJ2HzTzC2ZBD49yAf8z8SALTniW
UwGVjfXuv0VLFE97gmDqHM2akNRri7fflYJWdUmPHK7KvytC+P+bnSKngnreak6xxwfEN2FHba4a
wlJehcGx0GIaMmzDfQsBC/L1kHmTi6q3V9CGSDvzZYdRkLIGutd+zdDrrDuu/Bx19VoDExragZhg
d8ZwLcMbu16suokrB3euuF0M2IteIbtsSJ1pB9QvdyGjPrJfzn9DIGCOu4SVOWB/XA5P4XI8mPGn
6SHioYb76+Dw3riFM8nqqyqu6CJso00OYgG74d46A3m1yWKLmrXgvkkhSJlwKJYxth6OS/oEht//
cfptSi4sxo9jBHTAVwSt/fogSl0Y8ew1Os7HiBTbajGWwvWZpNcUvC9qsF94XMKkPGl/jpTaDUaU
+SVnN8AYB165GXeGSC1QV/89eVYCDPOqitgFWz6BNDKCGl/yMkstoJkiVuoouMc3vuGLUHw3iRNa
o6QpEFkV/OrI1uHWP0nyVHrvQTU0l/DmuISzpWMciC2wdbgQMDFhyOUrYcReLTRgE8a0lUxPQ6sW
xxCRtI/OH3Kuj4qQqujDSls5hrZ8LzqcfIrjb5VGamo7ppzhuGKQt5H/zu2/2nNVSwt7hWLVnFA5
zg4EIGt0TrA8AK4EmeyKwOZee1JTFZLZ0R6nkQFw6BS7odVAZUKIdWxJvrWd0cJCrKCnr/Qag4oW
iS49g6xO9hldXKjqagkUu1VGIbzGQ1KsJvTm58Jg6fKsByKf3eg4C9Q4xN5RmjMkMtVbrtdG3IG0
Lp3Qa0ZhOrpzD8k8CzWpcgf+S6uJD3oerVh8z1cr9Dq3PhLsaNItFXZWgRC/W6St0l0+b5PWbsCf
ajQWL64/FS0REEBKuxRbVoHADnEP6g5/aMAZ9OV2LGh5WlV2NRftQ5JxLoYhgQmu7ZZOOdkskP3I
t2deN+Rp7K7kU53v0Qt6tfiwg6fzrW2h/gD3H9ZrQzm+FdcUnuujXgnWvNvxTgxpJCrgRR1/5BfI
KFAH/itemsaNXeOpbMHodOfcYdl8gq2MdsXTZM3NEFX3XIcH/EoFJcfL47ZXZH1ZMqCWP2hhhAXD
0zzfMDwEkaoysRvmXjovI1sPrjjaklDbf0gfDGeUWggJ0KPAp/YWa6ZPwhaaU76oodisIQ4EIBrg
8DnKXCSadtmema0Y+DaXYgUxCa9D2napMZjkpfMqgfY8skm5i7KY0tqBd6hrQyIYSAeTNabgcDmd
a5nbML7Lf0zpyvmlkDppO/Pfiwx9OiJJBRyJhmPetnvu+3hSJEfOLHZjW6GX5f8HsJmvL4ARNv5q
IhCTjs7fzn5DxQQMpax8K8SSuhU324INEzJ3hTSLkj9/jq62C5BJs6kh/0958bRN5v18+X7G8q5v
J6wfdnDpxplXGsYO/flSru02nJxZJgOEEfrANO9cRBuOuZDjQodjom2qaEXQ06Y4qSzkho9N6SnS
M5D1R071yqTyu5RvQptA0NgglRd3BOH/hn31Ufzga6JKgRFstJsN0gmETkqQLzT+f9LIvYllMGVe
5aMYy82NJ1CMenk/Og+Puzphw5tCNWd5HvFHiHSF7GKBl0/wJFuegyfQyWkFLRnBn79e0LrOt9cx
w14XMvdo5+mtCfOb4tjd1mhGlWwQqEEYT93GTidK6scHfg84urt6OqbGhxDk5LI0VhQTzWlfESS6
Z2YHuXS8yyCgJYnf+cu+Dg8w4dX6gBXnCUnKM/PaviemmvSWF/yIG4nVLSk7lQTRYPXSvjv3LjdQ
ALanSiBRypUt13GXKOle0HohKcUkL6pyYGMWOZYzE/r5NUYcfFIFePgCHDpkzQg+PcSYmIkbEi73
8E2ehVZQYYOXJlAeTS4LsL45Y6+bJtHpuOpnidwKN07QOpNAGLIxM5MJ2fl1jVEYIdyaX3dLoGIu
jhKOMWsAm3RoKLfy5pWsIIfxdenmIV5gIwBn+MrMGhn4gOZFkPvqoa8GRkOn9nwzFXb1kEfhmL5e
KdJvd3TR+NEr8cEmx5CFz6I17ENcsFXPDUTtAgqi61jOAjiGUq4fjzfeRwwsKn0cagBLl5Fg3X3M
7MkJttSf7Gx9M1afYmCmvikmZVABUiEjBy8gPlag/H6tPj/ma0+KhNHVNhsVSeWu7XD2StM7nPL9
WUYzbBsFfscEmM6SBqnLZ3jAmmWvaACDIbiirSoeku6bah9I4aD1WFeNwa1VO7oUQGSU52mjBvhU
5/5tGwby60hGmdxfuM66g1lk3X1FvTecsuQSx9kDvG+TzS9mkvZttWlylxnaNUraTyZaQ9GhVnZX
SfYXHhxiT+KckfgMVHSEiPvmaE6xXtINssqP2fSFTFgs6OtTRukJI/MOn2WVNKyF4cq+MYSPEw9l
orFuKt2FFlteEup3NQwrAZJ1/y4RWFBakUmeP+PyUuRm6egjRYR/y2TMezKLz+VugcmRyEVYvSjN
8tg6wWOxp+cOZVmjW5Ik7pnoMtWFocy3f8WslrthcTtoCXmiLlvoOhzrDPe+By/LnbRIUbFPikC7
N2HRAVu77lNMDzLsGIr1kFknQ1TKWgP5kWntGL7MKIygMUxbsyBW0WkLoNFgRofINVJH9a7rV4Ya
vCJW7cGIZmpRS+UyqtvX7ZI4GRjb0T2Yf7eL5ttrhLk+4MDF3KCdSkSESX6ElLlyBqF52tug+jSX
VTEuExqBO4/6rlFs45sLNUyAEGuc+QBSgllw0rPTdEJ82kQSCD89YE9ZWaTPhAysQ7x23jteGUVn
y0XmAX+mcNTWSAMjXLS6Nu4v0xRTsysn++uEpGnmOhNZAqDx0LDdBzFkTVuXPU0MF9EpFjeZpo5c
+Hne8XbxDiBw/e0iAr7EnofPq+j3l2lqUF4PyFOMFlgPIYxLvyb+QfrUZfOZLa3LrvOGAKmboQE1
+rLldfkK6FbbJK6CeCVzNjia7iX9AMnhyzOf8k3tjkdfqZ1y+SwWUmLftEzXepBb+DMdw8qtB7lK
zk8Di+Ha2uSbB0/7cWMr8RWu8i0waffIAZ+X5s6So9ktjPXinJj0Xmc+FGETLLJjYpxC05+9/bL1
FwWaa5yL/7apP4gj751CNZhumtCZPRZ6oHbaPiODhDC5BcwPqrinzGPEugPPPT3A8FIcHgxz1iKg
1iVTKf5oPSFshD35q8/Uwy1ZMJrglScN3An5wmEsCjtcnl6M+Y6ID4EcAKnPnjhnhxoeOyeeb2hB
pG1eBWuA7hLdOCGKEh/QLAVFBtDqK18x2SoN7w2rEOELFPu9vqayMfrktDolxTZ2lJguNlChMZoO
ZfQD8jdmfnRhyWTGQrvV+GESruCyTUQrMFAPkHl5g4zwhdgxKcKyv2IFhNd/xSYuWo+ShyLhF8a7
NE9/7kEJGix2kfKH1hQziqaGqn435Iyu0f4Gh3zCpvF0g57wHk9BnfmBLrdd/0HBKjIDKl1vJba2
x6a8NTXGPJjWZE5/3R+fJGuKvH9aSZ0bbKv59Jr7KoQMHc1Ub0myRyCqQMH0AjoZn9sfBHtzqInR
rA8e0ZE8hclUFd4LRAh+6akVd8ayljcZVQU/RirzAYaxWieVepBxxHYIgvHwzkpYpvlhS3zTznSU
anh0zs5oQMNrq066KPeYjLD+6BsXiuBOnGjD9DxUZsHFhl/VDXBBukpIIg4BWRr4AIz+HLallsWF
znq9XjuWi+OvXEL+Ups163QLNshV77r7m4bFfZtT8kFpEejlnezyEzQ4FAF7YzWORwVjIm+oLv5o
nWio0O0kUHRCTgHVe7CQla557EyTqIBDS8g8yeI1FjAdraRloY21k1f1v9zzjtjnGKiZ1t376bmb
u+OCILVkV669h/YxxYTFXooPCsxVG7O+Vc1v82HBIeVX/TrpmiTcof4DsvGtmPQENWY9vLm+zcUT
rAgDc6KHfI/KlCs7K0CWarpuM0RNvpPArTgjOczs/sU9QGrmRm6BTESbsBNXZO5G+4qvBsPaJecf
XFbwJvZvT1/4w7T/I/CBR0W4utu/Zh7NupymWDsydauY1PCgYmxJwBlqJUwA1ZYl63EpDf7jMdsF
tPS/+HVloPiD+RrLwS5y/+tL6cqSKwoqXY9f6UxeZEwKlbDgKjQxfbVjpIEaaA6IsyOf77hy2fUG
+FIuhqZYIDMiPA4eMJ8R+7imC+eY8edVrIUEbgiCqO/Z7h/wcZBYn/CCYCl4HCppK4yh1r+uHgqM
AuwShBpDWOcSFHYYb3bMObYx2NsiVVOexR0exjzqdUFD5KgjACllwkOAxy99IdN2ylM99BgD4lz1
yfrB4+LeRY+nOXoYwPoBYtvUAMTCEzaMYAJpnTQxWX6UKVCogJ16OtDQmLt7tl4zJsCO8qTLA9H7
clNwzjnugFVvsG4AEe4wqE7xxALrw+dzJCPgFiH1mFxvsPpV1GrX9qq6Fi19GeUURx/+KwNayS5+
JN1HH4VG8N0qODP4aB96nhcvznwACbizCkd82dFSMn1Zs+G6SHK/bShITqZYfnLnogoW5s4WocAl
lx33xY+pI5GsR8UJc7kFHK7HAY034TpK770acxlMKuksBQjTv6hSxJKJ++2AIqikX4jaVvS4rKwT
FKGZkGn4qqqzQ2cR6k/Ml1JyNbChG2r5u9U1YWbA7buc/+MDrNgXZv3K1PPIqUSg5KqHrlAEeM2M
dxGHEdcO7XffyELboRVY3RmyI0pYaZ+5iho/L+mYhVpr+LCdlg4jN6CeQc5OZbYBKgkcXYSRJBP/
GQ77MuFbhu3pAhTC5q/i1eARAswnVNKwJXVd3vHF/6tEC4c6Zj/+IACHa+aEv4NOWAXkd44Dxghb
aMkRXI8vvSMmkHP/D1DvVhbviSNEKvMbT0F01iMmmu51ht6rNT7fCqKpKN8OcOW6MdG9WTjuB8jp
CBGms8dRilqXFfd8Y0yRYFavK5hVbzeqyUmxAC0XqxZwbhG8+Yx6txlyikvRMw7uYBYBf1FPrefK
wS7Dzuvady5az1ktflLoZ4sZDmQoFOsjwDKGzmRnan+p8Bz8eXpwdh5Rs0JxZcff3wdxMHAC8+NY
JaGFfSlr8PX2ePs71ZWHvRqyJDzQkGKq/fHQOJp5KqZuGB8DdteQCcNnYqyYvBPIdIlNfv5sWFoE
D9G4PXrp+3CjwWiAPP+xwRonswzbBkLnaIhDTm8T37VBUG3Dwg6Lf+s4oAUp6vJkpCo2USBNq9tR
rAll/drol+LNmbULnrndM6WB3ACf9hPGKSm2SM6siMp58K3+yh2SwWBk5dks1otfSkfCRQItFKe5
yWjWHd1WceQocdxVqI9y0LsWVk55smvN038Ca80aQefZviyR8xiEH0VNa7EovMgROWF4yhIzxs97
eNvvlZsN7AIKyuncT5jF3Xy7jtKtKFhXR/0Q/OoVMSt4kcZzrKJ0B70bxQQ2D0RBJAWAoklXYzFu
1aBmX93h3UZXIB1pwl7vxRjmq81sCybEShwK051lnrBDSAnpfpH2vnaKlZ616BtMdNc+SQenqAxd
cYhJDrSoDZBSUAzwv9x0kEMVoM+8OpuC6hIb7W7lDZBKlpBMK6uqrEC6Dj1JygE2rh2q90veInle
0Po3amZY4z3w7MQhY7JLCk4LMXH4ZHnRJ6ob0fnQRhfW2vAtkWeilft+HFFVFyTCc/Tr1KWw+Q1F
sQmPnMdbl0QQiEgjfSxaFtkQf6ghdxg8mos0dq/4AdKuLRTH8+yWA3eLQ2+mEF6u0ocDcZbBcX6F
1iESFOwcF3Me6tJj2tnYwFwWrDDbtLuXa2rSqCKQnimCx4bGp9yvq9HPhINofDSGbe8R2dX24GiG
i5IQ9KanpQy7utnrtlFgjc49/COTGEmtl4EkhcciEUleD1hGaMzoN9Otqdsbq9mCEh7ElLeoIMFE
hC0dtnpckWiUG+XLt03wE5nTuO1qzMpuQoVHR63AEKfbnYDLwdcK/hCVpaklE4TWjGD+ChIDJSLQ
JWH3JmlkdW9Yq7GSTnWRY5Dx1quhoWlwh0o/PZeHxI8OFE0aH3qDbXrV9ZMEIfFN+cBuIDf5WUY4
qUXDk/33apAtTdj0+Jl2xSuthmLbgHsIRzPmgoxeFKLgYjDB8WUE9IKsWLCsR9QzEjVWxn4cQwMk
YWQWwvKq/SR21zGC2n0Iyw562ODO9tg9Kw5MDP2iJ98U1197vVkoWPUWqXYym0XmmzmKl6qMKmti
aUtjA8GqxRh/4Oe1bPZrWmOdzhF6Cuhj77UFLX5UtFY9SqGH5Vbh1Oh05kwDMN29rCVPw9UhNfh9
/cPLQlPcoQfrIX8ghlidCAa0CZ78gBnQPKruuFTvhnUugh2tcUG9cyJ0mLZambjgJsclxZG54E/J
m9qVFR5RzYacEUnyNyDzUUY138hb97Yx+N/7KGp6cZHHwl9lQA4Doxyka5Wamjrd3dsM49SBLLUS
/PXxqNCrTskrJsklxMSqhGpGkeMyZPuS7PlI6rgoARGNHhe0HVs+0wwIhrKCC2DQoUMeUDbA4uXN
kojb0SAvf9r/D+2R+TqFRjirrWqhVD0y7oLXcz8uBGcmuy7SW1tagqnmoMPQVmiQu5pmk2bbQpB6
YVLJ70aobqVue6mmn3+P602n01hL5MbaF6RyNQ8YwSBhFV5bYg0+K1Cb5TUpnZxaoMwtIZNTT/cl
8cM695fLoyzVO9cIHdbvajc2Gfb2aUBafzz0jdKgl5aemsz1Pxj//gfZUEimtjevINr/s3fT7tPG
uen9TRA9WxpQuIggy9bAOpw4ZcD11Ji+bIo/RgoayvoTMHohhjxDciGX5Hh8aFf9cfX/FfFWm23f
imqDMcgzpgoj+oQunimWxxZ/Vh8FGpDsuKt77BxLcgOAuG0Tp3VQu5A5F5RpJuOx95rrThdTUuOs
pRlCgs3BR9gntwK/cKC939rNZqmwMgzDXU784jYM76/IT5G0nktMEmSX8D28ytam5xxdEIOZBYvv
nGgbyHnHdoQheowQ++o41QH2w4CgKNONzy7OfcAvNYiKuxGtRG/IYHTGL7ksN6TtUtnLW+52TKAJ
5jYV5KWqm/m0LKXqsQxFC2YRwmpJcdvtVuunD2qoY8+9baKMkiVTyZeoTPwWMlztzNQgwU3lO0av
Ksm9f43lq/XZd8WTb2VELg/bG4XdWNwMB6m3vXricmbHxil+qCejTe3dwz+tfx9HapRJN8wVtzB0
ikL5ZL8lQPgub+jL66GI6/XeGwAXy/AolLBZSamApQnexLdo2rv4kQ+iCm0fqyWepl6ZrsSsor9O
jXSFvhUUyKPyrYM5TLCtBEUTzLvYvFWJM2JVH/USmH+fNAH33zx+f9y6/I50NbhQD3iGiWrJftML
4YREh3zOOT1Nb45InknHwPHbrO+bz3db3kLCzstNERt9QGmUK8RSq8NFe6DpMm1xL49mwogoqZz2
BaEUCjiHlodig+aBf230Fop8EsoxLv+bu7NoATSNzTdxOOq2SKRd3Cw8kj9f2PWkyjigRjzOuNJp
Vj+LvJhxD8Djnpl49euQpltMFl16x6PxzF3ID+jgMYVwYmOmj8wi5FhfMl+okTuPO4n1WiY2lb3e
SmgpDkq430vAGzGVY2AfjEyYo+2uE/q7q91Rs7GR+bxi+4ZpOJb5EmWzyiucFsj0p9IlLZd1MTcI
Hsv+3JeuQenrLx8l8Y9KDGPVdv/c3T6EsDCbzJn4qnOXDPBezzDOZJ1LjifomelvqfqD/u8EsBwV
90OSDestnAJuYgNe//5Sj26WrXw/lwWcWJrG5Bmr8L7dgKB2PxAGJnc0SgI0bOpmMp0pDJT+w0v+
9+uGNCIxg7kdfCFtCFlzITdWr6GYADDJvOf+rCEmwPX8KI6qCCTheLeyU6JJDTG4dB+0MI6AvhH6
Kjo51iDLfPuhJiB7dhWX+dxdqPJysfB4vNeToR3METpXqHvdXUuIQvwkdELZSCb08Xt5OvJXF3CN
fpjbabPpRiLVPcsUV93Pf/mvRkp+6hVSZHncr9YW7jsepqOdKds/7qb09gOyUNJjPyAoNFmI1Mcb
i4qsjb2W/gt6ngF6CNjt+tNSLgVBF8h28yQDyKw9qqmcwwxK4rdKyImxSNV0VIeqqoGhvnc9BmsR
BeQbwSaOLcDMpSvQ5Ur+Fp8IlqCJFTCGQfz1CPjfIzOvONLtGS3FSUPl4AsfbR33Yz1+sIK7JaaS
bfKRdHcjqcIBVj9dab2nD7tN5rJPZ0/QVvbl0PmfvI9bG9t9zDJCoV0T7oDaknHboZ9Ew12e5iHW
LRwF5Oybq8ykp8Z96iVyb3jcysMsfKsta7rcddDg7lt7M9807M4DWzxpEtd0lSJRueywRtJLlM0v
gf3U/fcLmIqR6jk5f3Q2fRtv11m+zZHgCS29Axk/vRDct4n1q4LoSxHZlcRSRbQQefdfnEURyuH2
VKXWRB56vUujds3buu/Myb7ztMevGx5+UurKv7+Ng59sRZibib1XNzQGj8yyljbm6BCmcPWRLJTC
v7UxHe/6Hb26RD9L33rBAdO0UvSc49iSraY5bM6mULwRp+qdJzDpdx75htFBJ0NVkXehqR9heT75
3y+UFpOZEhPmnIUhpw0wNo5h7/sWzYwGE5+impNa6C3UdD9EuMGpngzCxDYrLnyszegccwX6HI94
bL/pW7WJQ/cIKjzQ2tHq8hrp6X+f6riKD3l1mwX0v65VpaZ4CAfDwKJLZD5oeLkldFsFq8Tl7X4a
HULwYBzcxSoOzn2R+m0nRl7XOCyOqIereRRXq2ZnIU9x55cFTTIUMJErGH3B0u+QiO1TnHr4pHP0
KGDaVz9hNOveu4bSQlzqbr6BpLETXkj7vVTO7GslSuW2iomRnNAttyLUYs3bSuKN9vhMXNNwWdt4
+uoWexHVjywkAs/ygz1+SdVgEANlHU43UV6j3uK3VOswgv0c3+xRD3Hs6qAlDkZiUT2uVXBB4Zpj
c5ZeDhSZIUolrlmMn5BkM0atflyM1qahM1NuAIgmQmrRqSTdTF32xYVHNoHdl1JR6k9y0VfX3b9j
O1379c3omA5f+jrwTudztzTPbt/kQ0VydUKkpo/kseEQtIZdTVAPWPFdgWixtIoCZGs6veW2VaCH
4X1t6+xVoZECE6pcTkDJxl6AuaWj9QJxoIwf/eJh8Ewd4wk5kk+QsrpWD7Twhiv6q5Jo4gQADcDi
G5ExxAO0stV24GRvstjYPt7mBV8qLIo2aDpX8Q0mYKzLaq1WH8BbabjwfZZlcNd3S6SStV6mZhuH
/c9noaV0sKDP416Y4lx9U1ou7F5aYzJJcc2fXQmiXH6zXznmgSlontcf6/sQAmrahqmtXgmH5JLe
wf3lS4ruMA6WpQFCHK3g/oEjuZwEC5tKzZ8T4OyfM/mwF5MUDaVLlYkgjzBIpQvCQHSht5hCx+vS
bKdRgw51KTeXaOrVBYSCab08OcSPHS2bNu5nxlUiqC9HqkBvP5LHUCm01qU6WXx+pd+cm75356fI
CUYNAvQ7/5JyrIH8bMnGSB5scNJdZMpfHayQCdc+v8m6J0bnujOmWlWwAkUYOaf2MA3MjcWon1aH
zSIJP16dYoCJUa6cZL5CZ9zKN84qSmaQmhuCqVVaSXvlS7ebKzwExldGcC42kzmtlDTmCTJX5e7z
cYkQhrZDIYiKulTyndyas0niddcSIH3X2PDNcpV0EEsOavCEDfu76Upc7RCheePamEdgWu91Or+R
PfgycnLQJXoomu7IUYSaPhV2HjvXZG2+GyISE+DaY5J8buxwrxD2o12j6FE20OFv45NKtbbNR/oD
R1yfqC+9HQt2OaF4DyvgK5kKORMZ7PygGW1ACVSAe8nwdQnfAr5/TIWtJyMQSp8hOwy1H5EsqHIk
156t0yQjEZzNbX38dYyD9d0qAH7pgcJS+TsICSKEAoz/M6jTxAxIt4e0IJcGsUajGND3DJ+ilSZ1
rDu8qw+EdJ9MuqXGnM5qtovpjPXXaWkm1jTxZV+imIxMmliGyzjlaBjviSn1vPlwxig+dUwHa0Rz
r9USg1R7q1S0edn4y2KeDSgv34/kUx4Qc1+Ir5Veuu6JqPLLoxy/B9s30Jv5c50+eRhgSKyMTxjp
KTMYGD6Gbk3DKn8F4cXPv2thq+XIp0bVBvZhP08wCAO+4kWBotC61eVcm4BRaypUwF2MVLKLtsj1
k7dQQk8ob5z/b3jfcRyVCIU9oaXaUOY+kcfEHeqrKmzm+UwTowAdQuvhPr/5x7kMYg2y3l48e5Js
kyj9axipvycSfBP3o6QryeR8dVhuHmrYBoVRiOoDQJ7+7yHlUWcmgWH7SrdABhuitWqIgaFVELGh
kim912zzS71tiVQ7XwaorInL1U7m23kU2GvuyuAoHOGCyOcGDOqwTCI46FSzMA2SVcOGGIvYmLYw
c8Mvi+U1UZdiodtoNleYaqWQcYzJn9uJR3POp2oG2qvglYFWI6YmiCIY5fULItbChEfO1FaZq07f
TKrXvQaCFLPIlVCEwdahmb8V5qlL/gl8jvKwxn9I6xEGD7GhNm4udwK83P6ARhD4avPVVX+M3eaH
s/Gw3JbJfmawkTUZr/KMEoGSYls2WrBIPfV5syptVAyGkhNix+QlNk99IX2wc7nB9gRRJdG5YDvU
Zpv8lCOq1q/BCiNbpb2TsW9QpbgzqSOXK4YqYbxUCdFh6q7IwTUwCigwGRCGzHAQrWzyNY10s9AQ
p/+TLgk6EDHWGVO9Gh7Ig5Spkchd3Nkpe+UGy/T8oMu+XSnf0Rts4oORDHHjVTWEj0UcM6tNaJwK
MAScghVw1tISFJtyX2Ds16kjIMxhUGxCDZmH9fZEU4iaMZ9mADHMSdlbUtki/qM29b0AhJ+/0CIh
0XkJEd2blKC/7fY6Rn2T3eNx9ixRcZBPUeLBlVLJcXpR15Dn7ybVYr7cMwtYhQith8dOzkH94xgd
Y5ZrUrS4ePundVnigBAhZeOsrrKQUz2JqjAxgZgLGo34KlNG+PpEDA0jYc9kI4JvG0Kh6voV2kuf
MpzH1CoqmyvwzZeIcvH8flXpAuoc823MPIPwxEcFY8p/rvjOONMPN459jCP7NZMfeY1BgcIHBz3e
VjquRr6ba0EOwsDzt+WCp+heVw9xSdjSfOS/PIv/wvsmt0+hL2pJYMkHgC41ZDQ2ezt2Ce7XVtuH
nVCQKmKzk88+rCo+jhgJ6/+pe27VFsRiIrU+DP7eSnJYoB8VktIzF/jaPBuuqOl4yI/6bs5ms+T0
hubKYRzoxAYf2bZTuVpOLrxuL8GTAR+4OnA7WLYrdab5630J3yP6k1d87ISfmY415e8/pCvoogYI
E6MIEazw7i5gMBKfVSe3NtnnfXHgADAi1iR0kMM6Re+6cbpPzGUdeTUQPwvuhuQGp5N+W4PtjzL6
rISV2u1jP2j+OACMrNmsJi/D3UfWCZhtU1RS5etDZjrZLe5TZhaU0KEg+EXfSGLFa4y1WvIJUH5c
tfcnw0RQj5ATbPJ+/hQU+ha8BnVGnKLQAYiYrN+Uev2ExhfTtrkI0yJDdp0P0ySHqZk5zOm/aVNd
4qCC56QTLZjZ0sfqGsSRv5LpOv5qt1Z5YnWn36EMzhqXHuN0BWzkMUwsuTc2Ec/0iFykNJST+mrs
suOcR5jw9xEIYpXeVkxRKEpbX9785/lOE47aUSD7qs79vMARGyl3ZiGbEqIm0ggTFQtxWzBtTAjP
3QPLDzcoEgCfxLgNJ5whrWfqn/iG8/Xoq9gaBquJWg6/MdDr3IIkwOGnG0JR+H5p2zkX6a+XMsJX
eRuGC1g7txywhxZEA48j8agVA3wHKH8M2tV8pMCKTWJoWASv2T52PH+c/7CVQKexm1CU8lUTlWnM
irZjH/EfNbStyVJSCNVnP8wu8H4Up2igKm8NTQJ8yHESwLU1mC795/kFcHUDtJC4hJN39t2M3pbQ
ML+vBYvvGwMIjr52ViBilmuGLnqeI+2bzDNctP9Hms7gdDo8Bmj/56bEDWBde1aKS3838y+3yEdI
mrbUB+N65HLxRtvNC36TbtncAK4oSF6+CqtaoZdUZ10moat61/Mr682GPWP8mfWMVrkRYrPecuL9
7QWH4HiCXemXHA4BR1aRe/r2VNWddano7fhzJJfQbYsUkGQ1PM/8ALpG0nbvW+I11ojuqftGUhvZ
lYl4D21J/7W84jWjoZLsQv8EAkn77z09fM82aiL/B8lOadpoO0MawykCrsY6FLWUmLSXx+X3l+rT
QkGaepkEkDz0jOzbf3fY+BQQOM1v2ODv70b0y+2RYCqSFsa14e6fiOiPP2UVLTs2V4PD4BhgOsq5
J4qqpb/hpbrfS4eVIP+MntLWcOu5zEL+kRvV+iv4zRovt8/D/lyGJCxdjOwHBYj+8JQ7c9UtW+cZ
09O3IfRIeUb2RjXSHd7wAdXq4wa1B2L4RwcFKha5Mj+pFvTO/tBhVoC6xBEwUenFSWk2vjKcqoE6
88eCjyBUr22X6qBeQMlND0jTDLasO7+rXOczzo9R5tgeppFn58AmI+JLsUaxAfVfiiCvVgRRbj2k
zMV2qlBTU2ZtVnm97pEiRgoFAeeXeQtK2sqLrNVTTsZ6rPW6h3/PGPwu6DY0Iyc7Ho6BKpYRNKpL
wgqCK/say8CYBmp7b6oWpy57PWzuQfwmhXJa0FqU0Nh7j+fSahf+cm0vgVgBAwi5vyFrfcZAd42T
CvLkNp+OOvkFlhlxaJk4yNdz94xpYdGjOrZ2Ki7cVzgkw8DbZwRfNuH2O/1NTB3PvPGz+yx/aWWR
pOrAU4kNsxnRnqOiX6fiLWAcfJBUrniKJyBiRhqwT6szkypWbKdo2kWRfEm8hUBaXdQkVS/tzlkc
1/C4b+F686glyfciykUE0fDuKaTRxBexU5HIQyZoACRYnzatdisHISplynKGIiRw4VvunHo8s6ik
taaZNtWY231o8rxR9BKEgcgj6y9sm3e/+TQ0SfxgmQwTmC1DS64qSrmZLyTZU1fXGk/z/iDwl59c
IRoMX6DjMvHW3CbrAYWkQqrF2whByVC9FsXmcYOPj7R5j9rvb5jcOtqyxDKuo3iH5+OEPLP7Wil8
2vzCSiKMhhV8AgHNiJ4YbLcqF1mvdV/hBjYsB8tfng3p/h+XqHc53yFvyd6K7UfP0UACngYDPuif
UI7edU0FNBxPbmlmZfRWL0ljbAW2L5ZQsW+Y5eZg32KOHhqIGt2s22ZoScz3mQ/j2D1drkCzKA/4
q9YlOVsGYrU3DzPsdQqK6YVMSNXUdUcRiPIPdCUHGRZtVBJybDVS0e2Gr6mES5VCAhuv5/XDg2qA
lOpVzt5uuSmIo85qhw7h/2y2AJtwsfodeHhNVyAnpnVsyxCnXBWL1+XGLkcZIxGq9rgvMEcspFj5
8ZuJpHVYf0nLFFjXuVcveXV/ccXIez1LLfpHjrlTGY/GxyhuJvNFdWXoFPPwhoHuUj8z6qGnVFUp
pH8qaq/zRikRYkn1Dgwq5wfXL/sFo6o2TUM64VZNRy3ePXhac+he9sLaddLtXEC3jJh72HvSCO9+
+sCj5LOOYwGksE5876t+4dVplxInbnaAVMIcaN87b4gp8oI4SaYXn+6uFQyv+N3BjZKG7XqeYY0U
J/URdJVySaG5KocjLPxIbwK7sThwHaHtA3pYQh9j2GFOIMGOzPf3CvqViJMB5wVp9eCb5EfTsW0U
qvy59sEyhOoJs4V1ltjAyj31Jn+FXYIa0NHQ69Ib/8uYaMZqAI7TSuPUA3YX2VJpzsEKE+iFiFKW
BnXTkeQvbe6/Wf911DwZbo7xr/9a3j5Xy88+61nv2g/BuuseIAbe0M/8UbjPDRHKnXZ2CiAbiL7s
xT7gR3250qtnZMYk8m7klt8Wvdae2v5YPq1JPh1QQgeKm+43BQox0QBbcExN+BhoWfII4FbtIsJs
4kDkPoE3xbHjDpDD4Syv7gjskNekpRTkXZ/BnSqIQXL554/Px67M1XvXiZF5rIhRXWnKTUlf9zzJ
CCtSDwureZtFrlY5VIPvebkH/xDLR0z6/QzfWN0nVhCifhrUOkmYcCI/1+JKY1yA8+E7sNlDLfHA
YWIuuHncgLRbadclPolok8zqWa344lGR1SocjfKxkpl1dAYdUghMFPAFBDw/JBatJghJwsaOCy7H
0X5iU2BeL6z00MMAvhC+UH2FsQWzIJ7738gKSphaZbYnCTTlwbBVwPY2R7V1ZCizTnBxukwfreR4
/EMdI1LrNl6DfPAVPA8A29FowftTwSvgZcegdL0+GIQf7U6UsgrA2BmjX8EYdKPnEx1E4r98njeN
x9j8vNmAB17VLFmaP4jghDBGg6MuAAVPAwhoevarcQu1s5pBzV9mXXq+JgX+Q7KNMApDUWJ7FXxo
az30nI8PVzCoFkWl3aobexqlfXaTxRHEPdNIfqk06WgDsvJiAcqCniisGXTVRGvIVAbRJ3Ck8rNV
1np1xAVvDFT4fcn+uLtxsFYpJr77xfA4RIbCOAz5mDfwHFBsem/1cQf9aBr+3yxiTfLmgty98Qtm
H74r6r3hQMorKLXx+eGK8rwyheUSbd6mqpq2HFJsISiqye/VsKvhJ3rDLhftv3/a0jQihRgpue46
7jnSQrdErIXaYNGjykrMQSrPz96YYa82I9+dbvbV3gMPj7L3cJ9C5FowWlUsLG8WeUQvY50MO+Dx
GaNHZb5++nHq+ItButCtDZBYZ8KW1f3P9fcDO4iImhEFIvz8QuiLCYADYW9BGKOqBgUJ1keiQerm
fsxkRL1sUGseudD3L3mVTDLtAV23Z8TiP0Kdq8QFuoSobBtQrKtkjCSxmBhrxmt1mMFRm+a+PzyK
wTC/f1Wc7W6tj8Me1S5276rLf9WWI+yRLOyY/La5KWbr1mD6ND1DigEznB6zHPxqgcIYlHv0mvOg
+IdJAADvqOMOgsLDOyNbuJGX5ThDEqmIZT8MDFre/V5+CjViRvl3rarhkCSc/ThgfTW/Bac5Satt
aD1Xd4hMk+gCAGiAop5vaCTMBS4IySO9Y59AZaglqYL1F5tg4KM3ss/BvHHj5YXfE2AJvbEbUATu
t4mtxFLgF89gAGBO/220S+RboKMibSWe6QiUUBRVw/CrKz9vXBjFxybpDm9r25NDQDUAMQ7YVB6j
sZpXAmj6oANQcwtxDXj3CIADPbTvzWV9N2cEqlmvnvJ9cGyA+uj1u2dYQO5gM0vXiAIBw2S/oQnT
3Z10RncVkOdgFiVzQxPA482D1m8wM6rM0yiUFNIIhLiIiSg2pp9zqFcum8i1lynRMrtSfny860XH
QY40mpsi8+byOV9bmmNpU31sicQQCUiYyvBa/Z1O0h7FEYyTD5YaSh2duDELBoyNE5ohBz3YBc2z
fu8aFMhc62GZY+DO34xO/jNbTZNqq6IyHf/Z+ae/MO6F8o3P5ozcfZA2qodnuZY4AyyYJUPQAFaw
OD2b4OEdjreQzcaC3/X3Lbk5DuYR9aeLDn357ADMFrY/LwQgS8ExXwAL3ZpfD04GxN+f+IE2uoRL
RWrkTg8DzGn01JxhKrafTTAR+/EpRkY+eOSm6DlwTwODmcnnSsPV7PdeVx9cJTartmVYNbjLjAE8
f3A3TF99vzOC6yvhgOHAlxMHwmOedDuomHZ/roOGd/1fU878iQIeiNY0flGMiq0dumzXQ4Re3EfO
YCcdH/So3orXmnX2uYYAyCv4AVPrk0NG3wfhum+eGdimhDN78Qf+bonTJqNSccpo48bKe7b9IBgm
zdOTJQRtgPW4iJhigpq7IVuldqdYw0HCLIXYUpTDZ8dPrX2nJ+XYy8scxyPJYO6xf3zssA9s9dQq
rKmr29BObOxtP+EWOjgel4nxLpkd2UY0tAYiCvQDYWYTnT+l38GkR2aDScUUS9V8pVvctwdjMqlg
L8Vij1SoKmHHaPZ6HkDkdMyeZDcj6fFXF2TlxFtBlyCqnY195v0UgX/n4hrDx5X+MaY1KPd8KATX
TeYzooMF0IYIz1cg0fyD3ONSOtQoXBzMlA5BWbzqdNbHI2ZYZuNEdlXj3rGOjFVjWlN1OfvC8wxR
rSDpGcj7Z9ecivmIskICQWbPr/eKQqCbJ9d+L3TkNXjlzho8vVaTQ3O3INxBKHUoZic16p3fkDrC
zyvBPhj/XX4Nq6NbT+ji5wNBuqO3YwaIq2wdAztssli1xFV2W/CIsnc7PGgryOQlO1tg1c03ycwu
Sx9TKY6UpBp0+1Mu91Gvdje0+yzQ+mZ1ec2w+TrkXjqvz5WShl9oYsZlIN9IPAYUvAnSMMJpfXJo
+SdOiRynC7Gnb5864MihZfJX+eqIL5GeOe18yw+v7uXWJKTqryAkumedY1MnXA7PLGVRVm6AbV6K
jlGWVUNu0m0+dLHFdzNDkINod5Bb5zL9CUFkM5Aved9SzWO8PAb9neST5Awmh2sNpKoN+y2EDqVh
ZTLPePPBqCqzg+N9cCQwCq4Wbq5WG5UXwzXV+2t4h+XLXqTEXDIKQDmvS7NhLkDEyEuGJtBYkYA3
WMYecQ5Z52RpDo/oP88pJQVVhF/LXuerSQIhfErQWqPgby6uzR7tULtHzB5J1n4x8fIdKkF0sgIf
9Cq6SiaRDYH+K+pE0h++KL5DjgPynTyNU7RmX9yZbKD312fa2d3fiOl372IUeShOYxAB54RGY8rU
4BBopLaZqJJPuO4LO5OVdScp0Bwdp8f0PKIoAq3AICB0yXVlF2JPBQO+gaz7DM140JjchAex1P1d
XN4u0HlSypXVen58+xkqtNyTc8t1K0FX1ftaoyecmOHfILG/s13bZblVhXP1eahx3MY193d4pLxU
xS6FBuXSalGteNIIiUigpkQW7e2UMU+SlUU9D55XBV4NB1QEA2A0aIuJh5CF9u8fbVcxneJCjVbR
W8Ky052p+VJcpznz6qbKms4pKISSazyAaYi0nMVOTtqfeMGoLz9IQqxSN0ULPb3bcML0dxpK0si3
6NCq0sKwOSTTNqAaIpVWNdN5TaFT+M5XTA7QEIcXmJJMC+vVaPz+HBIfA/CANFoQO2XtE3Dml1DR
y0EnEuBV6oBDqFNIsNNiK5YmLLNq/zz0pZVYc5DU0KxdRGT/SR/ULvnUP777D1mZCFv5okVl+CR/
gYys/d/d8RRkjXxbIqdqa0zzK/em8Q3t9l7GJNzq2piG0+0DOVZJqbN3KFpPdxl5G+rLX3mD2bkt
YSnvrp++WIR+W2nZ9B4/fg9tbK8HhKEWu1cqbJZ1kZcLLsMWUlLLCtjAyV9RniiQArHdylEOK7Pk
ODGRUI7khKdwkH3ewCYOdckeSxB/Cwj68XDomqvjrOi0QJtI4Sosucj3wSAc3N9Ora9CXs9HCvDB
0iSUr6ZvAp0duJWzw7mmTAkZsZXNlTWzCQzWxIjnB1jPp+RmOy7IhXNhw/Q/qZ0fLWxQKzhyHue5
sLc8+sTbhe36gYdAlDzqoZIXSDSy0YP10tCfIuMYmfnO9KvcNXNDb+l2UvzX2AvYlZaePJmJhHx+
16olVscJnspz3yxu2zQrHQSO2SEEBwCajq2FWU+VBT4RdNIO6bhlZp9kU/PSEfjl/FJs6NBoZsou
AG9vj+Jd0MZjFqf75hdNX5cyNy2TZdfIo+4sdOEChLrglaZirQZnoEdzmyf4A8dDsZEIKit9piGZ
IJfsbfX7ZkLTL0ZeY/vqJ6MiF5edBLWyaLpb9ntwQaY4R1p6h1C9EbgxX9Ls2DlctfM0wXfg+wF4
oqN1vCRmQZ1LXid+RNv0cnjnY70+z6kR4ITJY1/AakVq6nqMR5cyVzLT1tiH+HicABCSCnhLXQiK
aXtjuG558e4twC2YYkDrEny4pTPhkBjfBAKe/j8g1WP+sNM/fYeDg8SMBjdF5Xxnacat4turW7fE
F/3SwI2kzrdV9xEZ9/iSnBTCzis7J4qAFYFerowDOVvboG4BAI/CKOp8oMkeq1mjp/p3STHKU+GZ
tIJW+iXoCmcr2AlI7rs7rmDMT+MFHjQ9B4k7fJZ6yzYiwG6t6Pb0xudai3TR1GVRDRS/gY/9Cwod
G/HKW9qjnUAJUmNZ3Z1B0hpdKSsvzTuMSWXrHApIEevOCA46ocZcm3uWd3FheTA+xMXScBL9EtmC
rJ5q5LJlbfdLcHJYFntnCO9pyCl99MP19eAoPj7NI0TyCPTftBUBUKQcQfOoglMb8jZ2zpBf/w4F
NFdZnWeMw3DFDB3DPA5QrMtLkKoBd+WnUkOiIMgRyatakpesjnDfNZ0+cHcBggWCgmCdkCZUu96u
s8MBdvJOf7W3HXc4FMzh0eDxs2mkNCCqgEhQ3TzPxlwhAjumDrC8Pvh3/+Jca7rx/8baaRiomHwh
4ls1PQAMOWyFH9cQH73RH25fjStWHC05hsLcakWvqKdLafzXggyMAUbIrujMAvTi3mVQ46TY14po
4VGOWgfa9JQBFOa7w6uimSgb4TTKbq85br1BqLrmsXtSAlZTPfrBgHkWR1AHjyw0V5Qf73llp3Ne
UYpEZdAsDp1aZtWgMMMBPy2PXuER4dWI5+SPBtYbxt8ST7dU1L2CowWlZZAfTZK2QWJwHxG1lazu
IkyNJzZE22NIWIM5M0pO7crqlaF2zVtypNAmkaQXSKSQNzaga0pcmRPVroUAyDXqV8jw20TAFwws
AWkL0eTMdescJ6/3GxkmHR8rukjjwT5ho1l93mvXqsG8am6zomPvbHB44X+nmvWyRx3kj4eHPao5
kJNBA0cxNEPKjag9teL2hFLsfAeDtqGbYjbZspRj/d8st/gqBeloK6simKfDZIPP9k1vD7oScJIa
MvQKn851IbK793Wuhclbf5GEdNibHU6YSzIhDcUH0bSABTkT1eyW+TZso/bP+y1dPh+SAAHrPn6U
ftWTFAqegIyIe4mM6OjT9X79bJPJczMOgkIMHiqNAlrhn+K9vevA4a5+12U0QAr/YOGr8XmrpXJV
qVcwIMqKqeIKBbAjR2gaNXNc8XDZqOYCujA84HpwdPpY81oBBjn3vrR6+fqa2JPIXfNEPlUN/l2m
tPdsZ4r3AJ9aGwbnWthPNS0VPZ2pfbKRoct0OE7UR13Otad7/Qq8f5GBizQeEbUi2dFNaihXAmVq
eUcPJROYuPrDQvuO+j1ciamwWIl6w8rXDxfJzqOqr6E5UMCMTu69CQztQbBpE4MulqAc/eEka1Mf
8I9+oPdHGyCqGc/+dpx58YL+1CLYvOC9k5pUgAKQDcpQDySZnnGTKtvlOamdSrzM6eW9UcjGE2XQ
fxs33OcoNsjHRg0rrL3tjBjdofkA69zhJl6IRH0kMcK+lK+Pf9jqvaotvMBdwImTSM6MJGtwrthL
w7VE7fs4+JX3201YhDC0WA49UJRHXknJg6aZ8Aim3SsyCKRwVLgf469MZpXZHfpQFxnalztj4DvU
IeJzWjkOFFUZldYdeJa/Wm4Gsdo+825gUgNSAJiZwbJergVoR/VXyAZ5vxhdo835kipE8IqqIMQs
SraJuZ1HUMdEpMVk+nDObwF+/RFUkf5GXpDz75jy9Yo8iv8YX4NS1IabvHERAKSkOY8vT0jwWpA7
HaK/r6Q7TnAp1pIHU+Jeqqo9Ce+lp8WzzBxDUdx8XciiTCWJUXYb867gOW347FUOGb1Jd6B+CKsy
Ds9r5OOuQvV0fmu/eEN44+SUVK1XlWtUkpOFqBVCXHsHLREuucsb/3JknHCUqqje8JAcyOIPNENx
DP6qXPuux4JHTfZkhqoDhg7p7OT8fS49/PxtLdyJ7fBFd290iud3NPs/n6Q61apLaeFAHNdYNleY
FhTf5KHYAgXMN9RM2uu7c/VFJinYQGXJCJrudKVM1n1SAumqRogGFZUjFrt3X4Y2XRU1IWiZa0V4
jq6oRGzB147Ey8pPOTJNJhmXHipy3Wl1h+cdj03vZtxMtBVE67ZIAns9RsfdQ4xCX9rn6RzB2IDc
yqXN3UXMEHL4xHb9fIklhTdxB+3J+LRVoWiaDqPGpT5mT36ibw01uE6HiyQrbl+ommcnUDhXrRLY
btp0rjKiANh/X5KB/J7TmTDszF4CjR5gopM1umyFqo/xinqsPdUgqinJ/PNhEFvkM46kmy4LeGcU
N+VhBwH6M2T+zP/HBNiEEiy2xL6wiq912nykMm28hcRSwtS63lYyCXjOPnhesC0h1MWUiSa0dEzF
OPuakVQnePHhvP0E7tptEOmv77mmdu6L9123RnwRlGP7A6HbZnsZy5OnhSw2OKiYzl4Ub7eN/6ch
DKwGuBSZXSmYuWEJ0VCaEXy6e2Gkr9Juv48c3KUhI3LDJgD+ivUyMTt9Q6zn6S/khpsuVtMH5tvL
SiqV1pZBYVz2eV6e/u9ZCJ1k/LUMwZS0y4gB9CdQ3Jmo4OzOaGzTVu64ZRp406U+zX1U1bb/J6op
ZzlhGbBUR65usqOdjPqTCJLpxZonHGAt0MHmCJTm5sFnBSQcP60RvvRC9DzfVa1pYe+ksouviJ2I
y3SfI+Pht6X0aLJWillf4pjm+lD4w9yZ9ZeddeDmphyYETzSEWV8vchHzXRhZSBYjb2wBh8D+0Zu
qKJeCnWQDBNAZEmCRJhrijuFSBrrBoR1P1dpR3doW1SnUMhenfN+uOTCaeC26AmW51h8nxktJarV
0dZooyRuExaXKbD7nXJbT+qm5HqCx8LBCaMwoy4xO0L4ynwtma4/sqbFaup8fpsQQ0HPqytQb7NP
YQMhNJaOzhWekSewbYktqLL1r3mfwzVO/WmaG3mQ5DyDeV8QlJU6fCdLGIYaBo8paOXTRpJij1WJ
5tXbbG40OfUqWXnGi2ZbHqylDyMxIow7wdom/u5oJnMcy70uPZaFxH1Npdx9toelCQohVWA2ohDh
WHYmLADqkUd3NgcMOufFZEjREPeGzBpSLBmfnw+W+jSmRmFIMYemADp8IzqHfep90bz0uwHd9MWQ
42GeVt7aqlL/A+TTOSoEhIXuycUG2Y3oEKWUq0O5wHZhO8tkYyHgqqdsxAIxtO4MS8+T0vvYZPUe
scTcQNL0/zvtUVH6GJ+Dz24JyhcEw/jWRqFcW+7p53fuP5mwSivMMy3tzDEwORiBpCR8v/P7YwPB
vrF/5BOfCUD3oj1Q227VG8Zk+uynW/Y1JNuzqG1tcNfCio3cLz+RVqSZ+KF13PM+EzSdgQgR0YAU
857fSf35weMq/PLLC3Js4M9nNqHFWHvMIX2BkK1/O5PeIMXc8bgH1kLSrawj1gjmRGHB53HvHmZu
rKcf4vm5SQmXc/C5K6fhnzSvv3WyOTGwDbnl7pz9jUN5IvYhLrDGpbpOv9wlYiGd9lAxuO1gTY2J
WSdY/me0JrK4qS+6glDGJIFuG4GFGMs6oCOAnw8VCUMIfQ7KMCCU9tn7Mt97E/1FDTWhiPLH4GDa
PCx4Rg3qRMNahBs0nHJF99Qs3gEg5jxUweZInI6LEJiDVIPkslKShsU2oDF9KY3a9LEARM8ko71T
n0q8OAWLzNF4lOFCwH6FYcCUUpjvgLpLqjnguDQOwm7q4Ojl4X3JdHKTio4zMzuf74uIxElxwdka
HcimrxihgTMKf0TGntrC1awuYpEZmFYfFTuw6xeg8ANDk5yr5Im1khm074m/YyoJFNYD3233tBz8
2LZZw+SzGSmtWGoykoDtdHJkE98zl3r4aIio61vl1pXo42Rk0kV/QdXVbw9+HKuup7+VM5rAeBvN
GcBWBbNo2o0cBZuCEHG9qV2EjcnFzWQ8ONMNqA5dgsfLsQgXDwfg86wk63v0pg9IdZRFsoqQqEYj
JSj32kYEd9usUqsNLC23Woxxlri7oxmzTciGHmJQgRJKQThiur3npggjKgBcVZMTpf4vGcR23A+w
4whsGSb9pdcI0y3xs6AlcSN75INeASkWnI3/3ExefbHpmx1rsTO8tkDda6pTJ4Tr/NikdB2KzM7q
HuacGApnfr5FZHh4dazDlDi4w/ynnktsMsYHyMLmbf9ATtp7Tk8BGaUD0AO3BAKiKwbpwZkbed11
ZeBuiFpfjqHa8oGWsk7Ah9R8terq3J5/0qTkxEKfAJIVRFEnKWWcjGbf7gd5LAdm6x9LQEb8lo6s
fryCRdQPg1ebSIZ0omYRcVuqJiYgaplKaSWGd6yAmGVBCAYCcaaLGuXjLrjiFEd7t/okyfSVRZSU
26AWiF9rRIAucZuFVT8isSUdcpECsJ8tWtZqX0Hp7dTDMy9vP8cYd+OyBI3pIXyTfDS6FECPB/wn
eoJbyV/KvZsM4ck44iE69kh+UxINKnCNgTunLhBZOsjkTnLMcHjxGRTVN6xO6ODe77LyRE+EvHf7
UpieLHr3ldYb8hFcinqVsT+grUYp3H3bUejH548IBslM3Y03y9DghNSlUF7ebOVCkg8afF7FqktV
1wESSra3g0HGUPta4QJDIYJ/tEwKDC5izWvLrquL2oxSTP0mCObXeSWyRotWpfTqqXozMkx6v46v
z7D2YTp3n7ymegLSEn4BDuvIvxSegtzBRHvms/dGx0JhR5SLcRKguxz3kiAMmZvenIv0cC2sRieU
MZst++2K9BJFHg3FYK5w/h65RMePZMNGOfoVbn4UAq185DMqDbFA9fHVDN7a0hiz8UC/mmoN8QuY
WBHoeFeQHPAJsewcvqDxMjyqEddXGFiz5SL5sL1pDeMxEXONamphLNyEQ1zdv+Ov9/xv2ChEXDEa
10+pksMZGPfOl3saYuq1AvCQwGq1JgwnTe1ufoxKKQCNfUraEGnxwbtiex9W+6wi1pHMuuUn4C7b
USFghNz7YhXn3dFYlXaxTEStPvIlUgHfQ+zsDsBH3UURnzNO4ZOAOMX2uVHcKARpuXtU3UkhpHTL
pzTRuNenABT4ar2zgjF5tlyVTJ9+n140sAXKw1kffY4SHQAGebymFauPB9OOPjUjC7JFnzjj377M
KDMbzTtrnM5XmI1a4p+9ZmlmAP1LZ6OF5m6/bFgw4soGVKI+N49guA0CTY6XdoUfeTGZCI4xH+Jr
HEROBwwlajVFEHJ7Opmfjj48jGx/JERw/r52IuR9sqfuXreKn1vGmg/wlJ2LQEmvlp7aGcCbo+hS
m1S2vBTpnzmu790AIzwvRlviOtg3WUaNaJviD2R4R6DcBddFI56IzPq6Qd6ss8Rmvw8IWs+XBzEr
7BrI+9OWjr6ZAeEcUi02dwp1mbH5y0r4xSvl3rIR0bJaKIQfN5K6/osE0RPw+FPqsKIQmAhzV2TY
m+gWtysAiN5MX6+/QLKN8WzHycgFUCE57w/VsFV1UHoFOB1nqCYEYz5rKM/gPAVLj+GQT/QKS2h5
tTyNVoGlqK/nzZjMbucI9o5cds91sGJWGeTZ7Z8pjLL43EpjCh11w2xkdfhvi6G+QQZycJe8yICz
vOAfppRjFwmukWzAMxRM9bzypLpxCFLPsuuROG4B4XxenaPPz4zdlapNwSw86XucVvTQ4EZIojat
Y4v6qIS7uXfyGnH6zthD5UCZViS9PvBSIiP/D6498QB9ZXQnP3c+UzIgDF1yvMHBolz+YpwDxNvM
SyM3oioH5MDAFqk9e5Q2OEp/9l+cd1s7ROkSTdyhbxhsjtALWE8sz3voomRr7+hZUEATbC3mgOPd
cdA5MQ6jD7gjMUXN9eZV8hScmgzQo0lfcdrpdXf8Uacje7AjPsKiICza5t11lW0RBl+XBoyHujLa
Ip97l0Bgu8sWjD4nwwyUlCGffzVe476LSKxofEHmtA7C4NrklbeC2qfO11/uQNMOCGRVMZU4I8a8
gLqvhAR5+2cXsKfhJpT/zqW8T3TSCLB+eADzDIPi/ktutfUXIw39s7b2JWzPxR/64yQp48k7176Q
zOes+pndWpKbwhsPEsQaFTKUs/HLxvlVi2K8H2ceATCCxlLV/z/Si3B2TwbTC8+tXyA1MFA8HeXJ
glPyANr901UYGFT97zJKX8coTXeje33vxsTLK1kRUSXHg0VaPJjuYPKt+nbg0vuisaKSbiuekrLJ
bzni+Duq5Z6navPRM6Z1D4mFKSz7Ty5C0IVT5ODZ9C2cXNvCyi85sghiTZyJWGGDQI19XaJW6/Od
eayJLpyg71UkqBsCQrkwsW2+/spYAX8qtJvPWPERemnuuDwCE2ojG2zHeD/WCaukghdjn6U9CgzZ
LUJlhYmAeKFbpQfBpqt+Ml2lt2qeJ83vZdp8SB57u7jBMqpaxhNKQP83oLnE4VpTW5cx4PGWBAqk
aTFqNIudbCB+xaJx/C+w4isGDVON27r2LSmi06lFKlNj4h/DpK6AaRgy6SWSVo/SqnY8JeZ6fWMl
3Ni3V3hl/AGmsyg7KcMpG5oLU1qYnvQUdOW66Q8MBc5oxtOdXnRdO8lkrV2JFjXwCByuIas8ZU5+
fJw6UN5DPCa1/BYXI9StRbrz8PHex+r019piD0HK/2OzxOc2VlogidDaTUHs6dl62V8shulw1jip
SOZJYoZ01hDvVXukW5sW9lYtej8gEIJ6xfLV6ORSnvKtnuqC30U8+IzmrKkJSGF71o3OpoKmYlwE
O7WpM5PJBB/eiFcg2DDBKqXNGLDuo0+FhPfcYTmBmWM+PnGSlwlBD6ypJDNhQAbVvZwTCLd0MAiz
D69QTiAkm4Aw/xsuBDztqQIisa14GoKIITip5nkIwoTyAXD4q+IsulD5tNRoGnrLY/axXIYJPms4
sDOvWeHvUaUjH4W//Utk0IUs5uqJw0lwovCcPFzfhFC+Hwk60c8NJF3n4xg5w6K9fkK1SL1y7Xtn
+pbz2YGAIUtvU9kAOQOYIqHN3+xTmPh+hEnP9Jqzy72wy+KORnuExwGi/WdKuKk9E7b2aV83WbpO
IdZtLr2l8OjFvsV+Ej3P0PhwiQ6tA6BX5EDAmPRgMl1KjkNm8Tvvml1DPL/0Aw5DjebmwV7uyr6Y
9YHTtZDZrbITJ7PNmLDcN8H0evE8TlQTg3O3/bTJapEnqd/EDxW4906/oVIjbTc5roxRqhJzxHVd
WGbOsfVMW1QdrxYLkCLTY72u18LIrHd0lbvcZkhbY/oPup5BEZtbdt8vzw31MSuX3AGRlWtmhtZ7
Qqur/KvrDB+Q+jakfGaEtazNr9K5P/zyJVDhxIHHLVMUHfvWG7ByNwsV8yCxFl+VZXaFRmcDFtQ+
vw59uHOaKu5M56CeAjOd8Sxw+HkCljftBfJwZKpRsgAoU6dfNi0qUy02x1oWbMiqVHLNA0iaNUf2
6oy6zR+Kpj3DifxlNO3C4p6JiuhZYz+BRK2RF/2vmPBkxBdgh24m3C/QRiZXuDr+4gA2ROeMSdPe
m2dIPAX7rvnXedVfEXSMfAdQDmc1dbvKld3T43GANOhwgdIwr8irarwPmlMTFttnidwAlU54GYMX
4xY2coUsItFdEEigzSL2ZqbOfYEsIAWzYQhdv6e0rAvqmKZixsL3QYHYGibVQkErUQI0ntqZZXEo
cs1nfQ367M0jchEZd8Wa70zX4s5A1dMMYdhDFoTGwn80Hd+Xbt7IEuBNoD3zzVp86Nu7eeb9CeUu
9lq0TSKLR+2O5JWgbiBK+1VQQg4pvA+Ka//Tc0EZ4R/+0M8uXbKOh9ElxsbNc/1f4mma+f7RJ2S6
N4C4r8TcLpY1vLve80Csko/8zHUBS++55izE6zCJ7jwjOKwyzocgKrnJRE7TJxbZmHLrrmYDWb8e
dC/wfqj0Yz6g+kdgtLDjFaR0IzWE37gWFoQScpOKeitY3mILtfCv4sLJ0TXuzp1aQ/sibeSaOU1h
rs/uQ8lRNszwtA46XACvnzJQrye/n2IzXjGdIXAF5JougD+jjeN8fqON5ssgddphzl5kTBv07Smw
A5P1Qt13T19nUKco6PXa/nmKTaIOQl4orhodLwrHEOvgGM0v9GvURd/0vdXq+eyDyzZ4wWs/QfI5
i7ZWVi9hU966nfiBnocLCok+00dP4QEheF0dBnerKR3GcIRc41vX56sgv1mCQSAzuz5AyrUqIC3A
UFm86LXvPRWzfH2ZlCEziOS4GyDH+e8L2I8Bya7+ZXLpC89Bgja42rkhCRSZObi8cU1JShBgWHVv
tMqXv1V75PGimrz96DbL5D7JfDsjvkpD5HIVXa8cRLu3jHDC6I04Fo1+FwAVP3OYgKwpm6puNqNb
7trYr2V88uOLrIc3uuzm7jXNQflO/pQTfGdy2mO6yfA/kQ6QA0i004MfbEY9RqzSfvWvTgerBERp
r2RZnvTgPBlhL4X4ksWImPB4J2Nt7bArwQQDbgg3fnRGMjzXP6xsJhdau0NZqKu/C9cZd7yqUwwu
yut0RULtarzdV0KdE3KdFRNBOCoa2ss+436dU8BVcUm54Esu85JFaxDWxV1jhFXTti2r2XKHGD1B
C/qKnGJLxFAVMNMsrAtFcoyzqvOAuovTq7qplrUExhIMbgfHnxVQ2HpDdHa9NgrqgSc7Uu0ditn5
VbrD9rcYRJ3XJP+0lGAXs8+DZeEarAQYNi9YDJ2zzmaXXoNe7Ur2ieOt2usgjsGVcJQjC4b++k+i
CB2NWbcoZhjLdGY05fChz3oUFAidF7vchKIpL1juXf+TWTp7S+tdYwaN5ti/ioVQgpFlVyEZiBO7
HNT6JdneYQ7RPtNGLtfIf6u41oMXedfJKXAKYXY4AHkatBxTWwCtGKqSl1VeWuDMZypR2fKIixQW
kdvBIHDgGm6imFAFwt8zPODtim5gy5XkWD6/XzKLkfCek7wO6HxVUjdVcstx7ndIESxItMU+CRxC
eIxrAKvOy3vFa+fmbkU3QHG16GnA94bHz6lu8JEXP+sIWYyYSIiX8/RWYzXgnmHM0V85kJRU4mRs
p2Ubddww/aysyFoJYsQF0nArqGZjkZXFzwyM3z8q6ZncjZP7XVwWGR9xoj6/R9y9g5Pmx7W4luJE
fpyCsLBUHWBFxn0IpL5Jsa1fRHTyoAxViGVQJTJDho9uN+QVwo9Y9Dtj8RhQJrCIPpvCYqeMptDF
djT0aALJ2HmXZAv40a1RPp7bH49s8JOaQIDnDKAy/EalFadHU/WJRrU4uIsVT1ioRXTe8G6Sb24N
9iKftsoRN6kWmqvXmHI+uckvSUzkM9MwNvRQhHkroWZYL+XQCqHx18aLgdBHrDbVPWcNdzfmXnaa
5T333qSUtACQFVKRA2xu4cd+HMLAcd4T6B5dsW8fAOfdnr0Z460pf+tyT4ccHRwT5dwMYXTFmXEe
VWWQN5FtctV+rCNdBOECIDS1C7Ins3d5TsPmspo/2FJsPMr8cOTnkNffwr9wklxI0KZHM7i3oU98
H6W6rVvsMkP6X/zaV82r3PGfbBjN1FuTXV0WhiudrHLgN3sFcsgzq66B26XplRO6dzbmWTsCDYKl
gvxt8YxfXotikxVm84zapBfRCOV2OSQk8SZ3O5uh995TfXJ24dVx8c6jBkD4mkNZwaQIMkvbk1a4
8nCjqafpwjiyXI/9J2NamCMofZOtISUVdJsboj56bp0afUwy/dBrvjACsLtY/bfK9VcNQ9AFnpJv
+Etd2FtvYTQIksctiDCIu80Y0jsxaxLobYvqaKUofNHcGa2a21VEGlfJMpiQ2oJemeO6MTrfXVRs
ovzqunXNQWf+GSoQRBX2YhLTANiswni3lrZ/J8wRr+94NtOTgeo0SxZtC+WItCtwFYWLX2omRlTf
bmXUi7z8MkMaBp4JVw1y6DBma5P7skuE1mfCgZcgxEF2VaAqFo2AxAilSHJH3INuvUtu34NOgHuy
kUeCPcx33I0CunSGA5uVQnky+yy1PeBcqpmKxEflriBag7V8htDVUYU0KKw7BJeQqjWhGKc7T62X
7K5v63U8wfBTw2e3E8W2VN68nL2WoL4b5yccXt8kt2uv/gyemk1LqPsnDU4inYSVtLFuE0H0yXL6
w0vsGCSY0ko7FkVFRumUCw6xd39/cnKruJjDqTnXPxAL/koHfcUxj7LGSBfyJBr3RUPVILWRk8yL
ZM3rR2Z6O3ecKPNYbeSnIvk1SCfr+8ho8wC5y4BoAfAZhGxfJRamJtCQWIstE34r+wg37rm3Lk+1
ZslFG/0G6Z8DVN1pibCzVZsA0aOQ3Nkr3oU+PiqS8I1XQqQFIRIAk6UJSzUhbs8z2FuEH9n9L3OZ
6td9weVWsBsiaIJvSH7CbCIoSmAJLqXAs2VijJtk/8qwe1Iq71mhJgU2DXWvmLn2Pb/OxNjDhIcP
jhVGMvvWkNqLf9Nj5Rxx90mvfBB6L0LxiU02DAGX+fQ4LhsbOEJaHasOoVItgP62+zRUIz9tx7dC
PfzJSlCiSsfmH9qmoUTjth1x4e/0myCr0Lw4pD2Qn1MaLfhCXeI0C6amjKvXo/bkRkMYYzMHeH/x
9MYSRd1RUO/RTk64Gj7XBpgXHDAS+v9wmI62krOx8dxu0l9XJ9P53HEDuh/4jjKc8G19lq3DnBZp
Eaqx5hwYItlVxIUqgwEm2620JOVpeojH92ozfQLuQJR99eREbdRCElzLX7BN/brikz+jTSy5dn47
em7/uVFiD5uzEmqO8oQIlxiHZ61SLio0gd+4RdVGInk3nH5T3xiLdKmiZgkvbS5sO4PrQISPWefO
BK38/ZjGAZpCABfYm6uuniw2tmWWLknLs/XhONM+6QC8RkywmUwptCQbyrUexhpQdv9bkN4NF5l8
ZqHDKIhw9FL6Sm3F0swawYumzfq1V5OyeCRhP5xKLmhEA2Bmo0BXhWdQ/gkmi/HiJxpn00VjV2Ox
ptJN4FRnxoI4nT9lOYZlHVDuRHo1aKNDC6eJ2LhD52TdjzV/8WWjCGBDtxEcPiHT9FVKxr6/q3Ot
f6+VKXpzjc0t4w820iImrxWrO7UtErqPuqOd7MWOKV5DouLFlIN/7oRDHs86GscAbxZcD47myJ3I
DEy6vJ8ocIZN4vTMAZJVImk7EX4yoATJss0VS8f7W242/iT9MZlsGSVn2YxBDgkrk3fNSHiEIqXu
qeJTD8SoGvHJx+lQuSlyVuNJlfICbI0EMFDSF5hP3rWQWzTtm/sxKuIvvS2dye03a86DSsrw76eR
Ww09R/vB660pHyJsflelUdTunF8uKo2sW9YEz4EwfhCft2oltmfL6UfwpXCT4CBK0p9ZM1jqEBvl
hy/VdwQfxHdpLhyk/TQBof+OO2s5mx3WaBR8CZd5jrYJnNG1UfWI4eXYC+HoYsp3RU8vMv97iObO
DBkYdTqKaDPDnmKqCHy8v25vw9qNvF1GimLnwwJrSbyZmGFQ39sHIg1IZUB4isfyvRTWp1/WE/3N
ittVQmiAxnbhG8aHvAumnoxXUBAmbJOerx/M//qF9XJlmPEZR/dNnv3TYpA8B+bBPkRny7a1hV0W
Wj5VPyKzxXrrcrkGP+aST3bbchW6GG5KIupINv3lvbnCqWhUlugAuF7kZitgRocLeiH+KiwVMUlF
iyZRdQPnnCr7N6z3RXuZuep11i31g7ErHnFGZuqXRAG34jSACDv4j0sGSkOfnqfpQLkTiTUWKhks
PZto3iMHxwifh4KjDZazCx0vf2KJBkcperpCJIfqIMnwmnebnhYsZzUib1rSh58PsMmLN4AMNqow
7SssRpF7Ho2rWAmHD4/HYdUpa2JDzXGCWuQl7/fuOPHlb/726Ips+I6VLYjbeGgsM501YM38w+0S
x7SBi6UY2CMd7GHLPZtBBgRqGwzap2YxvkQYG6K/VeGw4Yckkcj3Kcw6tnW0YBzuuI5TGtlj6RUm
BnX3oEsRMVwYOkHC9f56HgO7glnoWqR5E46EqhG8nT3EFqsj4+0kJYT+PshMKKNnFcMQz15lemXT
S0a2UajO75cprwPWsjviW2KhOCzNd3cypRPrN/pgBim1p0wM9e0hKZZcQyGZOivbNW2Qz6qD+IJc
BTwoEAk+zsuoUpZs/8WYzDTgD7EUaXpd1cCtbsBy8aQcolBweiJpLJvBdZ4Nl4eWhI6e6Hw1D1Ct
tzHKdlawQ0XjhZDqcHenKDjNTfkyjqID3OAs9Rjw4M/MR+MqDZoG+QdiKdk7jX4fCjhYjhc+rPcL
TCHvBMFPhK8WPNgsIe/3pMyjzK4zuqc1h32LVRAku9z+r8MVeKpd6jwHfN1jNNKFSJKe7DiHcCkK
Z1/IsA941uAbTVag9J9bZFZeocNOe56WKqHIY31ax4I0VmS+jh+/6sogShVZ/otx02KEBRdD/sz5
mO7im14MtceV9qWt0EUHfuqWpDASSz86Eu7A4zeUON2aiNLgK5g0+TrK5VL7/8rECjWRz4WKVdjd
//NgjqyrU6eZi+0bZkBA1X0505E6YM0E1Hph9uj1oGp685O+pjxLkknigkckQ/gb6FoxAOKJUsb0
wSDFahuneE4O7Ycc+biinFHkv/gZ3VHQ5vFrjaFnuCJVOLygHHTte61e9D/pWNg0URnxC6Pzenaf
VfTF3AoQLizfeNonvGsaA2UBwbdLX2kfVl4OSmILpk9cJJOZ1kZCABEpDazaqG+8JCzUOfSOyucl
YjltZNmYsRl5WvqBR6mG+1TGx5rgatry7mh9FCdEqcYDgUT+FZ2FhtenQJqwDpzP4MuOplgpdTCG
xSsnvwMdqSifIYihGBVzhV60I0cWCMgPK4TOrrI2mYvtkJQnG8JEDTzOPsWAu1yRStpjil9HgiZn
8XbQ0+4wZnoYDzqa9d4o2hX5rIOaSPjzBydN1Y2AF5rfOHcd7F37biJqloD3fYF/MY/ZvdWV6ilu
fDEqyIFEFBsubcA9oTkRKTvCZAJbrx/CzCLU3RvaAk1QJ5iU9DrcFDL/XObEZWcriQSFkgqk9D57
JkUpw2J8EtdkjleNT0iUqGB3E2EQ29tNxIEbIZ4yC2xNDK/iY6AvkKujuFcHvizX50Uk4xloYPpG
e0g4IyY8D/89q2TgjSr5v3KyEkfdQPaQ/wprHB4W1mntazMo63GJrI/ocX8xBYq71m0ghSKJX2gj
qe3d39mq07Ctlt+54Zw8VtuSIeIQnjLdyoTXmyRR3/SpaoR9jlnyzapnUu8xdS9MmKRqmomMC5Wx
VvUGNvz2akuBy/vXcGIEzpkDyh54bcdDxHZqCAceWlHS7a32utnhjV8/kTWNAmBlA9UGFmabXxic
i37n9tGv6AwsHAJ+CiwNDOFuAMVWlmNJB6TUPt4KrHJdbLPl44wcErU/2xmiBJTmqCzRtFWOrbZD
Iyc4AnSfJXwxGqMga1xqdwOGLJizljDwYilZcN0aj2ozSgzBfGZ1Wosrip21vpt5tu44799wENvx
feViAU/H6NUjeqKA5FoUoUEXH8y7B0z/q8b0JWFNdrAEJiECRt2gIk6v38OgfAKv0Wi+LLA0YrHZ
gvO8FcURWVjkGUg7h3VCTsJ8AmakhZF77sB0yyaH6OkRzwlneD+r8FGMA/r9ZEtHIWH0Wm7SZDpy
6S/m7flbrOLz5ggRYwBGPYhppzSpy5JG0nTK4vdZ2sCn/oiVsQWVdegTC35ZW7/OmtsjPr6322ig
V+DBUDOTzTD4DllQdakmR4bbvHHwuNFKW9/fqNviEOUIM5V3wGOJJleT9aufxgPuuCCKer5U+ai8
J3gbACrTnRIKAV+BXnTcNGVKk/feVq2MWo8WP6q7LCnNobczKNCkk3PbwT4l0GXOJ/3ae9e5t9fz
uFXBoByVALncbblQ+NsIYW81DcLiNnPPX6vYCT/4rO6fZbSyCEPzSGuKtp2q9olfIsC1TPlIYipq
j4dDsAGbpMovqdKvmNMZybunETBzmDNfDTX3KYsc/qLYToNjjIzrnP4DDO5CZRFZnQjBIqH4idlm
UdGfgpfP7CThIvNadZ9P+yJbg8/mkDLSxn8ImUdmdzAT3PfkDWvtPfewHoer/uZjdkCq+100Ns9R
YZG5LJs+4Juw53Z6Q2ygKKYs7sqbEJ6zZEuZT2n6SBCLAUASJnjK2uKYzLfYyZp2PRXw5CXUsx6O
QTFtaiX8jJXh211kSXRco/c5dQQXkB+UlA1NOrhexTUM5l5Iw3FXz1i5fr9cgQT7LRTkB53WbNRH
BGmHySO7UcZR8QOfOYTTZ11xWkmy8327CZ6PKoTxOBwdkX0bARJIQlrLhI89PT6XAH3C6V60zkjB
J2DZh/bBosjMF0FfLCq8ZxsjWTmYkVsbj+aNcOmyUmgEe7BiBbpSAx4uCt+BRaZ24/YrrxVMMfce
F8A0PPGmzYgF1je9Q2UGLPoi4ck6QkGVtUgRcOzLDD07/s5o24q72aOJZHgZIIuyL8AwZh+eBFWB
OVLubUrACEjIyiDY/ltN1cIlnCTQ0nH3y0GODp8bTa9BknIvZPAP40idVRY9ErzTRzhgVyamcNjP
GQpYmPKWr2ckTnhBKrzK36LMsY+o+JOw/LsX3fsQNEquGAzKqHeBSGbUjZHMQ87EUtSiMlc4gmpz
8I++7mNLr4Qd5JJ/AYXLt7a2RjOYynPsNiU/xkwIZtaeFkfiDY5TRXXWcFoviaqZ0ZnvNekUnDpW
91zTIFpkLnk0l50MoBTg8a/8XapU3E4GcZiTMhNmAboqyln/vvagmuRxiNbCJBn8qNW/d46qBPLF
o+41Rt5o5oQZz8PSpojGH8aHUYbYlovrMii4JH8KqCSqUdNnzk9tpGDOioyg0ll/Z87zwJkRXIQ3
/IqERQg0c9akARnoClp3YnogDxnAvurqKAPz5D9WoBzOgpebyx3ML1xZ4+3JhW4PCZ+JncamgqAI
9uC21S247DlEN0zmn5BjSe118/8ADk3IkB5owstZzpsB3GQvdUTWAbT2s37UU22FfqKmwdaLGCsF
LcDNymm/nV/C9rsy04nMMmx4BEQMc8hg0QwNNUFqOOiCfL7UnQM6Q8wVFzHkBEZHn3yTswfdIPVD
Bp9Nlcadg67ptx9lry+n9g8S9D/X/OExa1OR0wXwHk+f3g2Bapi8qogy0A087Bc475NLrmKu/fr8
KnjJHMZJeDAbIGWWn9lrPZvtrKv3if7Ir36u3i0eqYjjdfXwE235Lx1K9005NwLiQ5/yCZD/YM5J
Ur5W+o/cUy1wYTZ8N1i9f74sa9Si2y4SNc4iRpt7DUjv9t8jCJ83DBbmmoZByL3sWJ9I5y6F/GsU
a+OQ6VHhgtfhsfcT99+tqEfh5GtYFynso9kJvbLfir1s9jHynkHVsTdozb9/vCKIIs5WJoQCFUyX
8wfq9KGV3DA1kMsopHwtX6fwJCENwfz9ro0Uah5pBSkJdwwgsC6C4lvArXpDPkJUz1Od+m+oVvWG
ikwsAuJTFc2mm1S3UYU9VKMxDv+1hnM9gNPBdegceuodY3xlecBSS3r4KZc6jv0VE/7d0rY8BWsa
BJSBN/QPbdQAjQb41NDVCH8EOW0Pf/VF43w1WFLgalOwiY6BFuqvA3FMwFxPiFzRWbE70OStG/ae
LMJH/0OFcNbzgFSjs4Al3+th7mWDncKIJP7V33zW2Cb68FbtgD942WbdNFdYk+Jw+Mao+Xy5gqWR
mdvuUujwkEoYd76lXoN4hrKVQ0xiIWpm6TqtffzXW8i+txzZFxF/42L0UkR0DrH4wxe+8V4uvAgA
L3XJ+L8JK8GQ9fMzEy4pmHA38udadgDxNxteF5wrVJI18Dap2agvEbltNwUqxgUos6Yx6dW5B4xU
OhhoDlxLjDxzp+mt0e1AhM2fHvpsIIglmcS2SHu4iJqJXgbEbBPfu7pad+pfBlEmVbRslNoV2C0H
m09j2Y3weL0MxZSazByjKSaZ/r/+6sKc8xPwKo+/eSlxwAU3QPD9aFWvj0dLTe7z3CVT8ML43bnu
VzOpGsLANY976ioxHEWqfL7GmGH1pgRUnc3lRzvIKOnVd43LVVdw22SwXZGqaDuevKkVVOirPSQK
Z4cvWgCCKKhQhQmYbgHLwzQ2W7XkDohbl1uGPAZjm9Z0SF2BYaB1KWzuHz2FFKKW431daTT/DJSn
8MH7b+dE66kd2N6RmAiXQ+PQKgGS4mxD6O2YlS0DqY07qXMy6t4xEA0t2Bh6cgtvtzVftWbkH5NQ
CplZkwSVZ2XkZHPnp4FSeAJy9/H4pIBNH216UilNM7t/+/xtocHgQ5pBtkXQLNM4ddo7wIuvo4Qq
8ncVh9WgO0GFNBFUPDoou5Kht1NHYGo7mYtDNRsDYcmkr8iyvtjBo6K+yVs8Kz9Au526CcJ1CjUr
quaB4FOBmnYpHDmJQ8L3UIsGci193dfIdn8m0zNYtW9GK6u5F7UmLdTQh+pv1ExaWTAjtPi/5S8P
V/lo2X5xDQT5yIEOoaSCz0hvmIUdfSepoTWmJF7WQb+XS66C/pIjGQ35tUUeOi8+s1PMO0R9pmE/
itYiYBc7O5nlkI5Iim1SUxGPrEN6SL3n/OMLbX62ECUFFun9IPCl5Cm6FjJUbSC+1UqvlyCiYqEC
SgUu/31CJqe1lm5wozMTLrSOqg+/JMRNIo8lY5F1XWlcX6A3eyCQa8Rqq3ld9UEkqrtxpniN2yD0
wxyiUWN6pAoxOEqF0VhoU0Crc4oHCKKN04bpy+YWFv4uRi8QuzN0PVE2LKHqLxpG5/Drf50W2Elv
dDIjmr/GtMwVe40CC+ib5X+kqhb6XMlHxyaDRU5HxVUs0RuERhuGHz3yLn/JtYzfDNxAdvLzHQAg
XgqGqOneOCI0NqxcFL3rbD56KO+WalTEkkMMBUMpVK/55junBVG+Usb92LpIU8AY33uyEFrppyMS
fevcGdk2gAHE+PsmLE4iADU8ZUDm83rmM3N6MmZv+rbm8pbMsXQaa3sb3K/BYsS6LKk+L6E31qLF
zW/JJijQSKTookl6/vVDwnILApwGw1IOBBdVv+xP/boDBMhIstG8S7gqQmF2FSj0TvFhDx0Bkdro
kTwYOR/ZW4ARKqrHQhVcd6zIDTPIOpHjzwG9X33YGVGgJ+MRtqoLWV6Kn0ObvIKWa1VAsDBztRkW
NaizK0eZxXRBQj1gj6IKngQEltHMIkzDPvzC3bT6Jz+VXEpJeyP5MoDzLdipUoWlhthKZqFC/459
nhe5D8HxMV9w9i6gxVMJDuX4hRijZCMeVISvJRnE/Lpe7Ebicu2QlfmMGcBBfahkOzxWRRmJaCwF
nji4A4dqWmyy67hKpWVDWz6n2UtrqjE3boDy8h6YVL01Al87/20b0Ky0gtieOek2ld7YAt0/hLg7
15qmOaQY++OWuRlo4OuYsPlkKDOb+Lro5Jr+LmUUWbDqqy0ni1YMIpL3izOJkGJg6RmuLiXSmRbS
JWQRKnQYCHL/UHTdY7lPrgbZTZcdYjH0bIPU5JNTE4jTbtZyXGXWxq4kmj/zsND2OpzLdwadUfo/
kEWH8P/AgwRLCUjABNe3tzIji/iVdeQDxIDqHDQX4cZXLrQB4l5A7UG4xKIjfB1NTwGaDwm7DTQi
Guhk2hcDwBTsHMqpHt3wXBOsG/9k4c3Llf4xSrtFb3PAZfss7ekMiuIkDY1X4thINOW5cdvFzJJ6
9fVek+TJka9YrLwJE0JMgnvWP3evyG3nDBYgZH0ler+1xxwKhGdwDeNb2fxhtjYv/njUvkdWrWEg
2mYSOtUkFW5yqmCEEZDHe/HqLTP2jDwVmMEN/7ZbjxuKGv3JTorGhiH5Z941/AGGZGVf4U2p8PQH
+WP29nBPurZpbiD+/JT2ojFEJ0Qj7E5jc16oUlS++MpSRDkcb/basl8lqOpAL8UzX4yxLIfXPL4L
dq9XKEIzFdB1RDegBoJ1fxcP4ksIGExCqsy+crLmvuyVidInwwH81lm1exC55TnX1BSDTwvp7xSQ
L9cc7nMPGB/MdSwBWrh8RK4UVaZWiB6ER1KVdwf4OpxtDGD5wBWDwJG2CnVZc3JI18FInWGxWN8s
bpTS6r0zYUtnw89irTo7gUbiI2t+7Yf4ZMw4Vv2pGgfoVghfXmUblDCf7JZ/uGd5EuAKaATv0bXV
5Mf4fVodE80TprVtxMhK3gE3xD0gQON0kl/MlyOrKypChuXD/xlGkjT1du9YoW7MelPP4Kq/pRri
Tfrrj+ZKX0dUTC+L3KThcfP91lS4cBsBhFn3XyDcMUAjEGnseq9I4062CLZ4MeVNufE0rJvV+8mp
0dsUUpgfCEjDyRJYHyuzDve2JRCxIqkmPnI/nA1/J3OtHU7scsd6yYNM9mdHK/kPRwUyordNUpEE
McQifJPUb6J8IewAbgRZuxCxQ3i0oV+FDHT5HnqyGYVjTKBFqVWkTzS7dIsPyxyaU6VbJqrIvqTT
C8rmdMwwcu2Z5Z/HS9Ik7kOME9N1uEyGs4t3WXQJLO+Ov0I7m8UiSO+u9l9APv1iFcZ/WUbaoVwc
GJ4atq+4YY/rnj6CqzSrrKYpmoANIL4xqBNgDZ0RGYHVf6EIwDO6Ono1NNj0tA8tpvWvCSMe+O/0
GNz/niPAkLfq/cxW3+lvjd3Pc8cjH5mq8aOFn85F5KMowFFrJl5Ngo+jIwagA3nXLztstTIJa7Gb
MLnEvToToYeimK8nDjTPVe/Wp5KIsOUJmGFCQF0bdNt2GbGyYm8QV8fb+usA3b45lpKzJ4zmVb6q
f+/EHq7wfnYN1NKo+l5908rS58cI6L8zaSqQdrxA06ZrYAVF56omEhYZiusnl/jFb4mW5Evafzk5
9XwXekA/tZ1IzqbjPynRiXjcy8FTkFt/5Cr0sMbuGCzxt8wq95+lRnUlAN+4KxIsdfGZ6uSFEt9h
P7LkitWCoUj3x/mzHsGNvWYNdTBMfmoJpMXbDMyBn+OudeQRJ22kTFH4Tg5QMGlPYxvvvpHATdjy
aVuVosWK/ZH/bj2x9Y1/TyIdOOzyRxA9/anvdXe+8bFX7A71bZMVF/Yf54WwuDVpPVVjS0YyZAGz
0MRnPIVV/h1Up52VFmJ4LP6qSeXoHJIvFn3UAsKDx0RIIXpmnwUv9QF90hB6j6FmS3N3pyXoITLj
7zOAyDlJpgR28e9BYD2a9abdqTWbR2/nQLny3yhcO/OdglW0Hc/UoJaNGHhTJZiszkEWrY1wNNG5
w1JZ4aKwJkR+NL5OwtOcB2Fk1cFf1AWBirovhxpb0Hevie76/5/7tELWgnKQVefa0aZwcp4vkNH+
j9ZKD0nGr2VL9sigW8EwHk6/ZiQUgVpWypYE5sMX42fqgZRe5bMXYLo8MKTl3sWK+A1UWwcLrc9U
Uh7fKXvhBET2jSZPgcxjsiUdV1CpJKYJOunyitMHk9fE1LRM+W3n8Mjz5YO8i8kAgUH57HngSUDh
3rhhod61/7C678nie/vr1/j19GqAl91FBhgX/j0tNzn9u6YbPm7NfmBCmyg7MoW4YuQD58nceYUO
e7NaU86PFMGC8N5jSdck7g3mhPvf1VmIXXS1yKVXxuDpqIM3zt5NB3Gh7zCookfaHuKcZk3zkCPj
BpTD2dCajZoAhV9MxFnR1GPYrG2G9+Oh4c+uUogMM8U54VJG1nBIoXyD6M9knm5J9cUHlA6naFpQ
TbmloUWCkaFr1gaC6Y1L3Oxinwj8xnoMi7Mzd2utL3gvX/VfkYGdED3haECGc57aDUaVpXaTV/EB
ow4Wu1KPCl7Eb6JIHfJ82wQGG7v09GQiv7zq6bIW3WHUxqM156g6DD26OoMWxnpfksl3U06J1+11
y6Y9VzPF2xpG4tq8sPLN89UpIKnSZ8YERueG64o6xWWkm9dmweN/Y8v46ZKM4U+VAU4cVVZISxYr
8YsK+r1UFUpzVuHIxIegCB/PqD01UOYkuTKw5NG98ccKSIKtZfxGPEEk+wTGbUl1U5qqqFCJm+FC
eNfTwmmQDWnAX24ifFt14h1NlZUSPXl659l2MzCvP5vZouXSGpKFKaNljCHXL18gqTrPywyBsWfr
gKHeOq2reV5wDgdCKWpix0f379FLrpbX4+Tfv9mSFj/W1KSO+EMCGi/S2bffOdSCjncIgeJay2/t
O6afnHkv0fJtcerxZpIKIuZB5zs5ct3BopQs090ZOuFyKdd+IIUsoxyBkmzlPdS36C1Ut+8FJoGm
whEaRdWyWyP+PX6QFuF04yjwN/17Uj4uM9fkv0yRFjtlR8KFR4SXQJaVdX50ovTbGXtJzWN1lJDf
eawH21fCW300FjBIDGRmEwfkepKkbllViIZyGx4mwzxzZMEE8zC83B5UJLKDnwCm+G6xDFJFFfiL
1pys4GQEjrIQKtpxqGbjT7a5guvTM8LGiVLhymSg+0XEHhiGQHF5SwNLllM7tM/Qj9xD3kuYOuzm
1u3KA/prLZDS9RciFedD3vK1SZ8j4dJIIG0uXOsRv+E5/rPOATYfx5YFWQv8BPg9O9MIrvMiQYWZ
mqFCfw6hzxl1CCxKb4EoHSqLiahPp4MZTcJhCg4rLSiWILk5b5/lNp0CQgfKIReOz/e2bWTZNHFH
r0Bez5ehq8xmZgRyEygz5p7dO8pOy8mSdApB+Kx5EMOf0TZGtiYFxYc1IcpxlsYnhPCFzhANNbZv
9nbNko8ftCuClU8c/ZnqcEHHrnkVQxvUafsNqmdIDGQ53nigmAq5qZLWAzfZzfKxQ8Ah8IXpMyD9
NHKoxmjHPZTzAmsXKjiwo00VRJ8oa+8YyiJBvWGejlbUg4rupYi29/tDho+w5C/pRcUrF3Ifrxu1
geBfhOC1Pteb/Pk/I9v/s7ZXGy9QriRs2tQXT4d1/SkJzcYwoniAzj88jW9pk8P4vOY32/3nBpng
iZYmlnXLDXE/BAf5oTvpp3Yfk4e6q+fG/JxwYY+KJI0aAGR9nBGaa42XIGwv6PKJcVNUgVd826VS
bXk8zK/Jgp7QD6P/xXHt3SCzX2XjQRA/GKuK8OOOI+rtfSW4XfZl0tUMt0gdkJVVOAEiFOk1fzU3
EtB7qFmwvLxWWG359bdgb9QO6EYo2Pk2FfxX5RT1vsJtE8Kc+tIxUNcb8hRnG1eceg4tIkuP4K8b
7KxQ+YDVw7chNqAWVjHIKGdNtM2GbCr3/1MNleYY0c5y3+WvQmwDZaeSssgQMCC8450qq04P6Y1u
fLpvCskKQW4a7JTalWye9eTVQvtpsv13vYpHPwd39zLPIYHbWQmLRCfQn70CRucA+VKRZ4HMIf7/
3nkYiPYUuwg+ntFiUl+zKWySH3etCgWalzrOl3vh5/BW8NzXteutmbvctfRuXkod5AZaHURYgHOm
yfobjSATNJWFeuE4pwwdtGZJcbkqCAtE3rY3/Jh006kgeOfuo5Yyurm8NMFMBDsXbOeWvnvufSKR
rXLZ6CGfhgqMAow4pOTuxhyNoo9OTo9fVuZ7RJtVMEePnymvcFjFRZ2vjAW2aeC9g8Ij28f/kxxE
j8n6SvzLeMOnRDOVM3F8tM5ielY+zKUnto40Yw4+BjcgwlPRvLdC7i3bv07wIcye1FYPc8rTsnkq
bbS8JOt+wXoZViNjYVZmPim0P52EYjz0eOaloQWC2eES2PcBSu7RmPtOzYkJTEKXNELKx8n79VxR
7kRyFl7aNQDiEAqPcVMimRLYxp7xxoRmHcxzkiN+Wv0QtGiQ1iDFi47aeh5bNkgbofgEiI+R+fPr
6IbFXGfmCOH1iL/MXq7cAalsFjPbH8YjkBHAseNtzqXlCsBpPBXUVMGmcPqDgjhgls5S24SruhOp
bKcsudgEN4yqLCyLSCI5yT2nMO4VRnPOs4accUorawQYVCNdCucbqzHHj9aCDiIXD9bY4M+gK3sV
J1WaJRncfnaI3NDBaKA24VhiAVbS1tdfk8vSWAL3YKRkdh3+Lv5EVywem9KWwPiQuPDjS5HTUa45
01eVRPX/R57SwA75LUZ/RGkrpRaDv91Ws/XZpxMW4dFW0k8AJGv5GSJ82ShC+QDARIGpo53+jbcL
Z/rv7GisJ+AsiVD1L+itjhVHe+20ViQEAOdYd/sasVFTo5L0w/eHoVmYXxB8AlC+RM1eC8Ykk1PL
p3iYrwmJdwWzkNBzUNDsuWEYMrnpSWz9cMbZjjp1iGH17RBOSySsPL0HNCyhprUekGR/BjuD8q//
Ha5g1DcFnp3NMJgYrpwjCrzmfbNWi9WW8ReNdV1r36aonlu/rG+Vsm2MuxnNdNtuI6S2lMY4ow4c
sUiME2CE/OGtT9PDj8HP9rBnYRvjk/W1+Q/6IO8w7l8wg5DKBYPF2eJn9EZlS+b2J70eRzppNJMj
uPxe4s5czrXRLY4ma+VOdFbp5u90Sw8Uj4ekjZjCrqBjX7zZlQiVfZzBWav6aNgPg16sLHE6ajlS
fZ01fYVk+EjpV4kNM32n2xokHQdOrvsKUGSJ6c6cPhBNdCWxycmu/tNxSFA5GLj8lxcINHtaoqO+
q4canwHiq770HTJv/SdIjsYodIp3qLsScUHSTQN0t61GxgskyHsG4CFa5ChWFYHYG8ijgzHYImNB
nEA3JnxtoSAxsm+KTsnS+u0t1yck7awqr0K7AUXVbIIThKMyZJfPlU8k8/dlB7goSWumvdFb78qK
VudYWQszmXm8GvQ83Kj3wHiudEx89BWtA0AKu2PWiyCgRgS9dV30cBeEBuVedSHTr7KvQiNci1xy
H9Wtnknyz2FZCR1fQDjP+UGm5j2gB9KXYQa8CwrzgBey22AJjAWmJiEQU8rJdZ3W1Ua5E1ZXEhMh
Y/Qmi1q6cD5V+fgxxapUhtaohOXtiJekWK09vHpqdXOmDh6e3s6ythKv5Teza4/aVZQ8qK627qQH
Dpf5GU0yn3B+TldcXTGece36jLBXxqmO2YpKFb8gxFgZniEV7rmxsPdXNoNbyKyTnmrUJJqgV+I6
7UKBlEcrGmcVmYHretvS93J/YLCFE++0r2tlOOdQ9ddgYcKOnPd2veRUxS0MB1ScNoC6+ZGu4FQ9
Lx7dT890oYLx90DfMc5T2ErwQTKx1NDxMpc1NL5m3ZbGO4jtPakDYZvxFm6t0BuBYxTsf9s0pYQc
cW1FxWH08MJ4OqX/zHphbRcI8B7xQgSOXaRAB/hPrvgXqsVWAEqdb2U7AKukD7HIsICv6PTiq00f
S639nG3V9Dv6rquzUDzVCvP/nKqUhHTV/GfkcCsaHj+97ZioLdXdHEHGkXr9bCu9+iV899OL8iWQ
qox8uX5PM7wLwf87vwS60QneqJ+ZwqUveP1Q1n+ZJxU3vM0xl+uKn+g1Xzo9HMV98UwCxFJh3QYe
H7RTOXMj0YiAxssssEevGJOZ/A8NRlCZ8/9uGu7exXm/3rE1HDOMtMYbih5aUYUOoTt7eX4OU/IB
rh/cLnX+e/Frxe96E8winc2zMkkoNmWmfnRcwVzcupxLmDuOFyuATMrd6lc6Um92L3tmdFFImrWx
D6SLU6Due0sbsx7kI0ue9m6Z1UGsiQka9JNFO42F45fIXJrdpO8IqJnAKi63rLA3O1Yx0Hbpeg3+
lNlcD3zBuqhnRvavJCZE4hWIbGB7wnLGji8zbqndKYzjXfFuF/x4R0LCNxFYOo8ioTPehYezjlyj
ioYj5bYNrXBpJR3gAvHX/mpJTnUbn41I3nuYxFVmzog+yeQJWograYh2whwWLz/M6vQ8/Z10OWdU
ILhReZ/JTYm8DibGZ/qdSiHL5uyifZA8+hyG313SKqolak98cs7UILTjA8vOg/pUuCHrWKSKklUK
CoEyShhDxbiuvUuJeps8Zf869Y/dCgj66LYmJZ5zuXiYPUBUJVYCm/Ft0tkm0BgOYs+FQrF/e0PX
s/FXFtNK82hfpaOPgH1halx3zV9+Xq3DPQ+/p2vHyKACskYSypQERnCScbZt9zoNTjLj4tjxq6kT
M4ds0my5KWvysfP+Mo9//b/MsNVivgiczk50zxtv/qwU6gMqA7VbHdNq2Bfc/0peMd8SM/GKP6Jw
Agbe7BEYZTaLEAmWtts8ChuNP8WTLnO+nt6nn3qJgWYtUof4nPB8tkQyRnqrhR/I3GKaZj1mfAKh
Ic06TJXfT87bTAfvh6/hZd4WL79/75l0sxw3nfi8bY9GQkc6qxn9ETx3HO34q2VRjnHKrgc5gQl6
lfi7j9h5SehfGrpNQjlPM6SF/B22Tx1niJKqIlsyepXO7iQrJ1vvLbSCB7qSRpEr0LA2AZgq5byp
7T2koYjjP/lSx5bMba94jQ6VZQnTBH82ZObIcQOo1AnCU7LdsrSQXo4S6dlvwsxCHS5XCMj6og40
Vs80WBiR5aurbG3e06i6ts17OunXlfvrJ1ceVCN88w7dAvNt8rg8Iykvva7wAc45jMm/l3eyDcP7
4ph8GuSI7PLGKsrpGIVO4z+T7vti286LolnHtkHnQqW5dcI9nuEbZxsOJirShJg5SP8xQaSQUS4M
BQzHZEjNdUWT9cs2NxVk5QEM6K/nIAU8UTBUK3ICRZw/8imGBsu25su6h6T2dcxiSQl5P6emuMZg
fGQ7qmJhgGllFO/l1izJUXiQHLjX4OWfI4JPYMukh+oGasNS8m/DhcwkcjWYtgIkz1lldZ9UufDA
kLJMidgs+hcImhHO/18gbP5UTBZN2u34fQ0nKP6NmZ5K6R6JgR4kLXtgKxGUIKnBhxB2EuXd58TE
w/gb38qq4Rgs2P9wQIe2h3/FfdXPtB+p6uKw6NRitZkVyZq7aXX6CtI2oQtS8+BzODVqNvEpGbkG
neK72KdAvgTPtz00zF7kBnA3x6ht6IxjPXuLVaWzTNElmdvS6ii/h8q371cW/Ci/TQwnz9Gr2PTb
qEdklyu5qT8U9ndnrGdTOZNMyLF9X2MI/AgpZqaUMLRW721b/KE9iLEnU4CW17NwYZw4lktnplDv
SWVali6EE9QgjonPJflRSsS5YLIUAnI3UZ5xB+OHTzY5tLO6cvJqSsI5M4XYsB0JY+JQJ3CeNz/A
V11dSQTlZ6sFZ/ERp56HdzTeQf5h3/4ZGE6Tt4IRgUzHC4/LlL/+wuW8HqlJLEmKr2fTjy2HIXwU
SVCPo/wzzodjznHXDpebhWvArgP5RfzJhKBzYluVx538dRu8OKotfYtGzMSadTjDqgoN/qU2X8vS
Bn5AeYhHvG2SUBrdk+RuU36/j72TUnueHDJRSbysQL8WExSUgRcOl8pcmhI8xX0193IVtKHXpHO7
Wasw3eP+Pem76aNh8KtoJM4QKCnjofsVQtxfINJ33gTCfFxP0yZoNMlfOqEuMJm8DndSqxKPlJpi
a/UnyUCHumVQhwrQxyc7yio8sK3MdD1XNdO0wKCvgOts3P30RZOxcuR01lXBUCdWogLTCW9vgEgu
zV4zqYK3poycZc5gaafWd2CIghx2lo5bT17kYkqe+95N/lSdHMHaCAj2qfeCebfbR+kTmzBWE399
8ER1sMo7V5YeaDANcHEg+mzhhDIIjFBMguPUUIweMS6evA9qiddHEg/BJIhm34NFWX5lWCNUzAFr
pXsBH7Ie5s4/KEPKUnlapuebus2vcGO7L0HBFNK3KPp7TEhAhw+kCFwUXUoMaVNlU+vPaoZ0r1tC
HxmQ79SB4K3Z2e4EWGwX5hYw3Rkpdf/YEDoRlePn49MwEu0AWtplLZzXuVXAw+DcbHR+acw9UOCY
x89YOdwk19AILPq52ZUSMmKK4iXSaGOkPmg/+gIrk7yZDPh9sGHFMHwkdQhoUoSOuQ3El7eSocIs
i7HR2PCmtFNgqEC52DjBsGOZtNSYETxGk93/nIn3/X2az7oxVs7Xd88d4zHXOrMxg9BfEobaMXeL
BU43p+CLhTyoGUXvkVVplr0vt7W7a38lSjCeYBijVeMXN0WUCrr3lJs/uGeMz2Bh6i48LPPSKcO2
r+m8wv+qVt+fLffNpyCLunl44F1yOLsGP0fX8TqnoQ8ReMS4gPDnboeTDdmr0KLVdZv42dZIsPm+
jsCpYxxIiJNUMiPT/jwn6wUQTtRFHQ6X63NBp5DsNzQQLQICwrkZVR+6EO03MoGLHr0+7QVnay/w
HPpczzQrWeObMn2jCB7GDamV0INgCchx9XbbfbN9rL5Z7pV+kr+fat1lyFOZRN4Jhz8EoUsWkuUG
35LeylJyw0DX02uwOJ5yU3CMxfXPUFiatc5+OygiAzi6zyBHwxjD4BgT7nxJYY7mQwkl7u8gmMCd
9/iRXezMJ9VhbfqkhiGo+n67wfZdo2e3CSzY5DktCXu3/hfE4o7EIhIumiaZcU5SmKlMMcmAop2L
EQYr+vB9Rpwacx9ACFU2xf0aXY0Cta9q2TojFX8aZ649AqlzSIYqRVbU8SJs/X2tfVSDjUDdQG4Q
PgSf5/DJgQo3Nz/kiPX7055KI8UI/XhS4PuHKS5PwQjaV+Fs539O/xPJUBzrmlHjQFcJ97h3K/yP
wcCWxj/urMvcnT6NUU9V2+IdVlal9neuMi5OXrcswsMWuO3yP5Wwia3H77VDno0FKs9anaShHC9d
+RDyvqi5djMmnPZC/eyqBfBhls5E5P7rXJMDzgGOzHy/mZLUiyikj7fCzZPbFrklwfcn0JsfVAUW
8fFWG6RQAO5tQGSBo2C/C4BhKUHjKNo5RlfRh1HeAwVVAxQIRr0kh1spaQDYIZ7EAZ8qnvvhQwSQ
mqlYqsXAz9k/TTXC2ijHzrvLKNlqTeeXYhrUIqh+0vuliGxOGNag4y19yetXSubcMpVSeDpl8L5z
irMlV53ZvOKo840P0KBsath4sFqYXNqc09pFNqBe2cYFK0upfrd/pjh+zktvHFseO8qWOJl+b6+y
kCaRd78hRVmgkRojPGrO0hP1W+7q2JQZRikTJbsYmzPrrECTioo9y+iNsgS/F6PpaR0KqwX+LRYP
ZUhwYE1HBNvUoIoyg/H4zj3pdBT/G1X9B0AHmDdkzcmuBvy3w7esh+vLMrg94WlLNmcC2eZz++Rq
vX4oFTDT1IGt0vP08qKs5ZxutctVH7n5g47UEeDR8E4K1lSxhuxB3NEDOZU4/h7FBVed4YBslkDh
10cRHm9jy3ivXakmUyoHZoWRExrvwZAdUCkSUFF0uTNsPWHuUiww1nQ6DFDLtZmx+9nyORllaXoh
CDhDpfP0kwiLU9/nR+XgTrgLt1YujrByNVIYpA8vtQomDh0HLq6ltcMZULeYJlFiOnLf6Ax1ksq2
y3igrjv7vBR10QBou3DMCzEs6vx24qiuc2HQMeTgPFVyrGgouOG2VjEPGBg6e5ZlT/GSIH04yLkY
67LQZfvO78Tu3OvQgee+CsJIuCd7z6xhGdHhDQWUQNJV9yDW0V2vxOubRujI2yKr9nPqBG4ZQK5R
/Ah4H1Qk5uQMad6q8G+KYMw8ENW7fzBiM+cOaHaMS6wS/gnpzFCwnFUVgwYZ5i39YrkT6q62LysK
ufnMqaMD3IWILpWyBzzWOUO40YeZCxo6UWFdpUitr7CAFj5rEKpGhZuUsvUWcmO7NmzYR1BCwWTn
qAgU76QJvuzDbNcWBMBwqLSYcUh+Fp3GgQMhXnl3PmLj4UsmROAGL6xEgWHRHzegL0sK5jhf+11W
4p7TX3Ity6wO1W53KDJagq1Xn5srtrb+gftZtKTxuyOPDU8ze3NeMmYXX3OYplMekQmExd38McL7
TWCgnF+dknGMd1r9UUQurqywAnXhiW1xLlwBTn9yWy/WLHvfOkRllye1K5aWhXKggMlytDDQftOi
AWETPjM1qaTTDoKMnwPAThEz3JTAYTIRxrzIKYbCc/vM/fuWDXXivFs/MALmx0qZKdYWXShJW6sh
40vfH8w3lk/MwRlgFMxjYH/Qp/Wq4LhbnHgFChPtFfrTft6Tnwmx4DZrKnwJmlR6R0g/0K1zh15l
LXT7FwoGosIx5ODNpfMK1ma/n4MjGGa8KU7TpAGykBBz7wyox2YXHpBts9RSbn4uTLA6rQrtOdUJ
NsHXOE+Jp4mhzOFNDjPtIt/sFtV07IhrvjE4yy/hds3cI91weeBFGC+rxNKOfjzjZ40DqMr2GN5+
qzeXc5AtXgXI1iF4OH5Nlgp1NtHv1MIIEXOoE+cP1h5jl71HpISHUa3cQrukgaCM1xaWSapmokU1
XLo4LhVv91BV6Rn/ju9y0axCvZxNftkiO79+fqFCdNqCdwFC4REf/q4HVUBN2D7kG+OJHotewaiA
+PjjHbCtATOsNt2pf3gMxmMRP5sSrZLe5KVCq8yb/uYsxpg8945EKpe2Z7n/1yTDiV4GoX1aBjvZ
WKHQbW9H11rQO3J20TK3Pa1EYXb7Duq6JGLUcbD2U3MOtuR76VqF+qny7T3VtKg7ovrjJmAc3E3U
Rb1nR9bDL8kxckXqzU0Sh1MExl4xk8zNSXAOy/NQ2cD6MH0T+nLqQK3oAkK4NbXPIz2l0jn+CfmP
b1MgWY/fUXGpLQy0ew2ac2RpKUDEhwVPWUx93+OlBqljXHcwGGuHGkAn3wm1ID+bqtVXEIeG4/6Q
AE9XIf3HpKmuzve7Y4SRYkHcWV1R7U5vWCkjiakDlEDYF3BVp4wegaYXp47xyRS6TcHFaDN4jvtF
KhXclPEz4XCl0FVM8s44calxcE2W2DRbSiAL2dsCqRT1x6Al/pC1ihzHgYToeo4mMkaSIMe+WJot
bjDA/+2rDTVb2thg3svHivCiSv98EiteFrCyi2+F72xAAbp11Z5t8ty4DWAxzzBGbgQKOYkeEyog
jWDk7y1aqP4O1emQOkC7uJyzPscxi8G2H0NHATzO+51gsh4ocFDdag4r54U+fU5NIEehBg+3b6v3
Q8CkeXBJ7CDm29TXPHvS18RYRFrUPTp+0l1Mq2RjRpXko85P5/RXGcOmIyK1Ywcikv6VoegScvKb
jbAXNlqKi1T/w3Yl9hRoNrf+fe/exerk+cTXakt24gt6QhE8cQYRPU6/qKB7w7+BcpuUCx4a3lAP
5qp83XNksbuiCPE1KgGuybPm1j5inr1d7zdovYPOIp32idDf9bEntZeejOJJBr/giO4f3tVhU5A9
Lo9esXEGvrIn7tF1mGVhBwEhbIBEe7V5XmXm4AdpZpPIiuvANtzbhUWDyU0+GZ8ksrEGEJS5WoFT
ihZbE6TrO1M/WKW4kItBAcwkbJlzmMzbm+VgZlXiChsVzCeobXpKpTYlrUbfkGqrhV8mINp1AVzB
E+/F/LJpwfWs+dlvM+he0xrTUvWf7FM1B/D57HX5KGGElvpBCNq6+yta1TD+8j693sg0slravBb5
rSn9oVA58Dbx6hCfEtUHKS/v/ravQAUdw88SUZSPPFj5kdD7j2qot1c0U7guTIcVPYoboxglMNHR
PY3WnhlXjtNqENJSko6GiMWUVWdJ0HnYyTl07VQnO3EYGs62Um12tesIlrSCgTIeytw2HJB9NGgu
71I+3TToimM84LCtlUgNyBU69832yImBUhPK9qFzV0IJMANjCoFzgZiYV/JNUNjJUEgsiLf5q53X
HWs8vcrUAzOAZAoILr/meMwHR3WxwiNMhpvHloahhk2stb6NTkcgERC0uzEzDyFCU7LsfehzD+z6
aGp8RfkCNyOe6KIOvnCuX8vJfENJ7x1czwTX6jz8NNE35xMdNeKDhdtFNRo0PUktJi9zWA0jsIWl
xKevnaJl6IRhIr+lkFcL1M6gq313k3o+Ia4FJed/BkqYPKsaaFXJtth1k0ZjruUHIbNQGIcBmRCv
AbiLO01mngNiV6dGdpeMtGnbJ3otuWSfrF3x1Ze4sBLQS6nZkNlBzbUtt41VnV6bxG0/Bx61+LpE
rvJaumLAXHLY4cncW0QjIo6QWKNzjSo5IYPiBbYu3PLL4Rjx1Ax8+29ezP79Y7DXFAnPrh7uHZYp
6lvKNveHz0sdtRJqJAsSGE4hpFqb5WPcODS8n4HvIUYSG3hoXA7gGSGEb9uDsoikVsHo+yOp6b5Y
BrJ6bo8qEwKTO9K9vfO3qDbWsLh+e2Hks4mamNCE/xVQHr3Evu9GP340bR04On6/aBPG7hRN4niR
9PjWqYq8eYLJGXSG2o/frLrHR0dezUNfQ9O5SHqDwHB+2Yt9TUzsA3V8/btD6guUJ8aFCa/SU6p9
OX0llw7B4FpmS7XGZ6lKtiQpw08SDhXeqNjqme9M/hHwRoSm+k8vT5VP8oEfgcCyhmhsuni/QGq+
dNLw23s/eaVAF9yNwlfxpyT/vRsGAE9/DJIHsnHpCwK9xYVKFpovgtAJ4T/KWHRNWtE75aCHPlOQ
EG3NCEsG+Dulq7TOXuLcojFshkyI/jZ3fMQXnIMWVmHGVZLFyOqh8rzrr57BA/tduGGvf8mdQB1G
Br5MWu+Adaj1pgCTnk4AyRhPp/AJIdUjDeXtfgKdbbyJRf1ivQPvH+fBRt0JVOq279jDbqEkokWD
MYUBrW0rIn2Q9tIOKre4A+886jy6kCJ8cPY2HBYtiHcgClOT2t8f9Y9MrIf25HJEFP96LYyvmYkj
+fxiAHqGhaHKMxmdIB0u9sBRXeargDgntNJtC4cEgfXpTRtYHX1xWsSNrQ7B1TmhGGDqNBCiSn79
k5zszvPpD31q337OUqZfHNyAoGbIT4mZuukqSczM0aeBPpY7wrNXWIICMUC/20aWdp967QDRJs/u
JS14Pg+iO3k4yxjShFjcO/JNc3XAGcG5Xb1iF5IUROXvPl6gS3bd3muJetCUn5x5y7OHms4EcoVb
7ABUrVOVnld2oPUNQy4YkbpkalqU2dQfz3007a90V6LYcPdywL4RYZuWKAZC2S04m5lfPW2Dsbsc
3lO5v9H/M/O8ss8ZGqvYci/DTP81MgxTSQxXr0ee1V49KJzJa2IdnSx/M6FGjTqRmEnuiF+ux6S5
Axfg0XSuBF1e/qO0gUQbl6tpE2wFrYJ3rMWJ6CSXqJlHvCN3EWyBR3jvZS55k0/d9YAU+5Ure1D3
F80FBTnXp31B1knyLrUnD8q4m1TUbGj3DqgZOWi1Hck79FGjY4p5uZ0Ix6cbeDBGlqaO5t0iKPq8
NqNGy8axEcsj4ZiAmB6ZiRjMculkjgXSOt9v5etjciRdG4GFTXPO/+zMsWbdH7QewOCqZo01Pwt3
HmMH/nPUriP2mxLki9qbkwgqd8hi6mledm3YFJWeVMp6jBA0vE+wMI/h+D3C4UEP3klDJ6UNUqNX
S4zNqWkqS9JHz05CgDX9f5yM2NPX+vBb8jJ21xbS0O6tP4akccVkihddq+4uPSsIKdvYyarh0KKa
0n1jZMLGa31v+iMzhVBnoNeGmCrfcThZp2HjVKBlLNvsWGwFOwaDIASe4KFyMXwo/b3vkq99B/6/
a0/SGGAmYlMV4rdG/AyWXQdJCJJTArF/BcrebFw06MpOueJXf9CkLKpMu8eI3oq73fr/SPtWv9t8
nre3HyA1uo54+SNxlH6sy2C9SdukaxysqBKibZ+/Kpd8VTW9Tu4DyMDtZFCMRV4ODNbiE37kMo2q
hnQdIzwbl1GXmNXU+CRUeKIFG5yWrZUdV+rfP7XbBYDo9I9lb1+i11f3vgfTIaIFEEAA0nI0Zms3
2dZx+CADeNiL0+Upa74dNgjQ5TZuJX6AI34c5ovbgb6GKrUiQrWI5P/FS9laXasR5aT9T2CXu43w
pg2Dw6Xc87GwdPMds/ZjW0sh3V25wKN0ZVYOC0GXljAT+gq0ZRzSS/EwKicY0iTMlaez5h35+28m
VQWkgHC16781tOxCUhzQD8Xy58Uhv5pBwUbFeNjBusV7JAq2fXNA0JVmU5KB4CwJ+VRhgiw1t+mG
9mhpfhpH6ebq6/Vfrg1h9dXfj6QGPquzewS7BwUijZ1c2SzSz1ohnU9wLJqzuzP9mNMRnhjedXuo
PA3EM2q2RkNQKXplh804x4fUUrJWvYadhiOBQ7IOEtKjY3rkEBBYtqduf7h9VR14NIkMhyoVWxth
stxJheWf9XDsb+OQvzz1HLBJJhyWngUJ7gQ+FQ8jd3HQMtOk4v2ZbFKJs20y+EDbjKygrVu24YhO
w0kmzk+Dy8GMTqnbaWFNTc+jl0AfmudcSSu/sEpea44qPJj6rzOkctn1i3djMNBTL/ZusLA4zDrW
e19Q4Xjf9DyZ84JTqvTPyPfwd8MiQk14nfKJV6Ypkst7XrIXv88LEmd7VzEwe8Eq1IKdwWAom88n
AOe99d8s9JsVh1AhUUiCjcOutrDSGhZDnvE2nKXC1pY62+qDhF/3bGOaaAT5k4oOjyLHBGXM6/gC
/DZuZp7xSEAGkvhj7IhhWh/Qe838zI/lhByA1H64CSml6zCotF0r1h4AUERb7X4494eJ/v4xHT/0
aZ3vejR2AbKBbjY9mxorg/ZN/XomEIVxYSBRqI5AUxDeiINf8G8EFwqTZJpKXT0SG4AqBIU+IR+5
H2ogYMJDj+yAiNmytIl6HvSgy/ytvCTaqgAqmajXahEKLwFEW1uSjR/FZhfhslNwSTcpAeTxkL9C
gEEFH9pXwmgejdAFTaOiLkhMWJ4DJtT8hf/TNk3bAccF/SWlpgGXPurKAMUvWQhG8kbg7tSwqHdD
oDfefha7/cmc48E+Tz5fm+/P+jHGwdEoQpxG4Nv99K7GLxKR5W8KYpYJA8PI423MqQ3SaP1tsRft
USCFKI/EQRLNuyBspqoh65T5TSn3U0fYNObxPuBvidm5hp83k7RFWmFpz0Q9qHGsFiJTlPGnjith
0nrwkJo+N1YDvIn91l91odxh3SFPVakEoPqNS7rtVEm9sodRhhFKuAFQhSU5IEvrHnTU2j0TqA3u
I1I/ZjW+SQloCRuEVmc5jP03NUEiht+fZIp+b8UJEEvkMGppyHyPQpRpqNX4ctZAFbJLes/Jp+rw
CdYfpk1p4kQuXOISn25BVdhhHxig82pv1e5lUdK0RkrCJxIwiWlEjyjbQLsztGgXQdlvcViHwuA1
pX0y3eE9ow575iVeOq0se5AvOj2OxbsfOBjKl/lpl97SI5YPI3I+hxabFCAaoh1hYJGX71jxycOQ
ZlIJdewfHZ0QAt4B+odEoPWKBZIMatqUo0x6LhXiflDVXMUyStVyDTqHnz4fYg42XVthADm6o6Fa
TQXlX4Wdvb+MLkAm7bfsLrBF1EuiHS0G81gWvJ5N1Jc8yhlbu9djwh11w2zlZVEj5mIFAKHWbKkP
cDw9xRxq3MAWbh9vSfaYQZQPJstlEtU6QaV+Z+7OX/bpbu4XF4U69km7llpd84MndTHdKAgmsW6W
ftjHvUPzUl2rg7twydCeHOZcpEi2yEdoxueyn6w/gG312L8tmjhNMrm0unTbhGNqTwUuQMx6mxxs
vwUJ7kAYLq6smCsyCNTPovOTOEz0OnrRZt8IoMyP6+Zhh9mEaPegH4m/XAqF+Yw/xCJ84R0HO4bj
4Ps7jWivFMfAbcdbfSBGMe1T1a2u4I9F9g++9yrXC1UqZO+/fcsRnxdSW/mYomZej8kDVJ9yr4FS
qCF32gGTZE6q2w4bZ04scKbOzjZaq1KHWmiLJoY7V+AwfqbG/sjZZzg7Acm08Obs67D4N0wuqL2A
gzupM3mxilExP+GRl4BuqGZBp+Le4/J9oa8KpFapikuY2ZqqLC5ocztymwdfbXOqC3LEMZJodjFx
YnKYE5v9vgG69WtMcZWalO2xMxHzC0mF7zU0TOdEu/X6PRIUsYZ7vTYKN6g528lcix5GPylZlezD
hx8bvceKmlRqdxtGY/HP5kMG30xUim0OSHK16e6QC+V2kZIOqYHlcmYhoDlTARgiwQbFl9Te4CBp
JuvqWzmxD8rbeMZbxE9a9fi0UMfKd9pij2wM/Yer32jdeAkEkTaEf5GGc8qv8y8X0sOkyoygkqEg
O8xnoyTo4CipX9rdTXvqiRfrk4lWUwLPn7+ccy+DYKbKT7Ywatqt72B8fbyHxiZQmE/tqT2HGTOW
RkubnaGHaPa5SdwFKOv3naI+f/WXQ/5IEAo5ZYWFhPN+Gx6Y9CHS4jy/S/VX468l2dDzIt3OfuDo
nnLwbmN/rLtEN68cxNLjBZGFba/SQE/0HcrFBANNZdzAfpSUJIbfb0ibTsfCY0Om6zeNazrKDXKT
eIVCqOepZxrbnvsdWqtZkbFvk+ZrqTv0Mwthm/sRvRZbN3LXgyKTkoFK8XoaOgAK2lvbqYNiN7bL
5I2rOf4JaNKdB/MpIJTlhRDoyflieCM7bg01VKjN3j6sU8ZDLpVk+qH3F/nMBunRJZFnvWpm1cgF
GZstwd2zr8kOXcxC/6yJrgnZoksBTNqJAShQE+3Z3bSyc+lsZu/9sPFIf/s7rlpdSrFaqsOfO9gn
JYEVBgQLYSgMJwZUPfifb94ScKyhjWeAp1D+5NlCwFWxo0znP0a4QwdH8BCCRQZe8Pq9gmxnSCCa
IyaFiLCW3Nd3y02Wp4N0R9x5xVpLDkfT333+hfBqYEWq9/WAUyVvfAT6HLg0LYuaP+G5Jk/d5Cbi
bKamtIPaonAd0rp1sZyQJHOFuHn8vf6KzGi8IQPFmhj6QZ5aygCVdHMVF3SfXWkgzZXq0goV1PCR
Dh5uCAjENt396Qr/XN8jxw25QrBvAdnq1zGQIy8yIv2dghYb6TToHaRi/R7cwKXNvTh5iGvmkiDB
Q2JxFNpM/5e3Cc7ZvhQOjeE5FtqLPeEfh54KJ15n5HBfbA7XwIObsF/tIxmkJImqyjZ+umUfVEY/
khuO+m3COJ+DGYYhg8YiX0xq/WL140NIH6ouIQ80vP3D8VrckwUszYoweZ2jnSlD6ixN8bIYX+wD
xU5Aws5zv2XE7TjSPKtxUMW1FosSrmLfW7Bwzlz1hJwJGSPZm/Trcwt4BE0OGd29mfC817klxrmJ
z+OGyCcGBR+CkBBlbwT/PkRQE6j4oeDh3QcoKW9PyUiG/5o/QaM0Vpibt+zSExzRi4EktnTtpMLF
YnP/cqlFwV5V//A3oVw9nrK6tcIpmWJaBWRU3vlBegwb9dRp7EDbIbdHUX4cJwrxaF9tdatONnxW
iH2q9YZ1N21VZ6DREokpzQtBAp9uUhZLqs+K/8cXacLb9D9anK/HZcszxTQBuwDnhr4eos6KFe+U
rRQdypAIHWb+nGL+T8XlTGWKeFwF1QaiI8k4hWrdQmZkrnZdCBkEvCeerTMIPBN61hP87bhTWwsO
46qGEeZMrCsNCv9W7aYmfbKg3sko/hQ1y504UkaV77g9+d3KriG7aIICJYkehtuHNpIbFWZXg3Ve
NTInzDqEhRsGuMUG7T83HNRxLx9UiLIssuKyg0gmUAGtO1jyZaGwEenia2cx7ofPy4Rw2fzsxs8c
dW0yOsXLUhUqsRO2AapDrN7aowj+OpThKHNSh47D1x2H8K70PBg6Fl9fFhLiM71NxMMerSXBJgKq
HmHvIWWmRM7NOpEEVBw54O+9R/1XpsNSeUX7HbTkYdFckgyMqDwQj5nJMby7jLusK+NrgAgGSajg
AMzipVquq3dWhuODXYZsrKGSG/A19J3PdVOAaboWlb7lMxt86AS4mtnAV/6p0B8CNvVjnfX0C+j+
XvhjoF9WPXOO1Uny5zdOPAybfdtzaSvBvNXq6g4Sg8tlJRHLdRhUHL5MIcY24LbCkg/U4tYEjZYh
aiLZkVVZ6iGXD0fZ3SrhTQtJt98A6SwYsprqB3tqUMe2N4zL9IKaSEM2bw8aCqjWx3cUg1UgKbvu
C/TcgJXEhfMr1hUkGDlaec0cFfd3PRcYYIO7C+7Z5yP0K+EWseqOZEodX2kp1ZV1mtwdKl6VkQ3k
EQY0Zx8szn/60O14wkU28x5T1YktBBVS7rZUfG2KQJz/wYG8NG1BkmaNNUPnUtYe4ROwp9m/yGT8
hsVpT07jOfSRv8fAcDD9rSKFyt6yzgcMo24I+U8wjSWXLPucSC92zi/V2UCfNQNMPdsJb0ycgXzo
T0vSdJZeF+jmCcQTrPig1DQJmk1coKcslGROBJUL02C7kDXGHikMx4IX37036cGZfYR0P49qPo04
9yrcee4AOQpILx0PPtdH808+ZrjaDruo5afcs7DxR424lt1DqR5K95RgAnteRG38ztPRI1jOHYFb
bVBvsbQmLEKCGnSZ7AhJ3Tp4ItOhPEnWupGj7n8bKkrTzopoYu8GaB9o11lI6XYLtDem0kZh8DwA
SIIZh315UKEqJJYI1bLOANDe98tiTuyG04b9IG81evsTOTg80zgYIVMauhCpMxBqcOabbas+9AiI
Ghi1pSyfQRkedPSuGDcwPUdSqnM3QT9zRPGj4SMVuQXmklHUuTifJWQeCmIbaWZg1RrpdPfk/QUQ
hgFuGrQLdNR3cBeqZwenlFIBHwnri5gg8EVhfyrvNmhgQqzcBGrDMnM1822ClcWJKWikdbt8KXcV
caBljA+vTESC6Qa2BMX9wKhhyNYbLkY+O7An4pjYwN0a/5z1WQ4fv8OSZCZtbZflIeRQ/Ql5blZR
QfSA2QUXnyoituEqPAExd/nN+j3yJxhUi/8A9xInZKyOyHgoUqsOyVQGiBj/pwfchBGGA7jv6vOc
vtreR7Lx6pLHpu4qK21er+DiPbKbEUbr86RmDWRwdz91mEMfh7yiyij9HHhz0ZcX0r8E8Kq512so
VeItF/qR7BoAEZ4vUiCdsS52gF9xUEvj3PqYmvMfOD5YsLVGxdTuiDZAlvxSyaQjgkl1BEw0VuIz
af1ntB3OhNRgfk1HleT63fz0g+EmPc9H1ZBFB45X++HewxNkY+kwX2JAfMA4fxacnLtBR2iLcqkf
ntO747IfUX7oyw7nsrN3/M8L3wb7UZlOuyBXtMre/kiUvgoKLW1489h5SG4SIYQgG/mXNZkUjklV
N4ctLkQ5GdVksVgYbCoxqo2EzSszsy4+VAcHrptxkiQbFjesei0PxFuIW/kVmi5fCnH02GvAgrM6
+Mqpx3CAU42BMCcQQ9NlSrIdZyOihpGSdtKlhwU99y2TQ1TDl2GD4hAWFpBU3nF8pWpnItaZhxjj
smooyzFT0Py4Htw2KaT3uLsO7FQ9dyO+c4CsTzXSM1u/LAeE0FCkZO9PCpW0f4mXCHXqHuInhcY1
XRvUNHlpBNS8KU6mF/QdS2oXN6E5tlzovNO+7tPKyMP0AhfHru9/k7deMOUZwEfWZDTif387rJ+d
HPg5xtRIXC+lkkdJpBzm8adt5xlSDftxzZSaTvnBSgsv8ieLn4qD5TSB0ISfYYL/6vtv1jJtrx4f
y36vJer3HOJXcbY7DK+T3X9fgv+l5SdvIkrKhXmpn5/kG9VSqeLqZob38CTNLIh7NCBrj5oNskgv
lqa4YbgEZRWITyTUh1EA3Z1lIqBqMTuD8McL/JQ2G1cLory5At2QCZ0tw9DeXcPk0xGWCb+ZmIZe
ioN0UaYYCcBrzZvVDEi3+cHYN50gh5FLjsxoicWIQ4DdJqjJeQ4Le7/VznTG+HKS2K1/Z1PpGxdk
zbPHFzdqmzKW+Ke9PQH99EuZoBH9VA20moFF13lwDAYVw/gZJu+8CmZZDqLoV00akACFw9w10tfk
IkWG2jZl61aBytrNA8adN3MSsCTqlzwmCx5osx/IyHiMLit4s66DX9e/givRqCmEsXt6F9t6KNS5
eVmcDGSY6cMEHPEVnbGKQ8muSizUo2bpUHX5Jg+jBPsUnEoc0uXPVrF32yKzQSxUTffrVo+/kYOj
fkRHK4rDtVkdEcP6JO6zypRoANNk77Qg7CDfI368jWsBs/4yv94siezb9hjRW2Gq37epSoTLUhNk
cr2naTZb8vnCvLt0WId89Py/ZcAoe7grY3kNhQxJ2q9xeudF/rXPDK3MOtPuckjybEZYPm94kbpU
W/jAvn0IFuPxCdLCgawc3T014NaiLaTApnExeyNUuB+yFaSzKEzuPz2OdWSXbYjkajqcGoqf3lGK
jRJXjH3KAdU3AxeK3qo22VW2S19w07dOxtXzbNi4LHe9bljMDEhOEbkPpcrkdeuoI52IrYji+jyK
+ciOBuAM72IQdFCxC0BruWnw+uS51ExTQJLBZ31jR/8jOs/SH0fgg/Xtz/vxjHMHrLCDnNJlwYaM
pbCs3wHddmLNC6PHSNZ8uH2e8uKSto6GoP+88CWKKou/BwmmRCMICaViOcH0mvsPY6PjAcBZLBkj
7TN0ji8ek7+zWmG+/1R8YDS/ayah5G8ExxgrItGPbqyRzgkcciy8QHRL2R7l0vfwT+CvUlHJ8bda
SxlfLtSEYB1D8UEQdoXTIww+/eKYgh9lwgqgEJHA4dlnsX3K6O9o/4aHWLU0L/iKR1ktrE+mVeMx
ZBwSQeJA2/np29JeG78zvZMEJ9BBaPU1nYfMuV0dYMA6xsl7LQl2yJXUcS309edZpv+/7O3m7kdE
xrR3s1tGNKqQEMI1bCY49MnKD/XoGp0Xn3+mg0HSmGTKFk1QHyelJQUjbAL3/axifDPlg5y1wbl+
TLALoiriefNybFwzBYv9TR0TtaOD84ojw3ZP89A5XOpWnkZwSY6091nI8AcMfUXC7K4hsiMWt6hK
aQ22fZhv5dtz6UMSw9SItjO27GdmAeAdInMYxXzXrDvk0wkpH8mhCCGSenF9n/p2wUe/6I0uxRMD
zs1K2xudCiDBKeilqmZYjmLvR+qbP7UChIfBD+k/uYJfypens3wR5qH7fWyVOPXdtHIlQWZclc5g
iSpzhCLVF9xjcYGtUHjqL6rGel05Csdr8yFVq0VDtG0DdXoslP3wYz/dcN0UwTwJspCADk0ptTd9
gkg9gIzt2Qp6oigV1nQz+lEfme/XnxWtSQK0c8wDKZw2v6hZmPe5UJYdHEINYpJ0fl/Zk3gR8vzt
Vw1thhu6MLLsT3TdfmY5ANRoen1ZDCTUwmLWLtxQI8xAbI8GJWyfYz72EdJr3G7iOMlXE5DB5JAT
3YC70Rz5Ag9nyOFl7TS4saalKJonyV2uHy25ETCEZi8fY65YPz3xBD/hNnDbZo/ULkM35WTuN7+o
YOjqDH8JT97fN/OdwR+DSb1Flqzl1cly1ld7AHCE06y66k543vj/DH1oGnDoiZvdYlAUrvMZT4uX
meOjFVcASBDm5qyLOzs8eOo91Kj4Z98n7T2m4akC1mZYMFHMbQr1vp3q/3HU9cfs7wyaH4/8wIGn
tRSnW0adh+acFqyaqQ9vlWJIwBOxYUFuOhR0LClXtbFZunB/VVy5NVWm/EjAUM11zTR3z7mabSnU
Hq/rZPYTRx+oiul/FjcuCBCdrogVypgo9Pq6dbWab1svzLo6U6p6yNKyW/hBmeCaDsTavQqSbEAa
QUMsGoqlKr33gKPu4qEdvDDOp7P5rRNSbXU2Djknzi+f7sTCQKyxRYQEOrLEoFK7BgQilWNU8xRz
QZGvuBJPJrXnh8rE2vOC0GTKRvN/9ZLh4vVSz2jm/3CasLForUvyP3skdhkN5fLrtDoFM4W3TXc7
j5s5FfPGxL/+FSVyoCQkFP+jNBfjJe9/YGBDOzQ1M81BvQl0b+Z4ZG7LgevInbsMXKlhedv6qHAE
1/sHXR3Nk4xLRl5mwsTYOs5N61XCxTqM7NsnCM7sEA4bfKs4IPzUAeizH2Tq2Xj+QBDSp/ODnvt1
797nfVF2nk582ln5IUXOiYQExr7fQwYWAuIXr2YOSaHQH66OhAiZTn1GFU5pXZ6CVsaLOvLhc/a2
Cq4TznxC4yFucwXtAcUZ1P2cfhuFZT8ZcRMfy09RBuoOrTTN9uwpKzCzz9I8pb2cFLNFxaCqtyZ2
dleknbelDM+95j0ZTxT3kHWzoJrOJfGexwh70U3eJTwmS0Jp2LRJ1fPJKi7jCHolWK5jBm8GQpnT
KAQsAWN7K1P3dxyFevkj6DEAGSktX4CNitw9NLcdZPhei6lVOL8Q7dxTuIOHlN/I7kSIAsdtk8zi
0emt7EiEACBXe0RR6NnIM9S6Kawa50M4eN5m0/GITxc0ALHajyfrHU8WoDEiFH2EvtYOijiPmPo6
L4+R4rxR1AJn4rnzgYgRtHeVSa+hWc26lvnj7DwkrX0zAHqdEbYQitvBAW/GGQpUXH+MHOO5iAIU
IH1XFiiyY48cUf+f8xdwG5tK4fdKkClG1DUbEiNmF1pAQR9redfu9MUPVQjxIQr9FWzCk6uXT2/r
2W+sNqCzxRmsYO/XnzLivw+cINSHF4sP/rJTnudFPF2Ug/SGHuTpZ5p3Pzo8gp4w0atTjTF7q34j
6mdn3zSDOGMsPYiE3UOr/rIeLp7i0k20ZUcJkQJ3/Jibjp/fHL2BoAuM8TlFjDQnqZW3FDZRZ1F3
27htVq+0dcrqGOL942eNKooQOnLfZyB+3WwdkB31JW3IxyzUUWRnnkBB7LmZTmTWiDny7Qv5myks
k8f9v/0qXtJApYYl2dbek4k1+m7aqiSASXHrqHMPGXB7V+5/KMVKDs3dDGZU3j9KMuT0Mp1KvaXp
ZtrDSuqH55EE0dppwJSf5zAevJn+UnmWgjNXBLoIZYiMBwi9NcQacjsmiZLIKPvEaGiZbZOP4PPu
sz3wECxLuzZjszj11BUO5n3g/5xX5Pq3hKrP4gQ3vcnj2PFvHY/6FEWzcnSKoUZWTEmZTBr5MCBI
TXVytG5OcLrUB1dzNBcP52RZzE2sS3uqwzuhiGzvLGExLiNB2tlSDqtfP/1B7iSIaTgmVqB8NAra
5XUuK/HoT+/geRR+GGqhB5dHi5uih7G7VazRHNo2qdYOuokHLuxMnptOl8BJdQHpRnkhAeHw0gJu
6xJABY1n+OKIiWheUW/aj1Vp3Lz0uYeU4fji87ks/cEjeXHgGWFoc1UEQyfcYCuGDLkMyNEElgrw
cfgvdBQPlykxZT/koLdLpN9bx6NHRz6xo7i82R8UREJ9cNONDRUWI6MOfDRt7yozqSD2a1VQvlTV
OnEt2jaYC3dx4jv3twpJ0xv++oclbcklx7VyV6LiopOwt1kiSVEQSHb6EN/5/hMaNvUUUO3L9gz+
S0zlaUy94QJBmDneT6GZCJxWWm/qBaSC9869vQNW7Kb5Znwf7NKDVVlH/Dd8yFtnD0f2Ln3GpBrR
W+16Smm6L144d8dfV7sfKFPBCgEczFde6DPCQf8AsdOEjYHCHH/QIeKNOH+2wRvxAo+FhLjRJ0ES
0WHv5jOSXbaccs25DP6I3nkIol9tybwYHzOh3+BE3RTl+hjYJia9dqYe/0XqJ/2Lw4meJvl0JquP
Sw5vDcKt0TFdg6voroXLHPhlkFWLEkOd4nomnSTu8vM38Ihq4oOIwYQm+y9zD5d+4VSB59s5AdFU
gE/MWyZBMoVAp2JzSRrd7IUKsSOQzz2Dm8oK+5Dry2BwAi/ftOIGoHcSCHH2o/0RloxEW8SMCHkp
YijuOdJXPwX8kGeXrvept7/4vAlh5tim7vaftb44WNlDVtGmP5LZktGlSBuyFYRhw9p3vf7ljxRL
2wR44BPV6DesEWyTLHBZ3a+O2QPsslgEeoYsR9WrZdaHmW1B3AWRasCaID5pqNP94E83aioRkzVw
IDP5TUKogB94B5RUHpB3Xos0k3AOHuwD/C8ztkTI85d+5ak8Np/FmhOziiV/ePyP3T1ytZg6Menz
F6Y2DoPikes5XqkiavKveGiC/N0wit2+qoT3BovZth+p4UiJLjb9tOgfsE1uJzNcLx75Q6f7wHmr
Fs0Y20his8Pw6CNBoWLT+MPcgsbCN0/74yw2ssf23OYYd4OrzT07sqKKv5NBbxFeQExxOxPkqFaD
akhrji7Yd7An3HvxCmG4ZHBv2GyQYVA6TChiwRPEe5REk0kpEGCRB8BkucYY1fv7X6sZtt75pwgn
KwyMNcL7LreLzQ2vtNtJI1qjbI3kacDHbIB86sKuQPvgXQw7bt4Y0Ejl8E6Ct28+M/Pf0nWt9qTv
s+yLLq/1lIrWc6AqY/NNKxV4rVNsThBKKXfZlmHTR7VSojEhj+uAmhNedix/qzJCnC5Cta7bHmMO
hXkrN9kyUyigpZloQWoesvlDhTaBgeXgbjDu0+4iuPVjHGsnisclkZ+qQQ4VdgGU7rOVU3rak5iR
UEl38msTLc1Fig0fvKAhGJnn5EyJse4xiFPXCIoO+FVvA8RfU58gzJ3ZQ50TUiFQy6iswFhFd7W9
uPQ0ThyzCRj5kS1E96fVFkA/QWC4GHQpwJtAnc6S+X3uABK06QumFo5krtdV/wcMJfPnIvDsoeTK
gIteV+aYAcYythBVP7DPbS5oHkUTg/jwbeeYtzpYNSPWiIxZNZoZEVccRPqewsoG/bWpR4ykY+XK
kYMl0EHBBnXH8mM6MGVhO1W/gFdjHpufx1CqtJFYi89oA49GVvy58ComfP5AZEG/1x9YMdtfqRUh
cFzV9HbY6TdOHNVedrYwhipOLP6/oe0j0QwveaZ3w6L3DD2rChxoTed2V7MMncEyK5H/NFeBSLTJ
UZACUnbH/kexe8HgO1GB/oL/SPlr2BabrBt7nOyyRLbgT12gM3lW+k380IZSSbhG+otxeZYKUHVE
tSrR89dkNXYPSWbJKqAV23GgIa2jf+W7ODB4cvGupnBdfhWlti/ERm5GGVRM19p/PqZnFiyLvoq7
waddNtONJfCV7eAxcvIJ9/yKp7crDxw8xgD/IBEbSGDamJZPnWQPGcdvHat53w4RKpYP4+mllqyn
k8NJuXWj79iJ5qOWWoVKj16QVhCCp4mZXKOtYVMcLN0DET1oG/N6yQCWJbdoBNwvSW7mc0l3bQYq
LTI+9n97VrmSOgEdNUozf+TN6N/n7lBU93yRnhMGHCdzzIb9ZCzkjamHCDC8oQhdf2gWW36h3M6y
0i+6Bq2k403RIGdeTHEG7d7IARaNXSklL7Jpgwb/b8aa3pzfgzPbEtCFSm8Pdsw9EP/1pplbhIgG
OgDXzCYbI/vwe+vgUb/f5EAWV3hCLPrL9i4R7jO2Xb+Svxi8yd4MYFWjMFdvmBI8ZGMaZbEc+Qto
XCjrlHodjAIOuFSs3+ilchMYKf6YPvJpcc6zF10JSIVmIo/2GB7S90E5CF9RzhLImicVObUY3Zns
hDoVawynqZAAPeovJZSaDgbYrRcx5D2Ujk1mI+ENlmGvgLTKVlAil/9M1ju6MnQJHPOerD6ZJ3v3
1g4QYKVk8bJwEvgyHLcnv1DBcW5DOKC+frVkmwyUYiBxnQIsOnRtNZOCoXUsb3uHF1IkuiYur+k+
xxNT7eXRiHWPcrKlRUiNZlycTip7BWtwi+/fLfYqw+dmCKhpeAeckyCjSfWnXtaEzhOWuYe8dc23
ktk9y8lezcs/DyOeUJfm1cAe4EXO6gSBtdchB5SX7ayfwckyni7qMUxQDZH074/ZobaThDCoKu/L
3bkXDyv1eDOfxsrXG2FuFQtAiPKbUBvm/hVcUjGsOhuDdh1eV6bG2U2UnmbrV5debMpMD0/sfI44
gL/CIKlqP6e5DkgOA+E3+FtGerFF5mSjljeT3YYTSieizlx/oYP3s0nfbC1FZhPkmUQB8KX+79pH
wH3tX2c/5dPBf3y0Nw8ykHhDbmEEmXxlS6gom2VIzi2tLYuReImDT9RQ4zhnv6Hqhjx39cnmcw5U
olDGv6Z3tJFAsfHePWr191l3cVxl2Ztr02s4/Q5CLeuZ1R5vQIg8K/1/xJWx/onjNXcYZogjnM/E
lC3qd0VK/kX/bnLpupwoWm9f6atQI8pgLYhns1k5RCxWIOjeTjnuYnIQgxr+eZJgoBOdE5U1VrEV
H1QwYBUvbnEL640U9StqBbU6NyKPY1IQ4yAARa8eTtEzO8i3co/4qvoDaE3teA4LTp1YQaYKXG5y
eZdu9xXgJi4tH3bl+MmofBtf7am3lusEaiMCKX7KO3x7v30bEfzpZMT49MXe2qnNervU32Z0jmvY
I3ofnYBBZruhquM7OXqunV0TlVH5uvFJZR3q73+QpSY8gxzonryh7hNI1zLgsvHmTc4IETis1NUt
EzU/0xZZcMzExN06xIuT8fjk3LtlIXibaStIM7Iu8OqOXSjLfFvA9r6KBzBIdQ/bW5FRwSPPi2BY
zAqJe0YrkBi77r4s3o3Nj/SJMAmY9r+DLK/hDlvsPV1d8sHrJtLDrGWlv9tHY+nTzLIlwFMQ+WnF
1HAappP1n2oX+fMkhrBVltGxfXRvFzxwH63V+1Oo4fdOe9hsMVEWEzHn4744d0tzwE+cyIM9I0SH
NOHgLzAUKEr0OV+oKMRdCWTzYYMBsvWqAC5hjBnal3JOZfkJkX31p1ALTtUiWrWC+ukwRL5A3a/B
o5Rt/25dnrOGRUotRYp9TMoVYMtpYM8vj5DP8VD9A3GGrTrYZTEF2TJGoiUsIvXmEQNdna+LXzjE
2qlQ/E0JEv5IQvDmDmP3r7F1o+WEBveRyBelnmrbLZ9C2XeYAoTxxfJqTyxFiGctbPw37UsnFmhP
Tg/6H7KAQlfmalEnTMyVHFjtIa0k0i6DdH46D6y4wFNtXvCx33TAbaC6MOYInV/jW2OEXjdNYQ1S
C007ROxjJSSgfLqRHeI5xzt5qOrfucgNyJFXugM/e1X/SeRT6jICbd1ZPN2UwfaR1VdIJzvDCJw2
GFEowBpFdDAYcH7LI2nT/LZHpJIxt/oKealgZ+Y7fcKkkBC3dEq/wchjGTtbvFPstF+SLxrqIFaC
RXFy2ck9Hod5K4Pb2rKYse8vIktOJcP2veBfIXD7ju8m1MEU/QKL5tEXCi411bL6Y2Fw/aZr0Z5f
C4qn8OZsY+XTX2AKmb7vtFJ7GitVjdy/PEkcgKpab6K2IiBwdYQMwj0hAigjk4uv0JXOJRfu7ilO
eMrH5T6TzQwQ5WR/GzEe12jLmCMkzUQPRKumWFLz/eDmjQXVhiaC6zE9aMMKJDuzhle8aWLueVp4
HFUKi6YolS2NiN5d4O5P9naUmfUJ3AMB0MnGgJD70CPZKmwDjDIjWxbAkFbUe+FWp+ZSvxLV3VDG
OpD+p5sdWNNKQN8MXNK2+mBDNWM/pyKFwP4HGge7C1fIXsRd8gFWOE7WYIdJV80VZMzeOaPbbHmk
fL2CiL1YDtJvXgdz65G69Xn4jyfEbNuarX/3g1VQh4tXt4XqXd6jo70pHcXRfrxSZKVt/LDFWBNF
yoFM5QfZiuTUwJVXVJYC2zG62mivztZ/W+3NkATavZ03PmssBd7tDLU8Qd9y43VpL8BFYvZ5fdwN
PhDjsZ+OU4ALo7iYn5AwYQ9o9oI/bWdVqQLGE/A4iSBKLZB8dPYWZ1q5uBnc6d8tqaafbj1z9GML
9n6m06CUHeeC/RocGZlE13A0oKGhco9pm0VJzR5msY71z5GULfqTQbk+3bL8ebNtzHeswKP+Qqs2
K+uEaNcFBny7btQADyBp6WupBT0p0R13AWsIbGHobHYbms2ML3QEgKB1HAgIZ37ViYNkxU2vtUPr
iVQUpq1ifmdBNeXBROHOoQVG+GOPnSTuBnsiZef13QIddtQUowNHsPhyLu53mjW2Yt+PJVd1bDt5
0y0No5YkFNXSTBU+nUUuC1GFAO3u2dtL2LdJLj2CEIkVG0zqStY1fqlbi4hVn/hfQXzegDrmvQAG
GVm8bGhuNUogCJhcx7jTlh+l+dwqHuRJ2NTr7L7AZ/Il74uBZuT7bdo/yHPrOquLF8VHQP7vg+JK
eDOVizfYwuyzFysdHsvMaM7EQGli4VhlWBnjB+3adBns7IAZzBdpaelAO95NtioM7n24lQSO4f1m
rLHxJYFxH/9GpFx3LnXfO9hbmFCFw7RAWWVBZqvZXIoqnnceU3LD9Hk7LqK6GRedYropMqvQvnBd
r+kHIj3hbxzgtH+RqPGmB5vd9FNUoIeRAu36HvI2YANqyo+3FnA0UKhd36mcvLsLBsMmQJ15vbG8
xqWzz7wTPlxUy6Ot9gSKmvKiM6x3xEA4D+3zpmGVgef52Kx+9G5L459bQihDXro3otPMmo88kyM9
CLl1qjsqKTFJ/27wvvLqhnmLi/3zl7dcJBecX7eCouYNjTYvWlpiaTlmXqPpK6pV5Cwm7rPSQ1lB
KRz1YO93IE5TyjTyGTdHQRp4C6PN48YRJ1v4VnxVV7rRVQMR95Mu0Q3iPCaWxtSnwNtmHf5Q6SqQ
Aj7IGyjz+WQV6zbsxFM4d5x4ZN0HIh2o1gMuM5N13AZ8oGwBaaHdSzoG8XFad3xOExbZLPEXxUga
iNB2nUw3ityEeY770OTUzSo14kkMZKuqbMTyotZsKU48bBQs2fDomJpNmgBwLyeYFWoTfl0Sb14/
kYKLp68JAWy55hCwGGvSSssQwjnMoIxO7m2f8VxBLPJaUbNOuHFAjRNGmzmUFhY4R1Uki8E5fIDv
LJQb6PBcw4Bl05lV06tj0gcPwz5GzCZl1RRqmMtmfH8GohEFCSH08f5TGBRAhNiKsFYwKV5mTa0T
Tz5h/2hxdGg2fuInJtKcRi2xRqNtn+eyhG8SOG1lwIl0sl2Xri4itSmwO9ZKo9fnf2EfcfAqWGmD
7S1YwSj2tAwl3ya411j6YQnIyz7HdbXWDkkzT8uiG9gmcmK7neShWmV+UTfIA7Hz2yzF1lih21nd
Q55j2F5HXwppbuBZVQxj4iHhk/jkcQ19WgZOokqh/qfsTvyfzpzo0p1DEcBrAt0ymGvKq099RZfa
ZKqAfHfNv5a3OvlqUwrqUKu/tUUK7RdelghMXyJfhPqT2DP7pUpop2k0sTegaJ6EU2ATKNn3qyPk
yME7p0PC1pEUryX3fX7mm8B1KW16KGbiXOnm7lOFm4oZdgHTVZk0cL8IWdmzsGCdu9Z7Ch3Jvyfm
OLoKE/AylbHAZaDbByEUb5ZH8HFNebmbogtRTB0D8EnMNUZ9hjPm5NWhqdpazQquRoEXV7CrLXUu
iDKF3sguOaRCKqiVpfTP0K7jWQ4Q6llbJ//trAb+xB/JzRPc+WARRZJxWuy1w3l1r4SdQSNzw1cw
xUdtJgpeKvGtDqFCxsXGLjzeSPP56zj1P8xnBfjPhq7d4Z63ue7DAK6r3w4YpcFd/EWj1GUZBxLy
GGaJHoSBNo5uHbRVhdKjfmxjbWsbj1hlLdOd6V41Rai1Bq+Xk/hcU94p3lPjOnbMrLXavuwMvkJn
zaYLcuV3LHn8/G+1XkwochAEqrJFe4Q9w2M/GpwbNmnrFW8Q1EJnkvOyE3+a3BB+MGKqd4kIz5FQ
9d7B9VIy9jR86aq1MH/99tTTn4UJFP0FrjbxDHlUyaRphC6AzIQfVa9L9wDRyARZaast5W2N/bZq
AFBy3AH6CqGYYpDJdOBOIVOCY6n2y15Vmw+RmuQ/OMgLzllQ6hPVYyW7/XMSGnrA4g+AGcAnOaI5
2h3LY67Lx7DkegqZ/hYjM626HxMsGzFq1z4u5Mj2gR/NQ5S516sQ5Jeua2g8QjCnTvR0xF2sG9BV
TUbsHsHwT6mpiM/TDpRTmUl917kDHTYyZflh+lX+j1FV0ObM2jLEx2OUYNf5omK46cqOMzeR/lpV
+V9KpOzyQTSzm9S7HndElDIeshcmqZFt3x/S9EYm4jTTNJiMha+naWVIF7iEjYF950uyNtpBaALw
igYa+64+IqFiFZQ9iuPyfo/mqAbqliCjK6sv6XVGE/1wvLRTzJIGewn919yWHcYUC4N25jSQw2ey
+Jlvl6W3S7Tnr/XOrhyl/EAFAx39/o8XndoQ3/sAjNNlUjXAoPNFVoJYRtv+95M6vLYm/tVtKhuV
FT8/Qbd0FSPJ+dF3QFfUWNKF5JogIpx2coo9TS55w9xKXrhUy/wOmkRvlHLXAuuTjOoA/V389HYz
hvrEl4Swr7ofL34bS6MKG5dSsxn8XOAzlHEcgSENRqxrTzlq/c2AB/LxEH274hJjbaxeXE9TLjDd
z/5d3xvsJrIa6eq3ZkBxXztNTWpJfj/zOzjDKYfKmqfH97jRJMI+ZqOk7n63Sv4/gMo74y8hkL9g
1QClMEpB3PEh9XLBTeMjl/gv5kVsGKdQ0GCbCDt/9F/fGK1P6XA0WZTfffwliuSCHGC8Nxgd+Ni7
Q4uZBTPEkEDXcvLEv4h+y5fWVsMbt/ymie53vEklPApa/tz9uasMjGjMR6YKMWSYzrCA7z9A5Mxn
ED4M8z9ux0uncFYncuwVjS20+IFbImkc1Q7ew76SG1kT4wxAmXEw9wYjWUidlFnJGV160HGkB0Kg
FzmFF8DdHSHriJIalcB3YpVmJCWXJGmF3jZZrjgK2Kkv9d9AUMpea4PGEhD1lMl7c8y4Ni3bbs/v
7TxVQKUqGwO/pYkiwCcMxbjaimmCamFxTorbpUmCdFxCcfUWbigQ3js5t0Xru+u6FZbyLjqTmWmJ
cZ2LIySytum1J0RsleMEu2rmYe7zwDpuOs9YVUiojfyAfUs9Ly3bCYULZAZx8ck2yG78ZqRtGK7a
FhEHodyazj/oDZedQLQ2k6p6w7kQTpMMFU3ArE+HuYk0qzkAhF9X7hx9yyDvTUEKAmAsotXpu2nm
+jcdKJHOBwG6K7/vo6FJa6UqB+P+Oc9E1imJsMM+gDUhW9qfGHmvpTH5PUXkteoKfzp+y+aBKwZJ
5uFH8uVxfomtW6oIZepuSvbF436jXkegC66GtN+blfa9hCRBl+RCTm1qxkT+jrMeIE9SkFNxc3OM
Jsro0dM7Ngvj9vJ6ex/1BKq8ndMbhlLt1VnvvjafWEV7gmjhWXkKJ/QLsCwpWil9bXzVe0q58gTt
/xGlQzmsU7hwYI+jZhxX3H9pch0RyID+2Eh75TBM+b2VXOdtYJElALzPajQxOrcpREJYizoJN6Xi
kQnQUmLmAeLUrQm+ap1mv0Zup2jVhevR9a4ZULn/A3De8YZgRtc8ph8qYefiBHU3muMnCZYEzzqP
jVNbEpRFRmZXyLoJlLIjAeTep7VIvZK32HrJ28FHXoiyCx8o5hbxyawVv5/XxY2moO7plapvv5GR
lj7uhu0+mwG3plFJ7vL9qL1bAibnZ5yB5n38XSKhnaq52VAAnE9kru3wC/9vnzP5rl8lXopQs99H
lpuSn9o+XJCC+sVgSnR+OC2InWrp6jeVnWw2jYY0iWn8dTXo9PJL85xdwBOfAsFzxm/o3Q4VgCV0
p4qRF0q9qtYyBsrobuma6Pw7w9nCY3BUn5Rp4fGjoRu4gAzPr74vSa4s/q6IcaoaGMMvqe2aRWHy
/sCYYnyThfzxVmYUjS5k7dfSsFDsQTGFkBk5MANcFlUTOltI9nEEKKjf8aUlx6Fv7RFwOgKjb13t
PJ/uLxOamKKuixtirSc1aNdQ17ssV5UARtmF6h6FPpZjfutYc/E8t5+TPFYY0YdwlLyL24xkBiVg
9flY0rwNZCRzrWsIOszUZeyoiIc+AymrP6hZzF54z7xRX76h2wVldZJT9axxzO7vsi5/fd8xZqlC
4RPfSIBuETPsVNZ4AK4dcZkqskXYicny8tlUBoRcoCk022ns+57RL39lcY00xVcXQPRvgwNoCIPf
OPmrFgqwA8osNEuKigCQW269XFLEl5VIsWiTBukpyNgGT8DLiVex9/XjTIQWmfWPELnR3wHW2nMM
YhEGzNMFoyLTLKXkkzCfhaMg4OfBD5oI2FaXuVfCo6SnH8oUv3WRPzuxQ96tvTnpUbIrXluA11zN
YxIF1PwNmhh1Ju7Y+Z6U6gg+aOLH+fbTWN4yar9dHMbLyCsQe6mi7Fh25ZdRsuBEQDRGKKYKT4Pf
dQflxkjZ+Oln4aRD14+L9deUrOxYaTZum1ZpWCLhi0F8tXP/GxIlKWqW2yCN++Gyv22Sa25ti/F3
noA/Vytyubm3staso71DBc9Me1aLLVQKtppBMr5LHsZj3PJih4Y5XUJ3K/mSyIWANu1B0CwcV4kF
DNhdt+4eq8vjQo2PWcPD9xBn2+fMNqtS9o+dqQVAHtrXJ0OJST/WDdF8ZZhLG7dWKZUgTecjIbuV
ry91aXaXB/glhYipHr1YxfMx1dDF4Omrm1hC+SSqPATHMhpzOM32UIFURZIpaab1QnqLpUUvK5aJ
taXTcftp38eqOygjXS1+lPMvepFLHeiHru3VrR4RD9oUbAVjzVm8Z99jaHY9+1aPG6z4iMdbTjsB
tiRLpn9JmCEXgKG+vFC2HcsfxoGYA159FRkoSwZc8uNPpwZAVzMjYCWMfj5QV7NZlFhIvaLGUA+/
xMoFY6LeQEf9OJBPVRrOWZBhyDMUUUxAX8k6OH81rjNV8aFprre4nhUmqLGbWRm/FyzGbkgdMMwt
BEnQI4wfOh0C7jaQmkR0Wt28dI4wsgGGjKrLyae5cGAg6KElEXSm9jwuCCQMM9gcwAy24Ezy1VaX
H/98Gyn1K8ZNFldUPouspZTiuIIAaD2aTwKyu7i1Jc7GFZDwmOoVS6eWOIgO+RkJkwng8A1rUNQo
c0EHGuBnIu89EJ1ePVG8ZHidiSJQ2T6A/B887EZyiI3NjWjlenzjFjJqd/Qnzch3uJT7eoNds4TD
CYH+WlK8ltUoatJ3UIwiDEanrprA93wLZwWzTYYYzTJFBFaoysCqElYfb8aOUtDhHKdidfQL2xv7
dbENIYGKZ7wMH2q4BV0NnM25JKb1yzxe7bXkkj7pfdpIDoQsn7JvG8l7iWW1ZXG+EvD5BrVfWSiR
YVeRCbWcUPfmVbEYOqa3ujYQtIa0iobHfOnZtk6KZxRhJIuN28SEtXXurFzdYgVJqkL+FBE7eL8g
G4g/wamIFFmTWTJNHznb2httnscJLy1lJZMWLME4hOyjqEbLy45d1KGobFu7zYS/PiIuEbHWjTY9
ndQNGEo0MiL5tIT4/TWTkvs0/EHdtuGloNo4305ovZJv+y3EkELds6+LllfPvBQqS9TIZDnVHJqS
3yIom7ndwE9hlzHk2UGB0pMQ6zqLjcdktGVZ+dHaAx5aQfpPewpGvzg5IpgW3hAP9BNAZNw6xSZq
WYQRjoEFlex9aVuDT/qo5ykbuVwGMiiNreNA9/fx9iYyKE8f6jFHzsVd2tMn2snH4H0NRJXTc+R7
qQ9ztleQhELYzaAJAYj/w1OmwHzSmmcHkAAbp0SN7jUGfxbazpIaIoCd6N5ddL/UFdhdP7a05Erk
bUWIrJ6tbpBCeAtbz0UfIpzyEtkBgHlBVNvgPyzpPMjdZEnklDd8ViHhe71ieLt6u1Z6v7e4bmX6
RJFfPNho5GMRZaTBn7YlMYFoHpm6JQzkz4I5gkMTJuTWxqlwHTVmdZL2G4vJkfQvEtkE63AtJs9B
JmeGuExIPJk6DgVz5iYxYmgFR8+oU7pA32GPAenUwJ8JWHkeO5BZsrv4PpaTuZN07ja0ghgDSD60
ap+w1rzEWElHrnyZeLdEs4e3OBuX7H+zj2rB3AZBvN9sgz4d1vu+uG3R0NqCBcRGn8n+hbzJLUuf
ORCLC3pI2NacHihT//A7q2XvHKcRe2wRUcA4tvhn85Mns7POd2ClP0nbIZWXDtdwxOCgnciYqujK
F40wx6lk+aSqJj3xiWOBjY+reM0fzZsrSHrpAaHi0/F9Rs81RAFZaEAzxoPXeNIFsirQfN4M6iCH
zKKsfF1thptp0W8NIgOg73PlrXzatVdJPvsiEE1bljn8XW+oIinRHPCkhQ330HSAlrDtuZX/WZar
r775nK32a7jyC0CgraeZTAdZ62ikHOhXou3l5NvGlg9HyOOSfH1G7BGGqHf2Vi/GPnNv1dXiR2ay
tvzJpz86sMMbbv+4dob7rJh2TrLKSEkShDlwfvXAnFKLAp9Q/NsnOLt7hzcbI60Es0gmopkFypxD
i6BCzGP10l8ZSo30MAqm0lY83Ja7MSKV4ieF4HP4MZ23Tza/Q0B9KeF/AHV30F7FkJUT3PbRB3O4
LYi/AFUJFxBuqhJsow6FG9zb8IsAomtjvqzbeo5z5gyAtg6kpPP4M+mAD3Z95wmEBnPq6TD1KWMC
cl8zZDT0ADk2wlKZOz6p5NyBGFZSCBDutG8D9FZ4TugaAga2+L5iPHkvOucW7ht26KxdBhh44K3E
flQCpXsA8bRd6+E7J8+RJXWZ97uFcsxpCHtMBNMWlEztf/uirgU28+5DayG3y2V3DOBEOYVPV4sZ
1P//AR+eHmKdqkYlJb3r7u4tGuTagovmpfmbDgnjh1ONePPAjDHM29ShIlB4p4mubQ2JkNafbqJo
7m9UWRYrXKzuuycTcc40IRrKNqnuUMBUOJIeJ5KWXD3aYRMX4ZQRpolm3/7FYJOBR+per0Q6Qs9X
71zkPdWRD5CzDXvF82AgpG6e7zOMfcgd+bAUq9CcSHmu0cjk5l2JZpibRfkzDPu+exLZyKeBRd3Q
0SijcnhbqFAgcOOz5pdKsp7yqtDDzuOBdu/61x+0oWt6bcJhrnDRQ4aWn8cbY+fbunVRS5+YcvZW
JxYMaHDWIJgAIxbsmCigWWrDPejshJCVjtUG/SQEIPyIZm15AX1ScR/2vZUODRxukXlHwF07coWv
KCrVszcGuojajNyevBcuwyztOHFkgNKVbLQwnN/VHeCtpBPQmlpWEVsEmSw8Lh0BXFphMIoVWHEc
RBfJ8ffejOIDSrFDrXGOamdyBQKZnMzmqXvzBBp8CoYiaUEphutyRYPblDYPfz3w2JWyMFu8hzHH
a61JDkqzSgUZPEXtS35gEpSMSWFOh1IUItB4DWmqIci+4v84nnlLcko1yyVvUpGXK8fO2Yz89h4m
Jn/mcCW9krSIN+PVtj8lZl5w/4hEl5I8uvKiw7CE5WHM7yEQuzwf0lIgTbbQWJeq66U6Kc/xP+4x
xlw6OHL2d1bbaTDlDs7rk9K4Gk8dFKKdsnAjitmLu7i1meJG3AsJKVyMWnf0xUl1gvCWInmx7QHK
QsP7H2pxyeoBV9W21FBM6mD5Kvwp95JsWO4bO7C47kgxq/DnnbRX9XT+w1IWwlaM0fFAKAqILOT2
Ov+fsiUNaECWyAJA6nKMsQbddxTb1Y5X4diKuQw5qXtWRiqWmCspPpX8JJbV6N2HUNsOyUr6y/LS
jyq34QYW5ZwMieUayGNa8DbsKUw74cB1TNEyFlrtmryjGfoC8Et+f/Ya8ExY13ouQ2uAtdBwxGq5
THuw3JrCNNHtth2dexpRTLgBN8cKwqq8gI+gHgDpYcq0DHeRoMtsUFBqO2s0vvbvAit34aMF/vlz
2kuw9lET5LOnFQY1cww+VCbaJVb4n/YgDxWmj2u0a5LM9LyQmIK5PdR8p6JKeU2Dr6NKqOUAwrfh
WtIlIJGlrZtVC6DAeYXbCQGhbXt2a6JRD6h3LfZyRth1o6L32WVcTuyPe7uocp3QqrkTB6NezVe6
UNXx4QrUw+UC6MLzOlv/bALdBuWzZD2Ts+DeVVUuj/uxaPvLiRklXr5MHAANlvLmoGtviccWyKLC
BMGjj1VZvN3HIL7QJrmKDwj9eoXiid0sKAo1UoOwNw24wqYpgup+mnsFPy93KIQXoVdxykvmNEhy
SY0trrp1BGZUpTGHGjYML1dIipUTh/1dt9VKNcAjvXOWO4XmzKEeMHj1+JRSNa2mjaMgkcJTtiKe
arQt7rq9HazSj1HIlUsFJDZE8XYPxVu7kiH27KDfD02KpJuRCrFLKTnsQ1NVKl4nKmF34tod9Nuk
7wqhhyt0kdvc9XsGqY8gqGPM7PLssjQjGT1487rR6ctnJgwtS9X0GU7koYY1LO4V6kVC0P5Bu21p
BwrGT7sDvL5XG48R5+5btWb44Kq+JfHUckuSB1uJN+ySpim3vvCI1Q1PjPu6p/dU/yGdPCEX51fO
TcoJqHTp6rIq8UwzbIsLWyQ2gkGHPDZS+G6aKzzpEpsatEY2Op78vhxrDknDv3J3KzjA5owP5H5C
ncdOC7crLit/W9U/iT4HGwwODR3JftwmDpvTAnZu65EOOjc6Hlyyj0Qr/KJeFKZJoR6NRSAW27lo
odrCyTsCbAs2UKwaEJYM8Y28g8aMb8+zSH2p9GuiLV8WnnYHS/Y8GaVyKm19rIa7K+/Euv/itZVQ
7lEMAlOtaCCIhQ3VELTWfjovZoTeWkxCF1A3gmfQdSrnuk8lMetS9M+amgoFme6JuVB2Cd2Wx/Kz
8UQ5tYicmDW5t/5EempJkOLdP33EQTTihTF/aOXIv9lXZqkrRUK1COfrIGPhcEzApT0dAasCxkBv
A5gZusMioKFMopQ+z8nJjrLjSQWto0wrPrj4djWi6oYjj8nvrE5jvtVVh+HR9stxIv+9LnbUMut0
F3r0aMbwOoNhS1gB9rYcqOjpkSut9jCFVlP9O2rDfScnjjSxSzu57ewuAoTwW2vjb+Xct9wxFDs/
JjSFTnwMqDPRRgjjxhhedV/EXU3egQ56cEp8vli/Vd8pcAmIPjpNylssBrTQYII8mWM23ji5PNm/
wZILEG9aoNRyDH5uLKEGfwmGfC4RvmBIxi2dsjcFOPq+naJQg1vflPM5if1U306i5Vyy+sCKnlWL
5ZXaBYAQhMw8pRS0bapkoAoMtAXptFDFm0DLsrKk90JqDT/O/6DWtWdBAjPDGDB77IVm+ejVwl0s
tRUYnVHXqUqnDM60kWFuCd0oHXX7Vg8K2FNdsI2Z3kd5J5gcilOL/m2effaoc/X0f2s+qk0Vn+lU
4fp7jw6rjMuKpPYexICTQMtkiQdYq2yPWDnXcOyaiZ9SwXfjLEWzpiSnBuTl0bIXZQ/F43lhz4Lc
M3WlKF+rOnHz9TA9YBRAWVjC1rh/kvVig9eRDVQ7orR2zUFYDdeR/gTGWgwal14Y7cfVE/4YZH0z
4E1oiepWOwyKh3KEECaIjWOP5npISwO1OtkOMI26jA1MIVlvKK1q2TB2DTkG0FvKC+g4yIfKiwPP
kiBLRqfnD0eIvxdZtl7WcRWnH1ejSSqmAJ6vdKLIo26ZvuWBOvWozsh1Wy3QhAxxWwGS1zpB8eGf
eaSXS7iYxpHXJIxf/BNr/EKNXtEy+AWN+5ABikduYPETMX1SvLUcGerv44ZGt+O7U+IdDPrk5HwD
lA2QejblnTqgFi17UBwZyFSzK6QnuVTXad3bdBuRccqFNC3/Eb3axVaiHo4pC7f9eoYWRGTsHNsD
lrDbbU76+/lfZHQEHnJ8TC8x6gw7aK5hqaxTdf2OGQFfwoD0pAZmy/03y6P6a+DCcqARzTzrnAfC
369mZqvrEuLKL/QDUbv+PM43OQBaRB5UCHBE1Gs5uAOECJPk7vzKeRCe0Fd++UzpaQTzhBwIi4KN
wOsKLBpjzlPelPKp1bFvMiTM+WjxOhBbnKmecpXKlyj8NLXE4/kZ2w0wkFYXlxtTsHCCxvkLzDQi
ujHeIucb28+YE5BGPDwVvr5Dk11vfHJpAapLcw1s4+9ZDOGoLKHVB9Crjh9P/0hV3t+6tFyf+a5C
zAxVU1qjFHJ8Y/5YxtCgFWh0/wsaUGkpHGiboEbt9OCuOJzLvYxIEHYOKNVw1BTaUE8IWLcUoveL
MkoroRBSY13GswKg74w4jGQetwfn4UAJSYuoLITSK6yB5NciQNtgfkSZypzQwUTRtpldS7sYwiLf
RILGG9RFkF8IAKWiHz7m9f1oypU63VLJ3qkyvURVj73cMcMHgK7E13tOPV561J27iAtdWG1Xq84I
LbZDwrLR8I7rBQ0Il4Xlh9g8uIb4P2Pe9RlRcyJ6ivylw506aKUgtC71wJ/wxdlQudmoQxgDyMWs
xVFuZzGujQfWau5gTPjM10wkOdlAxI0QKweqCn0sU3uVGkDn9wn3C/mvsFKkBLv0vQf2bEQYryRK
ULt+3SAFQy+h8Ppcvu45Ymp/TD55h+4NVJ/7bp8xX90xkfhdUMOWJW3sPUtTZ1OH2k46CuQLsmX2
rLAqMdOZ8gJBxovuMrDK6gKG322/R3m4YjGu0zDe+gNZiwsL0y5fTU8c24knkXDR6raztXgi6C2z
cUQ1JVQBYzJPXJf6XPLNcvGr/MFIvqUF06BAz5ozK0Lv3H1S/BYo3BGdRr6PTaieoJpp53fGIKxP
iPY39KtEbhq9L9j8hFF2kNGu12+fuGrSOMYuq/GDvZbjDrBB7D0x3n+BSsICiCiQk5hwhEuQWkss
Y1VHVt+EX7XSCMFDg6GEDfv6f992Wh/yoJM0R5ofbbjXDy6mHESgPDEMtpVBJOCPOhfbAfTAX3pn
F8AyrHBeXfKI/DqQpEIF5KIWX0RlgXaq3F6qjDojyrzgFh+6AAMaYkYaaYIt9sT/Haug3z8qrcS7
luyD0L8WqBOxe+SWy+wZWrHQz9xoEXidT2ZM5c/aEH7gIM177xygCBxAOy6svkOf2dB8TpGySoYk
Ou8faQDkZ0ORbCLDUXy0lNDBI93rfZQu5j3hYm/tJLCylhIHFzfWTmUQhKLV+fsd+8/q4VynZshA
WeuLe2+s4xWIGziyVXkksortddBPzISX+hQXJVNyS4cC4pWdwkd4XemHPgJGic+liXRT6KynA3dA
oP11GG6IDHtyhOpsDIVWjW7+wxzzonGX+bqJlwVXzwFCSn9Ok4cpFc/08TXUVENERGOcwqpiXG9j
z18pu+CpZKCvIUOIM77hp3r5nUxAOXCF88o78SpL1C5TWX8DrMHW8i9jGO22nML87R9VyDolzUAg
AlG3I2JDT+Dk24yYXJkMawxW7dA43kNvri3S0rTsvAvtfaO6TwoFEuw+IHic5FCIL1k6c4+41NXl
WpdbaBa7CmdfBROwj0+7jfaLfm7Q3hi+deSSnKaUC8Cd3KodM8qBIDUe4gi1zqeRz84LsZih+8Yd
4IH+Svi757kegbv3SuCkIGAXm8WXn+yimGm8SyufvK271Hmc1IM2KV9zlazrW0CKNchdrsTCi5lR
Oww2arqMXtFYOu8KcQ1gW3/cITgvNPdmEclIOepacvj/mbHVwwm5Zi1FD0WqYWBHyNQUz3UIWwbO
VLTIxQbvFVxrbfT+f75DoSm1UCko1aC1isjv9U3NBRL69MC85mKJQPLoP0DbcYhUgsWK48mwiN/F
k3onKf4l1s/x98OjBAcW8yMft/iwY/3Urc8A+SWBfiQHrcct/rAeBjtx4bjQfwElDhKYI1IbVxiG
/YldPt8okqsr2vcDSlsQZxmXThJixtjdutKS5Ku3X85BC49jQak1Li1Ng7kSNrk+mAqf/fpQ3T5l
qskIL5SKhIlOcl+gqgzOLE61WWDtz6BcHn1ZeZ9aY/r49ygGK+uoGd7KoOYkvnl8hCla49JkzPyd
ve7VyfXHKIOibMGuzZVVYIQqAcAvyrMDcjzIuH+MQFk/hSXZwN9dnZQgIZOvqYkVN+BCdN1FwBQB
xqP6BS2UniYP4phzabam1B66/tI/WluxBQq6Zsy5quXU6PV55l+epQIher2m65Ecu/UeXDNnZ1s/
rGeWDLWoqPzFzE3rME0LcENQWvLeu3FCKlfXZEP7CCzx1VFKFcxmWK5SJsFnaDo+SwzejzSogtF7
VCziNUtT3IaH5X1Vt/e7zVBvejb00Y3bAqgMxfwlJ5ZBjSqpEWBlpozqcmy2v4in7vew8UwPiIFo
dfryR9RzbDiX27O+sig5J/LNTt0LWNNfV2TM6x7QwJ2kvqIAkn9C3cTJJ0iukWDDIMrAcILXEhts
2fQhuJ4Crai7VDpFxrFH4REYG0Y04sP8GkLEnxeLL2183edHRiKvlt3C6IkyzHRbheeMkyf1VzgI
rIGTkQnvcszbypyYcVYPXd21cO/ewzv3h8q2pFxZ3/yoyWgWizSmjomgE4MmFfGr3M8HyC4oFghS
GNafrAiyoFxzaGoed3RrGCCKcUvc2mKSUdaPSDisOVqAiorkvm2YRbbzsZ9tIlKekxAU/hh0hyos
SrPd9PZLmMVoPRaNrth1LENaOwt9wGaZELX1uKC4D6dgeWadSReV3MVigUFPHYheo5qv3Mv29NVK
JoXvaKXkPc2+kNB7A1XKT/R4LcLjihs7ZxkVKCUnQEVrUoBgiIcb8FKdf0ESdmFdX2S7zFNkHWpM
e4IElA4KhuUdAtRw+X0aujiWzDGo1KenVJ/dGjjPRO9uA313ctuI7PGJjDw1RWt6I6m3e8auAY6E
+M0364cvSI2oQid2ImNyEl4GLrSpZI3b5Ikc4vH0HZ3riNFey4iVyXG2P4bFLEd0sPnZiNJWw7Ex
vcjB2LvzQmErpB+fBo94PlERbIhYadBaKHxfCkLrGIyBOzrIYXbxlMQnITiCvU3Wzr/jerVyn9zE
gntEJZ60f/jnsytRphYOt/M2vVDYrMWEK5yjWS5sfp3fl8iP9ocVzmmv4yFdR/ftD7FoL7nqVZjc
FANaOTkLdVqWra+4IUT/ZLEFR0Q3xFmUGYnjQLhFXaLhp7XqCSkM0xSGn/OcgF5L9ljWXVJvTXsb
+bsa+yV1950VqunGMlcRg/iBfE1TkgV5QHuPK4ochafLz13JlkAtQcS90dLpU9c+SzcE/5U/HwmP
BsczhEGHghgb8BCaseQj/MjBdcrNLBruO3ajQNIj6sEfZhJ/9fsT+jvGQQOQXtV7thWFpEiVdeiM
CMqqdXW0Ue28e92RHNYLZ66keP16t0RWf7aDnMoudEFUNQr4gtjUyvBCCHcfr3jz2NbQI0KdobBl
ziztz6XpkGskTwyRALO1KVDv0oy6QmRmjUFgb9KUxKwvhvA9lWh3Z/DOt/NhMqKgftk/l50uXGfE
T2rwLYua0hUbWpz7LmPWI6x0x/NqHKMK3JPh5xbmWVBX4HbTuP5RDlvFszjquM2Fa8ese20cD1Ia
Y9d8Jq0pIjJxAo9j50wCc6J2xXXxRmCmQ62Gjc8gUooYNz3xN5g1BpsgulBjSAJzNr2SX8iKgf5a
e8kM1/i0R39Z/fuYURogO1eGP1u1opwP8/demi9u7hideczeZRQak2D+llZx9B55XqGobpkrqJCS
RAA7NGAzWCn72V767+DiqoLiJ4EC1PF6FtnXoV6oq2Ncyt29FEcTdE6G/XcOwckBxMO+oIL0qRid
nfw42pDReZMb/oGBGla6yvC04xEYYIHb7DtVvcnE1Hto25qdRbxDNLAT2TTQhQ2nZPqx5Tq+uehN
yYxrY0mNNKlVMmh+oRbMLSMuSYqvaVDXgGd0bfZRwZmv7VElrQuVI7+UlqKJhcS/Mrv2E8SxUV9Z
GC3nxy3IYHk84u1qn6uWgwulPc+Ji0ewNTVGxxixMZJ8QvfU9MwsBVk0w1ExX0vfUTj8nymueya9
LJ+W48ZaMlVi3WaFRwWEG9IMc2ugfL/ivabwOLZem2iScWLM0OveNSFplXkKqftJl7F2O3gZL7Sz
qJ6U7Xg4AkJy2HhMVnu21WyjuLYPiMhH8tnixAybU+DMUCD1DlnhyDR+SVMM17n5xKs1YCX5qeIb
sexhjazcwirSAu58QuSrag2MbMct/nNxuUWyyRR0A3J1k2Ws/ocYa4v7jEmMeGoYVyvURjL1Q5lI
k/ExO4ZMig595jMAg4HaK+wwlZUX55DCA5WgNCHZ6TtnLhuW01FS6+cAQ5sOJXq6PUrdzgiLwoQs
wQuPW7J8tZo/klZ9s+xqQdzXLseKf5D9XAcTJibZzhqKVXnQLislI1ueRPPGgPcyBS0SCeTJwTnc
gxud1uuMM0qdRVgmprP3zrTwzwkI4ssyMpTPY76OOV6qf6in/NHTldID1oBco6o1rFgEru/OvcEh
KFyKRD23sCyZnqh/pUKhZ3zHL5twowEQ31yVG0+iFgFAOwWeAJ+dv3JPxliZcxV59zbgWPKlgubz
2nHrjjsXq2NwxbDBh0j6Kkb8qfkGehqlkR9u2kySzTQyWNbMSBEpPlxOcC+eoO+w8jmE2UEYB0gt
C5/P6nCoLR3+FuT/Fh1y1uAOkaD1doTgYmsEML2qdMpMuJmPO9YCuWAU6TqDy2AjpNFgIvlz5Zlg
IBWfOVsmNI+Qe4otWYnF6rr8VomN15uruqbj5yx4g+vWBBaBnH9n36Dsp6G652tIkh+AV7X4XPt1
zqAbWwdu/P/58XbFPnJ2ZbEvREVnEcr5UzgzQsoeCWd66aWEkRfythagsXwOKtedbdA5aE16lJ5G
3ZPrkyPj/rkZTzseotRIEcNXi8wow3jbUIeB0q9VqWoIihboaR0kjagtb3ilab5Y02wRRzTo5sIE
AUinZfRGJP9tVwS6Ndp5atuX52tfhFWriCXHne3oemY8F337fiE5/B5REkcxQZ5wYdlX5s7kPrJ+
YKb7yXA8JCaE8PNxgzbMM9E4dg7U9KZ4UZyXLQttyfH6C1fhdt0NZKWCb7N6JO4eX768XB+6jWg6
z2tFnx3M6rpyKpwbpEvpFJCIi/Q5fFYw4qCPB1aid/uRjRHXAFPvoyYWui5pfohwzqKzQefTQHsB
Ur09P4gRKSh7QC2JpkJw87EgKqUROmyPGs3vbAhDKafKx9F3mMeHCrdt6RMHTI/phUQ5eYll8zWb
eik7w7UXhcXteyYT9TC3UbmrCHqoxN1OIavspeZNlscA2O6Ah+F4jkIStkvUzp7n/UlX5l0xlpbM
RptKjouAX7N+q8iB9aVt/59PLUI38hsQ+rTPXC7s9TttGL+UM1X/YWahnB/KlHpzW4rbAFIRPkQd
D1iKl7VUVu82XNgF3oIwHu0NXMXpkh4iblyOyzJH4N6LP9ReTouU0MZVn2kiSEnyDjypoIfUV3uN
Y8Q1RLu1Ssm52eN6N1zTbR8r44xbVmRf7vD1MVPjZiEipvoH6ISBajcJRMO0XJA4Ang89C+OKh8O
CeWGuqJfjlMOmDRiEoq1SEI0pM/l5R1ADsuVym7lE8zQBT9r5sYPW0jvlQSrvtdf7GYDyaBxMCQU
3cZ4RvSWNNSpzllWTQKxdzeeRPYSpmzrVNy7QLdnSmmJIMaEw6YhgJvI/zLI0kQBmgXBJIvv5gcJ
gwFVlTVusH/g0WOf7Hyk4t9rYFSxYRml30TDtqWIcXYl+/oPno6Mwo/a5/sc+NU+zqR/Miu19MAX
x6Tu+UyKKwFI9RwIZf7r3QNIZ/fH8bAfOQLWKdbOHmdGIHJkJ1uxV2p+FxbnHme8fT1zEeXg+sev
gvxscYsRVefvi8S/B7xedcUwDTkdXkcshMB/DhFKvn1QJ/HcsSPGjAjm4cEpy1C76qy0+cZYyYRe
o6nLvVAgA13uJLxJFgNYkCaUqVqQIVGjGkaHwDkfmWVPFFeKixmofVdctUL4hbiE9ZxTOcAlwLkC
AnTFNohjtMS5PRlTX6sKtGxQMmY87edQd9C0Q50mmxERDy9ubk6CfkH3FYbRk8raOJX6Egzauut8
SS9MW7wKvi6mYtQw9KeDrtaHutXUnqYuT2XblaZzxZg9n5YeGvrRGV8x2WJHTfEUDh+zyb8W0wDs
EuABg5Bes0ug+KawLo7ysrVg9XFoqKRTeXMkslXGjjFuR9+S+PaaYLLw7KNmuBURV/VWZQDQzGJG
DOEmPUbN6C1x2Y/rKskt8QF10kWvS2XUHsIVMPuyEynvsgRTrsF1GiGyS3R2TVV05xvxbLUizvJa
bAONgsMKw7oyf4qkTXyi+hdEXFp1VpWQkTl4c3GkzuofrvbDhnc7KJxmlFeJiwa1yXUzSlIxeeZH
Dux90z8E8+faYV92nfPd3glQm3dBtnqfTeY8IsJ0IgnaQUR3qfR1KeWBPYKAXUJE48Fe2b/WCNDG
/DZ3tgVxaQTnRllIMvw0VjT7Et+VnwYFObJzk6TO33XGF+HGSN7TqoIKnF4409DBWdwIv6RtrKfk
aEHGZyB1UR40idpqlYtvNRhj7Q6cNoyos7MkTbBj4I2j4EFzZEVE8mr8/WYtnw8OsdU6WC1KJglW
42ZV0ME46TZdiRUykbUJdHuCTPyiZYK1i4SLUzP3o+81D9Ypj4b0iMWANCHd0YAufUpH8RSqixO/
V6qENn/pq1xaz99U1pocrLPTZNcE3+UdGndFSrViaQ7r8i9DAzxz4aPe4JZ7SGFZyRGqWKKFSaxV
EqiOZkc5OE0QC0IIlCL2G7Jo4VAV9aXD2wVsmOUtJcjE66qJZCQQSpkoyMe19K57BRlKJKJGW6sl
qg6iEVTYd4Cs37Pg0G5v+ybVy77ojuTmH96W2O2DJ2h8+BEDxuvhjWuFePu78f/I85Em7cxL4fqq
Y8u84oCzRZXi3MibUo+4bFZG+G0uLC0na9PcoglzNdeOSizy8MRllfZB+Y3SFhjf2ybJWaiw3l+q
dC5w5xVWyIoX1903wAu7wKfNSnkck/UaehzyQFYvw0CBpPEPik6tglZJEE1Q5Abq9ulawGeqOYCY
ddSuYPanq7/b9TKToKX6qHSs0VFdM12V4E8F+CT9Zz0k3KRTbTzunmI+mXsHUhLT2gUojilg8u0M
ua+/khIadq4p0vV3XaUhwXM7JPfW9as5FmkViad+awU0isMmvkbp4FlWbYskcs673dG3yrnXqOYa
M6GKRQS/bpxR2gSPIh60GyOY72bVHnKI7s8EweySjNquibpGHTHB51w5pQ7EuEdz7MbQE1/jcoFW
YRhS5GHO6VLwCP9Jg90acLOD52+pNqNTFDFNPfp7eqOUV8X78LbeKYlNFIWSWhXBgZzE5w3AzqUX
pvBrRyq9cDtU+QYqTV8r8emOQZNzZPD19byJnAa5bxVB7OWyDI9qBOl4xokP0NZC+smoG0jNoUtB
tjiNdyhMnGA6w8Z4cgWFNphihyDs1S3wwWXAEeg5W5k6srZ5CyTDoQbjWEIgPbLT41payjMGHt3k
z289yVLGV+mUu26hOV2zphapY9ZEgH/fBFwP57ZEgszxnHH6GY8M+Lo4XqC8S/p7jo0uql4e4UWb
cdshinapPxxDC+SG8VgNj2h39pmgyaEL8Pz14FWWpuzCX61SaWqI1WM0g1+SLRHU4/au9FHBXVV5
DnnAmjrV5FKyp/4r9ZfuXMXLpemZgtnkyot9s20LDMV6dajJR7BoAj+R9l4PNGVxa5h56nQ276bj
HRxmqW+J+O59cJhy7UUXLctS7IBxkyUF8didYSoGdMxfh4mgy44HNiDf4UveKGdhF0ZM+h90zbkb
4Q9rwlaFz41Fp1vV/vGgGCLaN8jgOBeA8e7ozVflUiqv2Oey8Io9H2I1CF2GhlB2paJgqQvzEXau
BkN5BU49qfwmtc08/c/tsCO7NlemTFJBYv5ytmvAEu8OAeRtHrlJvgre033q8s+jbT0M64g0VDgn
sPN0zFVogVdTS61aCgtCgHAyeCyP4Xi/rJA119Aor3IFB60ihzymU4afuXmq/e87ZHjWjEzBzqAw
7H105KvlKDMSN3SLwmAqy6tBubL0d21kqiO1I6wH473sVwuTdokBn/L9PioLkTRgAbktIjmb/5G1
A3q/pctontP2oKkI52oZJhUIKkSDAqa+IXzXmveLlIb6BGiuDaZVwzaDsdGCfn8l43pAuIrT+vGe
uBWf0jGszVIE2Y9umMFduaNThkBMf471xXWpUU62hrMDK5y3bWLMPuKiNc+8Xu3K+7OlVCCwlWi2
Ci1IlV2Q9FDfmjdxv87xRTSqEZrTszvFJz4Hglr4hLvqaA2iA+izaPJ0+m2BXDOiRYjdbcZsiRHb
El8mfYeNkzDzxnnT13X2NheY7FnBM+WbsLVqoFYxmpxdWp/PJW6kscSsuR7X23IgW812N3N37mfM
96eEX3B2SUDakyL6OZeXH5bFL+oW3PQB/QGM84vY+8rJjk71N3lkoz1fTUQnI5WuOU4OFHvwFN1L
NOzVVzg7G/jl1CoNZkJEiy/Rh4wSVn0rIRDpYASiiM/sgp+sbiFZe6Xms0KYbRNmw8S735pv3e5F
b6uP+m1GeH5v92Q9NGup/sqCB/GaZbHr04GUQLqO8ftI575myuQxFH7rhhUAswaKjyYQ/Ck9nZNZ
6Qv98m68n0mWfbypXsW/nRwt9pIDrBEgDbZNkGC+eWcHGFkuDP2Znz0nXx3VkjmFLvhF+PtggWgb
IOoi/gS+woGai7MsNJh1bb87NT/w1Tw82zC9E6iLOsqjEKjwleuPbNKJfYd1KX2UG5Vyrt5DjkEa
HGiRjluwngpwEmDsmuLEK2qsBds+raTbBIlvuW/5IFT8Pvpqxe2AzzsRSZ0nMzf3WLTks/U+XDqZ
LT2NJ9QYWZkBu/PHEpJ5Ymekkhiu42KZ3NHLI7wkGtpozUhkHvFnAtQxuRjb/h1tynMOKNmUFT7/
a6muDb6v8yQcgs69CpOp2MAObegy5I311IIRFFLP+ApldthzMsiv++8j+4Ahd9gtXpYCM0Ya66FT
WtMh6DKUWwNfaXDa8lMxx1eh+nXkP0ugZ3sYU5sVrP7WX/WPqxLowN4KTbmAuEsknQJRLazpCach
7g0VLuFz509JO5LMuaQA9IipRroeanIpnuSgujxEw4M6sSgjG9nDuBm97cnEmVlN+SrOCYtbhbgR
weB35UjH89d2VmABcEF1Du/iSXt1KAuddrCG8hb+pb0YTtg8Av4BJ/WPzxg2ddKl+YgBYoUpbiI+
U8vY+sNZM30/om/XcWqcfVw0SreP6j97BARf+EiNere+/G0O5w3sLl7czseCnT3SJUkbk6bS7j13
240nLi8RqoAyBKcbdoWcNDGXDJbk2lsWF2UOi1/xXW2ifQdRvRihy9dCP1bRtujm7mTClXHkhoHw
mCNXZII3xVu/tBSpdaXItYPczyWk2Wv0X6zO7Jy4mhTkCev51QB3M3f1nwyO/qWdjHd9pFZ5JfUM
2EDFWPf3KYNsWOYtzyxBsCToyWj2lT6Z33RY3bFoDA+VaTBliM92m1AlSNasRuk1MjEDXuxiI+pR
64/BklxS3iYMRvUpWIb7Mowf48o3v02D5j4HfGicg6Xe4x+OHojkfP+09j9qbUcOx0ciELFBrK9I
j/ffkFZnDvQpE7/MgiVy+Q4rS/BymaYT0/b44e1ynDlfJhnVQJDfgUL76OiehYHjxMq7YcYD3PZP
/nbHR9ERKjvwhsN5wD4esnDSTQMOJy4FLcwsZy3ntBZTd0+AcRhRFYIIGLTGUjuS0E0V40Y/qPl0
d0Nh+LgHtVK/8nWA7kTL4tAxt8NBBhOlW9tXVE9Wv34zE1ihF+oHebsw3wO6gib1HgQ0hn62Fe6N
VNqDrU+1kAVnJFYMj18xoJsXnJLMpHX0S3yM2rKmgM2yWS+nJF0EvDHZniXvRwRVlqSXfTYmS0HT
iK4qxux3zR11hNfpGc0N9ZoPtp/f6rFDIst5pQiPrnva1mJIuYv0jIHQc8dvFyuXILympbS1ttDW
qCbO8tF9mG638LoEje7s8LMcUfIuGyymVcX+/t7UR6RGgTW75rqDUxkijHc2bWpJYgzI4t/7fKDC
CBayRMezYqe6g3YF5uZ7Z5FyEeDSY3fnCPTkcrGuISMA9gMvBWAGjCdadaiVnHwrqAxACtN8raKp
w3y9cy6cqqAmVAa7kLTd/8RgkrvQbyU1hb8hFCIxvZc03EMM/u5H0gGW2Eds2y7GzL4rPb8JKifK
hc9H8UWVzAu37sjT6Z+X2oz7lZYhC97Q4zlhPJiF+N0Gs7hTNqBqTutsuTObCAt5agdp+6NiOLmA
qKKFQ9W8+1y+PUy6u8ghGg2SCfGQTlIlbnZiXDN1It7Py/t9hj+1o4qTHi1I9K1WhkAGTZKt01tF
IDh7AwtJ/S1K5jm6mHJe6BiouTs4mn5sEGUgAv5D9KTD3uc2VAU16Uv7qPlYPrQxoLkbhStPLJ5F
nMhz6DKChH7odwgdx9q10NADOkN6wKf1ICDbtSjHqxxuoUEwG+VIyYXLIOfeOx31JMDxjsgtxMU2
cwXzLA3s3T7Yi8L0sgDUPKNHG7sA6Hxz+mJEfkC51wq2vCRsHljRr10snSbYa1BTu0US9Y9PTn8b
499I9K2uTrlB25Y8SbXxIFI1vsfjDRK2CuQsgSoRrANv/WPGz5+ZBigU7X/NYky7T54drUjzaAqi
9O0+pDD9lO975AwZA+mLSgK+N8OwLNEUVP97ngt7SgfzsTtbRN6vJHBbr3n3EWjkIVoLtwN2cSmL
MQ+KuzLLRFwFx65LbcXZ7/qzU95YX27HJe+GiwTB9gnF70km/zDCu7LhbyxnAF8Sn8lox2smwNTz
QZjj7Nnt7hZXNQYlQy+5ppY1+v5UfWOl2TiGr6aQ0CxXyxkuJuHkAishX5y5/XJ1p3JJw32ungL9
USl73aLx6FxYjKpyosp9MvFiWi3GnInCeOvXuboRfow50YBsRTWh6c/fz1WTV2NAYH9I3nuPWTjk
0YINbwBMLRWZeEf8TH1/eZjQa+3imD2NxTe3jL1hwMgu0Tb0NC5QrjEhBFcCwE+/d+zSOWhzyI6L
uLfwWjmtmelkreBuHlv+Be0tMe1e1OVQG4s5UzwaJNyxk0C5yg0wJwgmWuo1jEEQEnjNqIBSzEQN
w/+vYniJ4763vtIcXIMCvr5OBRo6PlWdokcRv6q8b4kdwcThLrqnFBpoftcSEX5XO8oiUVH7PlhC
rbukDfS5cSoTCww+zJFf11xtGTnRVn4Zo+yxIe13s6GmA8AY+B0p/VISmPYrb4aj+0F+qytX3GNd
hZTLV/5ho+2raKYMh9RXPSWnoa7VfBwixZFanPwHdtz1cqG3Q5f859JVdvCof7RwIiklhnE2HX5X
Xf9e6OGxJbxQDttpy6yMv0gVZd4Ey+DRg/66oD2vLGLCrJ88VulWT1FcJmf5ij5zkDrJ7QR97ZN+
e+gKemoxr7zxqISidA+mWL8DqHvPgZYnefBaePXpu+zxErezMdiJZG9IgS71n2pvC6giU60SLDHO
ThrhjnBY2wLTQIlfBYMgTCLczWTs1RY1WkGmlCNqDFBMi/8mvtH14Y+de1NffdhI2C+p6z5ck52C
xqhUfdJzn788t0lLqwirwDQIePLiCcn73wTTZu+q0LXIRcYANotwcNTYKmknz7YFjQBNx3EIUBj5
DUDmIS7ArdNwElQUlm88jE/tL2Yu14pRNnQlnLS8O4oVze4SH9vyaqTd+ddrVluVd0xs/ESgVVRD
CI7+va1zfKVumFt1kMzURWJ5+zXACXLxGpq8rRpv8eVKGc4pGcsiYB3QBIuQuhfgoQrZ2YijNvUw
6c/XbpessI6jkKZiTeQMIxw7eBpSnBfvaLpYAOkfMRBGMF5hSG/D06zu9ocj9roBFvEpzlBNQt7z
dcvhDQjZEVoJcdInihUbCrprh4nQISoEOfvLblsYW6OfqihvbN69WueLxLYb+YCX1fk6JM/+oIkW
P0XhyzDSnbr1cgPgEShxYtZIKLXqvnBAxFQcEAMCsg+FwWUsFlYj9LRqpdWC7K/qQDuvw+FZLCd/
tfTeqPAMLbcFcKX79NkdSWU+7B1U1KqMesBHLPy+ysSVSHdYV490EU7ZTDDGwlGwKQXrKuRFny3G
BuzlZ8l05p+L/1gEaVHahcMDWlafxbj46KmvOgRHhRl+EuMujrdw5eqjO0HEgiJaVbIPSUFACjvw
YagMC2ZaD0XLs0wE9mbQNxUn3JrKry1DMp5X3EVSqrBV3ylaaJO/3Q4PjfeOypM8PybRprcG0pZ0
aUjMLo1uQGynBY1+Jte84dfdj8tyMMrTe6y3AfB/KzQt4kQJXzNl2kc1ECp1Mkd4L4xX6nvG27En
xiK2DSVo0TymYiklSJXXBNEeSs+f2XORS4cRCk5XscDFwC2QYFdCwt8f7dyMcKS57s+h5/P1A58y
Kt+BhDZaSNrpV/YweAtqjLN6ROafX9z7D3qM0TO+9DUo7wdLo3+iupHsknNuBNaPdn3AkrLK2TOW
nnbQ1NwieTYW6vx+R6sldLgyb8oNDYWIJTKkB5DjtCqbnkPuiKuHS+gf9qL6z3zmKAuZlWiu/YRb
Jzybf6TgIywna4ocNubq81Y8GMGTK3jfB8cgLQmK8LHsrIeG7+GVwLE54b2qq3at/62fwiPL/MJg
8IhRrXhU3sIIBPPu2kzhgyxociFCX4EnJ1rB/f23SU9Lj/4EVRtg97VosRPzmkXRBlKyOtuZgYEi
Vh+EFpH/Y0Do3+anWJCF5GcRAlopH7yyOaNo6wt+Bfivr/O7Q2J1+ucfqV98hqsYI/Sx6xZqDwI3
nP1d1rj3tmV04bcQPNr+mNE0aO771kKo0ITrcYk7NCi6JwHttWZYl+kZsAP6fXX7QSSqZGX1JQGU
uZtoNtmMSeXaibGdcy5cq42JJn/wKhc6rPB9+lS4UpgDWu/wKaPh+JN91UO8AGaF11+P/BKYnF+I
r/utJ/FSFzQFTcyvV+RCf4Rnf6fTL8logr5sT1yib9YaagMwmBT2vBdUI7XScXwJrG9zbPiGvBLu
Nhtu5uG6ul7Xz+yBKYkS2uIybkstsCfQzCcIlxd1lCe5tLZ5zISfysXeUD3x8BTGqdAcos/7lxWQ
OELYOrnFXI6FyI/XjaOB413Qh23cWrZfXQGfXbw6ZaodzCr4Y3vUV2zILKmXioGwOkcfJEdGrn6v
ggKiJ3VXT0vEk3+vyW5IT40Y5Lu6ZuPBtLeYQAojqh9JWEsw4d9/K19QFaKzpI/UpfQM7n6ffdW+
dHnlux7XhS8j0ebUc9WT2Bq5RyUWS7J2G8+82rdN3HsrahHEUuVmbX6gyKeWj2u/HQ8wSMuP1w8Q
gZXu+9A6tGQWSUVzEdlR0dzxSBhSLIftKN4GOUqz2lhbhaOspI0DuQs/E+8Y2Cr/XZ3UO3bCM9Y6
Ae8G7dQt3vu1BllRhlLQL/fNRN3htIrR1dwS2RaYBxpjWBknCKVEX7clYN7k9BW12uaCUvLiPorE
H0MVDf1C30J3m54EoNOQ96tS34FrSJbWT6YRZBNsrhtw6bzXboFtzShhZiluzlq2JrehJDy3uF1u
AOrbIsH2AEAbJptFLLFweMBiVc/bsjXFecmzL3QGHVO4SXm6UBQ54LdrF7TTkQEmxxqIhy0ENTdJ
45qKDva3kM+G7zmFXUhN4vxV+JUid4YYEwRg6swoRBo0FQrkAet60KjxybtlYeuaRRtt7ISTM3t+
euUWv8iD7XwyWZgxoFDFCkDlbPA+t1qeEau3y53Bkzwgvx+E0v2juJsNEFGYVgMwSHzwcPwsXmka
gbDxsKKs9omLKYsbrJpul1yYFGIeUhAwsyY5dPkMKOdpJpNECVRXegP3Bb9on7A7r+b/c9IE1Wd8
smoRmA1EF/wodJyYpiQC62hax/dBTOLDfaQEXbna0rAIzjFrao1VqLzEyLjcBELHiI7SbyEJMcVj
zAkAlV3lg8IFzq+ro+sSn7qkdIrEkgkoVt+i/Z7gHoyJOCSmc5DgWWE6ylgnC98j+PtU3zLcFv9+
TNmU6C5ljeaZm7aCFyuSvuZcMkqwQpJv394iPNjx34aNRFXQBmsbeeHlK0J9JaiahIB8PRD8DL9s
b+d6hnrleuHuwvPmmA/Q1uPKPXUFLOgeCRMnmNrvh0PpyW6ZNtevNMXG3KuShZCkfT/Co7DCscMk
pNMn58ZQ85/cMyn+EdHZW8BACoEN65/itAFkw2i9CZyWeOzMZ0Ti0WusqhY7+lb21lGuebW4Yvjo
i9JvfhbjYsVB4iV8ZhSo0LXuVvl9PtAEwbsp97EntbpQpsYY1mZiBz2VGHRzgs6+N6PQ9l47WTuC
/A4jshSgq8hnueRfuiZmTaZlYp2GSCUbIRvQmiEz+K8BGKQ4tFkOlNLQDcN0KqurrLTGfmaAm6Bt
xbQU4Edw3eNjJHd57NCV0OxVsIbyYfySq6pZHOsuHpzSvKUbcxPqusPYYLWFmNH2wz3sioo6Iseh
lqJRi6SrnyPltq7pSvfNKYAk1wT8U8VEoc/eTyrK18GSzmLFHRi43MkrDRP0JGWnVbgBOcssrRBv
SE7qG8rILapq8OY6lyTG2ap2mpIzZk+v2MN/WrYK5w7x/j+9rcXY3TAulHJ7RQTEULnTR46P206l
/upjk3AQduMcyrMybuRmYo5BSxnk4QEnP5XDbLHwGd9HnF8RNMiohO25zNfGdU7Yl0Fa1DyNS7dK
pBZbIWpVtiT5FYlIbY9twYDFaf6Cikmfm6AQuCKpdtmMOZt2lMVC8Ive7jasvBpMI5hJmzOfaRxn
S1X9Huiu4IHOfAL7CGK3hR07q61MFqc+fuIYlOqpgH3PfRbkRRNcdJiQbBLtdBhOTpa2HXTGswI1
i6VzeUDsz2nI4iVqtQfio5x+zWPuvESM/SZ4XtvABujnAYTgs4DSUnjTThfpqwwgQeXJo2kzdRAT
99KImHZXUGCH36BtOiFzUkDkCYrfr+UiQ4MOI+GRZ8UZKbOx6r8jD+nMuOG7ajYmtv+2LN1iA6Q/
z/vgafg/PSrHSNHBNJXi8rFZv8pVcwbcPqjsZx+YfjaB7bBKehqbTq5gq9maeyVde/f8xZia9d6G
tyiNJpINZZhzAycbrAfY68uOXa99yO/MOYX+e0gGswnqlBGp8IvXdvPZLe/phMloB5YuJNgx5t7a
Oal+QTPisfQ5cEnS98PnVmyXWICwZmiwLxy0ef87Zklh/3ggnn9zWey1FVOrexH4qYFhNY6uZMGY
XWDrfRt7wWtzGCUzZUdOYmmm4Xvuu6fc6PzOrseRpD0qg9JYwXuujsSqVeTfnoraWGgAWc+Ovw84
TxGUkF+Ff4bxIeoJXrJoVEXvl23fzCwlYNldc5iwppKmv+TkgHwmJhotpt0vtX118upouABf5Tkc
pIi8IPhiU1+cAw0WKDV7uRN3ZTOd9RPlEhU8dp5SGQ1FFU8ZhCS8lzFGP7h+T7HigpT3Va/c/DQ/
WSQnqznShabu5ML5QtW7QelA+n38ntxZ45PzyspqTtt7AolOiPgYewCvyDWZ0fug17HmO2Um/LHU
myMT9wwffmDrSiFfT/pOnSVGo3aQJnZFsv/mv3d0dP0YC4fRPuLgZkskDRJhw/A7lwb8TKk89f1R
AmVsBmhCNBqFLlTzspEXae0EHdv5dCqf3bPPxF9mvvEBRHur3ml0pfJJz2Q9tJwNaSou76hrElLF
vU/jLJr1xsZf50DEtiK/M3aiyulrjcUW2FctolDtb/EykN9aKbxGD38kmKqs19lDvc4/pcmhH8wo
tlvao8vKEewtH/v23PdqkzTndIZKvZO5oFgivumnilGBFHCTjyHWZIau5M1QCWfKaTq+z8FNoG3m
/rFcJqi+LGa+rIUgsH0Om7tNxkar8GeuOvOcfcltrhZgawkLCt8dDyk3HyMFI0cvUcfU6KLdj3r0
NGzn/aH65hraDmo0ehTv11IpwXZt3UDm1J5B5XVA6G85M2ePOpudSYXEHrKL2TbwEU51ERH+SteK
iaPPGwc4Nbzo79+3kbVF/cJJJER/bKGLNPS8hiUUlj9C+Qd7d//qyOQiJRPuyIeKeIAY+/U3fVND
SEle29SHP9lg9c4l5W3jpVq7DTs0Wu+9xet8kiN/I2/wtLqaeJokBF+UHkq7s4ixqe18arbvglTY
rIMb0mY+8QL5UtP8XPCriWNAWMy1wvGV5bhqYt9RVmSgz/nsnu8Xq9vNdxYgP5LnU/9zYqKwfhgb
J/RyAwxp5shHI0QCQzSfC/EstrDvoqhS53eTW8b9Q4JzR6FL7/MSHmDAL9yUlHlTEdvGMORGn6Oi
yLYUXsrzRI/S8rr/VQY+i7gx/iwfZdWlOSZqa0G8J8d3EDoB7nAxmAndj5gVTsIupYYpatUnZETi
dv2P22sXzBnXpdsGWXMXhZGg30fwZfGWFIwqj/ZP1aZkO+Ci/Ke51VD8Y+J0bimyLlMI+2i62INq
kwwI2DOc8wzVwILMnnHi28nYw4wxeH22rayDCUI6m+rKQdg6K5HCqMvJ7XnctXHd7/wktPdth5zF
MCUD3bD8FFE3jy8EA8AVlZEHkcKfoDpRjj1V/aDX4lEtEAdcUeJgJxbFwf39se7ZphWDhKuXIwbw
YieRmU6M7WK2cwqjsWIVmfrI3n+tGIms702D0wxtZk6KQTDJEMR8IfiFTBK9Gqe2LMqx3xZlRk2a
f8EIDM2/XjZLIuM5eHpMbh/bIofoQbgeYr9H/KBgI00zPl57lZRXCiPwFSNa/rlWyfwsLHNQTmDT
faeOjfWSgGbqeOmWY6ygZxwpwfb0LtWRh6dRszZXBaY9rsmN29Toc8lWzmUS0r+52Bzspt5WNUti
gTCQnj15mBx3+SUqF1RB82/siYRO0lsTisqyZxLXNUas/MbQPExoBVuDmM+yNSR3TnEyeJh7vc3W
HdYfcK5xEqxav3ZCravTyCtSh5vTe8OBucVmIjHdDmaDlnTPGEbFaNP1mZnx9wy52/rtGW08S+NS
UM7TFBKIiMrtONrbNdOEd5JeGBKvQKty+LpfWVPar0gJ/n9q3nh/iEkzq5p5YbNa8o3lbhNEiAid
Hax3HBelkPvPOo4LrIz3YnFTy48YL2gBiCCZ969H3kTqXjhXMothg/MabWZo8K3VOREu4y0+tH4E
ajVT/QtGU1He98rfrU7jppxV4GwG0Ai7ymbklZCHMju9DarA6pcy/Pew2+3bpIdRuXvFZ70rEQ02
5BzGfbrK5IkQ5//h8/1D+JFms934XtSGP/Y3k+PMCdKG9JxasI2+hbJIXSxO9/kuYjuyKkcc7yqh
awggzZyXT9RBuaWb1IYhgdFl6/zEeWzzQTv/42Y4YQQ4YMv1ys2iKrQS5xAgSEdbNUdLRbZoWoLE
uwM7tmwaUapuRvgHywvMUMsQAK91jXDDlCdzEr4OQu2QUDp+usVTEGUctpL/kS0T+TVx/cTmB5OF
EVkIlrhXb8j9GkzD5Xcs1p0p6rTHW0NIKGnE5TeUHBog8PLNRs2bKEC7Knady6oK/8gjHup1RdG4
flDyMCmmT4zwM6wfwUVf88Tp0wo37Ta85v0O3Pvc4LODrj0M5m9Fp77k3yFqxnsmtNDDbkPIkBAT
GA2N6Sm3goohmYeNrw6K3IwEkhoynI3Pd5EC3yelg0HvHmJL18a4NZPnqeSY4uXAxViTwgCYctdk
ixVVCgI9uAuzGykAa1BZi5yCEF+S9pk63RePwD6MzT+QmkZK6Q2CnPZax8Nwn+0FBkQtCYHGiwwE
cl+8J8oKqUNdOdkiDQV4HM74x5Y2+uQCDNsDVFQg4aj4i5t2/7Ile8Lk7EnC8vE4kH3s2VKTJO5T
/fZcxlh49fvwwyfNYyqwxm0+8Hs3GcuHBGUwIMx1b0b4VjkoFzuYwDyvCsyPjGa1QcJOdgN9z5pj
TbDv7Bo8t38dT0HyFA9y/0kMh19lqgohuqNMM6659AMQ/TJd6LJk+oyj8g21q/XLKJxE3A5XoMbE
IRVt+Qtf2c8hM3/xswqdW1v7wMf9e8legtyN4KVNuwFPy+5T+l/5AlUeIc3DeeollAOr9bNI8+xY
FmXSuaE6Z8bbWUjjrc2kqHY9yiUJsQKX+SCpWeaVKuSp1jNFvSszs2VvKryLUEGYuJpUetnDV7lT
vgVGvDOLY6vTxyoGhv4uuYDlNUt20eHluXA5qEhw1BhGPy5On3tRraT36kO0o8Rqg3Cm8YJE4xh8
xjAcpTX1BNcIcUP/q9F+1jcN2KOGO+0BnmitTjUX0EHtDy1b/JYgQ/LUdZv+rlV9hwMkTXBVsZ/V
VzvhaH4IQpZ3ycfFvr7NiNj9Cqwq/coil/wANYGO8E7M4C18XfSdQ8U3LE/n0L58VGuOzyg7yd1m
AkKE9ERuOKL/xv6n4gktfeICsPNB1gN2A6DqUTMcM85ub+sYqvIaxp//2mR2sfdXkQ4276RTM9gC
0zzqFJN7V3YRd1V1MsCHDG+wlwqqtvSKCFsi0g5gYle69ljja3NAnMGHKjKvvqG/MH+k988B3AHa
W6Ue7iJB6RT7/+orC5Hsz7q4DcnlAzvuCQBNjyX8QLJ6eBDLxh4d4JzCxhy9Nd5mF2/ChTlwNY3k
XZ0z0qLXYKGvd3WjYcdxReRJl8K+9BA6PVHzV8oNgu5ZhTueyvsy2kADqdQbNntievvRwzi7piOK
V/PnjW43FGeAZMek6WCdHef1isBxCfIHlyblWsi1BYtfyPYQDg8EaFvETibU/iYYAjWail8hrZT3
sMi0FDY76cWtKe9EqKDPwNQxRcqHfw76/QLbLTSrmdlznnwUyewALOulzFp5keWMHfme91n7GGoD
eHFACYqkHY80B02lwelRW4ktIhrqkNBkjWMWjjceBvEYM/0JnbKzIMmWy0wyadc0LfCQ4L/GRZvU
VuawhxEOA9ndWsOhHp38j6vHmQAPF1CqiuAgG8c4W84MmDWAF8vmu3nYlDhXRoDxhz9gEYp+4M1B
2QdfSVY/dO4mT7fiw+xIvKnaJbNQvSx4Y6hlmuluHL/O8am9/w/ysIP2HZikAYqbSQNleF5otHV8
bSJUSFlxnJSWe9HBToGERhTgIAMWDGprXQrhE/FwzeZ7zIr85QW6dEaICDjAoJmViULuGIs0/dNx
/RcS2+0KA/DvpukYHgd3GqiueXgrtkLI7bd+BAkPVmJykR16JUbl6M0pWpY0MpymBjdXuVkkjp59
bmodFFHq1maQcvqaEWJeS4UPvz8WlVvC9lLjN7+tmCro9v8aC2OYkKJqIkM+NDF9Dih/Nb9Sv6AC
7WxvmI9tmEqU7/MzPLnan5KLh+JrJ52rY6OON9hI9GqfuuWZe+bUSo01e56QTC9WzqP+7/5XWG8t
9iksFGKbFCVM1QEVQjUJR2fHc6yTWDqFxHZZVDYYd+C03D33o0+7T6mxwXFKy/ZncCOpqjJBG86C
q7c1DNsoizA1c6h6sjV2IbclS9bO6j40NGfJiXRqHr14Z+/j9a6e1ojuu2g34kVVLXES7cHLf4zt
uy60+M2QS31HmMslnBmGMcZftgurTaLfSZBNouAXx0We3o6byE9gd0qPIuLjA2fnWlkX39VGChCk
boUL1JTWF+R2ZlGeKwx1yU19hyOMg5vAX0/qw3PSe5gIf1EQErjmnhXaQHih2dqtzBnSRm+IJBTf
eXEzGaB8at5W2Ag74BrbnMa0yGutYq2Iwd25+/tDHO9Bhsu13VlfLGeeaptQiCDufczY/le/Ul2h
3e+hfLV8NnVlGuNy6phocj+3BX/2rxfAwv4PvKzxAvvGXNT0bzJL580hEyIaYmtHvp8l+r7AIwzL
JP9pbBpDz5fds4yNJyF5u+pBoQOpCo0nOjsbpwsGrZU7TnLekMNcA95MMf52OZ1st9M1A0G1uDzS
dOTw63rxS3zKpsDqBMXEMqmmXTeNOcuDJ2vj0igyqMfuA/i8PKAMT0eQ/GtXdnRD2oOHXJfG9JoL
EeJlg3iw4A8I0eNyxJ8rL3ni1wz2BaDeHpo9BRn8xiZizX2+9eSYEKEplM2AGbUl+u2CIqtjsVP+
0Vk1v2sOXgJNLPLDOaIyljQc13Tu3zpj27TvylB7ZXB5Q46/F8MUt4toO8oXlxckVIBsHI99utoI
jZaI0b3oVp8IhjqGzn6vgoiQSYR2jBGC954sUrGyUAgFx1O4lFpChWzbhR1woUHymA2T0QZ1S9XT
8LaM3tokehdCP/QB+04a+5ZqkQ576qZamgmPuxyGg3oamZ844u/SvCe+58JfVcB3/BIGD7LdxFG+
d+ER1BgYQWROOTOAyigCgh3PoCVkSamgjL1ZexBDGLiINAi3d9897gdgYsBmF4kGDBKKy6cEtqO9
I4Nczbp01TORmQF6sCRw2S/UAwfI5NBrAXuI9ZF8V4SZUu+MBa+V0Bnwa18rRFChC7g3NCoI+Bp4
JWjtE/zVEkwH5X4k9AAYQ935DtNb4FVBJBX+FmdDM5yixzfOJIZc5F7cVwCv2x7wwN5aHFr9fqDT
rMS8QvixnCpENTJLm7iuxgJxq4EI/MU+hfiYIz1+NHasSFU4qJnx0fhDbUE6MrYm6KkFvhrjSl6U
oGh/MktMqlkbVzCZctT9JPC2DEQu4zgIV47Vv8DogzdTWlfDPXBCiCoSAvsXv8YCbcvjO8d9WM3n
AbVjKnOYoY1GOOREtpVPHGqtmMqiO5t3cGOPshtRbtd+5ZyQDe9lYFNWh080LnjqJXqV6DbG5vXV
4hlz43AN9+pOE5qnTkw7cPqLD8DVyEe46sCYx6IjvxnYzsYoawgL3KP8+SGRsUHL//xI4qIMcd4C
mFeD5DQqIprOAcJXUPToscAbdDY3UtSEIOKusVhAORA1Rw/yh7bpfqr9zJ8pzjj3q1ownd9PMAlI
kLB4rFAWBnDod7Jrx4/kEjdwmD0zcY3WLoUrBr2Er6ebew1xPLnhfMq/ZPGmpBOLlncJ9OtPsy/7
c8MM9ftJRQFQAEgXlOoEEM8TVp8LY8ft8hOJRAqDbVpu9F6BavBZej8Xx5Jwb8uXMurYr1Qnrm9O
GbJDMmI/WHOO9/Vf0gsRHTVBKfDVVZwtdog/KgQVpUT+QqNryE4psKxogfiRUpJM09l1W1tYLEia
fMqKMljijg41nI/cnaRS9OSBuss+tmme+6j5AFwU6NeXd9HyFDoqL+LXJPXL4qB4fJlx3sRYLIHU
VgfNm6hbzZZd7334BjDYK6qD+lkfEDzUHDZ9zbpJhzU7ukT5SdjPh0bybAMq75+UgFGrHN0ctBsv
oK0/ioixCccu4y3orzPiMFACHieTf2rGMgY0tKsBVtbwbNB5gTaVWXL+MpUlkG18dMEpNrOynwF7
en410HAvP3wuRiKhHKv46xFX4W/mIPH1JcItw99oiaNmh3KKXeBVcxndt0gTZ273Bc5bJ+baoAf5
3lFJrRhQm2veczZF5bBEx+Owa9fkEeib1IifQx9fzdorZ4tGGduBWKcRxjUWEktzHJRUSbLZjYaM
Xxelew4VGEFejbrWt5Potz6gU84iGjgB2dbqqphqWcBeuPQIjnWqeW7KhGvRWZDxDT4Bq8sqPZa/
0l9OGmhIBxZ+wNnt7+4YsxaEPQZBSedjHzgnH2vVcBouxMDC8n9rUcmyvVXYMbRqcXxkM6htcjhb
MluY9oWhwGx799hTDR8IghofkdKh+AziiektSRVB/mkhk3SOyZIpu8PMPqVTKvI3oCFcPDbjDBIf
bM4U2T8FAGWQzI9nRCggv/D/jEjBGzFDsp5yMfsV6DFfBsNTG+KDMON9xcu2rzHGr6VJGCR8yAw8
yyXb4m60KX6LfJQdKwdwKpiZTrm4AtfdNENZpH7bndOvIslAmDiIlmcTPmo3zk7K8WEaYTAvL9b1
sD9C2n1McWbw1AI2gCmcqB1Qgw5qG9Wf6+51MXRjzEWd8zMi4cQdwN0kP36yu18/JQyLrt5QUP61
/N0OMpOCShtlVyXkxe+qOSlIXQ+HjtDITceQhgKnk6H7eiaFF/bRyfc7Di7H9NmnjFfFC5XFuXgb
qmhR2tQxJT1zp5sTCpjgYm3e8He5tfCNLBbiY1hSjux0qM231/3GERZNa+3vqpAjEiN7Modp6Raa
YPU5ALjEltH7WMoJ0iYJCcGiZXcbjJbAZjmZNmR9zpPy3+HjE0O4y50RLd/SFOjuHzfCF2niNPfc
sP3h1OFVq0MDLXMkby8lYjxHvGP1lW9orVISBzYn2j7Pnc4dDOdo3oREyiYvUYpT61a657dphSP7
g/0dtHewN8K8no++lWyBFHbRnAcSfFdAocKC6Q3hoznnYH948Mkv7vxXKFehVHsYP5+uImWlX0LV
gn+si3kFBQYFodHwhjIlXbvWqeO/o/UyZrtVHqi7ts8VEKA+Rs0Qh4b9dG/+4uG42KX/2k2VbqSD
kywIGMst+J0hv71ldtFYS+Y/Nfof7NU4LneXh6GjWGYbbXhDx/FqLpMLh78x5mZASn6WH+ooVnmh
QipcdLRUSrrG5TbMszUZ4qEOaY5rIn73lf58fk+YUtEbtRsyUQjBT5TT8SNX2YabeOGvcbRe8DCC
eLvTweLWVCXejCGCFMbaWKRw85/eKqYZ3zK7siXi89ZaPfC/15GTtxwZGNefLsdxpXI2UETRmI8Y
icDg+XHMTsTtrBav8dPHHUFQSv2f9kuBv6XtBbfCQrLvCt1mFFVd/AbWvpYPzCPWlNDWcshPGSAK
LJlAM+jyP0W+05foKlcTfCalnlfmaq6WlOsG0wbxDrLawvdTpU7Kls2xqZicRtOVAq1Aba93OB28
LUAXZ4FweQGWKSmML9PM0DUM4sekiGeiM9EnEmnTZWze9EnQeoKzO+XEX3/EjRGpCQnpvi/THkd+
yppho0m3UCqVie8cTDVIsMJXtcCVgewdN8DeJUBsGVdAzdPYs/+YFHRqQdDdIzmw0NQo4vXP2Ws8
u44qc17xE7tpNgzmtJwpVu4u2r6xvbLV5zwe5mcWvjM1ShG2AwdZPxLJT5jkMmshbLdEKLTqKZq2
8rX02bnVBrAjMkDln7CI6LbKgbxKexfr2w1If4MLJuz+QoonwlpaI2j/GmSTZheR2ChM1KcxT9tC
q85bKuDlRd+vuftLLnfZwD9rqsNJ5wfSN/PElx59l63jpirMJvimj1mRdDhFoT9lGpAXzIvyNAtS
+1s3ZdrkWO1pF9XcG3PJDpfLfS+LtxCnRdK1Lb++hpwcbKYy41kMt0llZp+bYK0YxXahASO8vQga
FT0D4sbfjHDtvXLskQtpB6Jyr0XzF8YS/Lczckm7ilqvwlxFs+ykFkRERLFy/Ze0+oMg6jHZV6fr
VYhRFdRiR2aT8rbXylR0v4LLZt1Mq8jB2BRB4kz24d1DhHPAkgOXroXZjqsP32WHm1cnMfb8UK7P
ywpEYLhzcvxEA/Dxbt1dSW+BmQ4iNfoAdwOCI5z0xt+aYIKMq9OU/PlikZZ39nLDt7ZRusJ+XhOr
amwm7+wdZqMUCI7FVlS196oumSOk7i1l/X1AEsBWjOw9RXBljXTek4Co1DsyRn3U8EWFvVxCANqu
KNWnkqu+56dJkRBwOJ9+wdgeBLFmNkWrHJ4VF4CfNOvYkMZHQ8L19YNItWmHlUjMjxm/+0aII9HG
+8EMI0XH+IeRVVA23GLxVn1pOErnLmLFKlMRDYnp8/2wukOA3Yj2Dm+uTKKAsH8BaOJYHOWw/B13
YT1nIBlXVxEtBUOW9worZFcy5+JYDNrHRgRDEywYEviQz2BPgzUKZtcvOh02Shhmi+2TjY0fhyHS
rXxtQS25BLsQw/J8yaDQ9T99Ay6GFSKKredayZ3bFQum6acugoVxtOPaKnZT4F+8WeMrMVb5/jYF
IorCXgMraoOjZR0oUY0E8qTthH8gFCKS5i4+fHtfQQlYTzj1nbFgNKXVVSnGnb8BIzs7NTYPxB5V
xi9XE9DSHHx4NVSAhSqVgcIh4rA914EFoNMQoWvfSKbx0P8fy4bDcttLnOZXRED79TjTiChKQyBH
8/iDPHOwPrO5yzFqZVHJ+Pt+d6/N6bd3JjX29YiHIRFMoON+CVQsjs6tRDIRYkFpVZ0aofxSzfqp
A19T8Adr7JEH6ugbcCwVO7/LrJ3ZxNYNr0WtmiFGP803009X2rvFO2HHAr4hcVBhCF7w5V5Z3brD
kC7RJM9Bq5CKPoGGAexbGaJ+p+nmVcLuFEiRpHmcTS+q7OPLJLsbnm21Czx17wFUl7PouACT4BAg
e3MERzXOLuf+FnXYRfP8/aEQJEHKKnRL5Zs/gMp/T9+UgSUSBU/S7TGLveJL1VrhzhEJUY3UiTGj
Fm/YPWKf1i41m6shh2sq2HrWlspaHYfxDQtCzLNH32aQRdKf/KeM5agOnpW0Fh5krneSKE6L30CH
Kj9f+NuThSEjvK/cg8KQP92fipnSX0dC6qsrJ5XXC7+v2d8CWkJBueqDvFPGjnok9DnI8mbD+yzl
RZKH7z+WhlmigSg0nvecDVewcyh5+oZNnmieici/Bs5fEWk4oq96VA8S/0o2gwHpJSRGDm/mLgdq
qxDFstfBUYxPlA63bO0//9dHNn30sqrfYAInoCTUXqyFzAuNIrFZ2cnMjpBO5JcwMB492iJjMcHw
UwYa8K9MvGhoYd+3LMwVLvUL/qamBMrwA3Vup5rvEhz0c8s2+sE/aIhtusKLBFOlwz55emwmvUVU
7Jh4xsVavSNUeqGDrZT/y6lun9L7oSWhOcq4SNMWSMUGzgwU5a/uZit/AQYZTbq+b+etgeo/xj8F
VWWt2rJPGtlQqV0Lishfz6qQd3I9DbyFP/3UvE3yGc7u0AkPI7o3QpqjOzzc3Q9ps4HN9cEGbcmF
nncvRoS9xi4qKeeu/gjVSc+xxRQUJeO0qSHhL1fEWE8AVNtjq/502tqWHbmpt3PjYqSZDAR5h2Ea
sh16MSI1UEPNZYVz7EHdcipGwBfntHAw+kbE0+u01SycMnJbGCJXCb7/2e5EcjOXynoXqHe+QydL
rAaglR0/tPh6h/cDba/M/ISFKjYFky931jton/RCjyUhauEh41RSgY2pvUa0gYKAcCeDYSz+6Q6s
wLNloYVRRalPOi+au+1jve/wmIyq5426OXBqCsXR4ieXgngfU0glDi9GlhR+5hK4hBdk4O/kjCrU
2txuC1m3DFLE7WTv/4TYQ2tu9T44Oy1+cgFOM5wpvWO+jViv2qV4YjPsfywCkFDQitR+6AwRvpnu
EVlFgDzZoXQR4qZ8H1mRLjwBHdMVEpyS2XX4M/L6p08aI8FYEXfWqTzDahDhA4BtMPkbJcMfNwf9
coWnPZrGwy2O8DHOlZ7hY9BdjsVSOHWaPGyuaDmKt6w9MVZJ4Q/QM+hARcALqeuU+kmcBvJ89Owg
g24jkdsPxo+Bw+yUpU1LTGFNydSEO9KA/pRnUmBNC66diLDy+mxQRCItq+SQOKJpy7Pdp78x94S3
qPCx+vba+eVoJXLDc5qKRLp51+zW7SE1vfEPiIGISiSRXgFnK5xsDCPi8pV7qS9eJCZtJyn5jxZk
KBHSaJnu5hU0aZoj/NiuWpi7dAwg43W4t8n8CAor7vAf4cTztCdJ57FlgShmJIRjpWNxSOKPwGpF
X7eQpA7+BHrnAbVNUUu8wjeVtrirbhV+EPZ2dhDoHSkuFGmmpOBjMEwMPwDJlIn/8+m0j/5bY8wY
PHH4X1T1YRFTe3NsH4/NDrdIQ0r+cJdGYelf7AqGM95ROfrqpfFI7HbEemMbjUtV5VE8cxo3UoUd
0c2+czdpmDlkMMf3TI4pt/GkxqtgKsOIvHnZbLA9pyEZa46D1t58jQNeMhATc/BhnWh7MYNwOR74
mfBPFNjnIwF/nworhsOcA5LI/4pL12kiIs7qjeVE/M46idliAfDCSdQsv0dDnF4olGvd2f9UpgVV
JyndelxhIfdI4YCWtMVAqy9aEtY/0LP6YNWgqk1xOY0iUCv6DGEZc2w8v8sRZWcC19i5MJ9CL5b1
BJkHkM4phI7xY6df7T0KYfwJkaXGjvb6WwjV1IesMIUt7bnWOmoYiMZy3jtaavH3GFEFb0tQpQQQ
NqiZs4/cLpYilAAGlgcbePKSrBMexoZKj8YMdxWp9FLxWeG3/hhKESZZZY5cHWAvPzDZaPVgItk5
yfE145cMPxld+VVzykX5ocBy/Kuq3bhHKNHETEFwQT4lwZ4Aad5fAOUK7kpQ1qOjV3qL48C2WTaV
VMTciQWomllHMfbGyJRHq/80ZO03HGbNsr0hPMqigdzg9qVlBfRd/vd/bKrpnSXCjI51AU7qlnee
Zm2MRrKWm4Sn7+KHeQLz9Bad/TqPEjSX0X08aj7C8g9SYuZumnV/qafjEQ7HCHFLalVIfAYS6kuj
Tj0LTvi7J659I7rTiQ78cWAQ843syMy+cQ8yOoWcVp0i41glGqq26anpUFWsQE+eU2EJQhOgapEl
aNOsoGjIC0YOkYRELH7TzikuVNTSC5D3k2fMTjMJ55GpD15FKBzoaJT70xfqUDF1cNCoD99lt6BV
zioW6m3MlJdX/UKGsavhd+ttxf/XQ3i+dEhp9dw75ArJX/33qpH6mi0/oKYDDpCX33DHs6OyviU/
ryNCn8wP/TZqZZjy5PAFwjTFTZtApBsHNVoAnc6MXBXChet17197RTYbl0opw6yoc2n/0eKfja8X
AnHkUHvQeaUWl+EnQ4WOFj4Q1s3V6z6nTytYXNuciB21QWkiK2ZuGpPGHec/o0GFjPUwzYnidymS
H5n/pNl0QXP+JmTQA8wGICWliXTw3++ZVu/bSfmp0lMy22AFOW+wIQxMeLCFQQUk87V2EG0AdBeL
VER2/MpfAmoiK/JRGE1X5943uJzhy4lq3/4185H9zwfNje/IEAEySfljLEfVph+x7u9Yao/pxcHJ
E9HkJAgCmQlODb4bGb0PgNjZIG9YQwtI5K9beQYcwM6NSogkKqMGVCGRY8pMZ5cUzbVpo2yqRGe5
qISNa9NnK6YkeLnxY3MGoRJDp6XSQ1Ul4t9tGdnxTY5yxjxdnc8WOROsYfXFq1jK9L37moKbs0T3
aDJOUBMvI9qXwOeR63j3D4gaF6YhwIZTd8WGO0QC6MSIpokc+IlJkkig3k//yQ1cn1/Ty9OF/Fs7
RnWPFyW5OpJOLT/MliBNeQVbkpQweF+OrfaNegxvg+yVu9waQ0EECZ0wO4C/DMBV21HIpj0xauhw
WC+my+xFXsNH+NGgO3OFzLFHd2sSIPsIWqCniSOfqHqx8nlNaMEjUrfwvgJ7nmOzrwV0vfHbpIeG
LcCEWWWGBimc4xO2UqVE3SWXitNQk/nS1rkJ/Jcw/iCY04a9nWvp2xxQjrr9zJ96HWTL29DY8Ztf
AHfqdNZ+4ijlbQx+chrk77qQnQb0bvhyTO7VU1a6J45A3WPjtYMGZP6hOHuQ0lIzL4ZVcQqYzuF6
tPxeq0iOtwwg85lzLiErHpQOZ4u64cnpdy7V51DRtRjJCQgzbGNja21lJzVkXMSDuR7u77q32sOn
cFSpgCBfzAcbfgmlfMKS+5OZ/kKNf5E3PgBMo6js3AWTolybAMNWbWMyShUWG3OiqdKD+7GBeKmj
eLcxNbMw5uFK44BMfuZWi8HK/TZXeSED8ErCqnSI/r2bUGDyf679J29E4zqQcxOxyWsDEbN5cXyk
H0uriHG5wBgKvU53tA/G6lgGHUhIomUOHqzMeXZT7/RwxsFX1sbhzSkO3XogVzeVJXiUsm7gEgcC
PyKk8AVDjx/a6vcsrMZC2oq/OKukIqCK7DrpekAZhDxj4lwP8yB3SowtTkGkYHkunjCNg/L00Isv
BC4BmwvLZbyi1UqnAvn90MTBklLutj24w4f2A91XS7ATXnrVPDRbKKq9cKmTKWSIjxlm0ggecn++
P4pA7NmErZ5CZzlDOeaL7BFon0PQSVwn1veCxPpz2J2s/3s/VpeasHQSp/LAXe9CHOR4HOZlHZy+
qOUwFNOsJPX7WW9nltSqOtvouvAhbOUPEbfbrWOChVDB/BJmxKtYRhc+RVr1WQFx6IsUwVsQJR98
uymGOHd2wOgsB52slynzAlHJdHRfLFcIbi418IT2NyM9vBwt7WGcXfIlj3JN+khR2UONv9i0i9H4
lc3EJMBW986FrwNEejM6nJhdc9mhjXFBTJ2YP7mhbjrHzCF2fY30J5xK8H81MYGULfqpkNy/yw98
h/EFWugqCLWWUpkVfICrU7HpLA9HsX2aunscyxCOonzUQlxXbpveJ2VBBOiKXZWvDOVNBE08nTh6
RXCyTSQZsL3B0mwqvjkDvsNGwgRMu0TMgveJ9DsVaZyNUJ+hSUEU5K4/vt3Jde5FlqmrJttE7gXd
beS4ilhsg89cNbxngsdjMhhJLHrajhcr5FW6GfBO0qPgYcP0NfnUFCWUTzczKUv/FugbykOIGbuK
+UFRHzat8tdY7sPaovQmble87vyL15HPMX6UzfTM8X6wN1FYWVxIN47NlHRXGVt3MPWgm1jhLcOS
Ah2aAnXeszOiYVOWYyhh3fN8i5YgGKL+79Q2KRjwgKUzH7eTYTrjqHad+zB/wvPRUGxsZbk/7OYH
ct1xrC+QZSsto0PzbwW/eSnQ2MKcYdrsaf/mbM3YA8+tXn3FicxEOgMk8VzNPDCWMBV62VAhY8Un
/zPN5Np8TK40QXvQ0ludx2qn8/oMAlb/vXSbsahtP7v9Irfi7FWTCQPTZFNFySlfIQ3PEfsPw70n
UtIe0yNyMTG01uqLIwJ9UjBLhLDg4+zbvRZ9rr3BgQzvn+CYy2UsoyBzXavHqbN63cU+Jg9Zg1e+
dDddoO90DqSccPcNk6ZY9Zw22AqebSwJ4rlSuTaK9A2EiOfjdBt0sFKW7h5y+ovbaAxbOnqF8mB0
rQO0qZczjmsTQiOIRcAcNUfVbXMp8VZm7nDfXeOivn5LbPR51QXN/P82E6NSuD9h6G/kPIKd577F
oUU1GI5OAmn/Fvr2koPMedhSi8ceOueN/yCMS17yicuFVN7J3zu1nbx8KGcxdLLKm0/OYx2WVlrl
H1C/OgeBKG6HCdSXGntLXnnWl8Hq5Dq9bmQIBflyZD4De3/UZIkwvE2jTX330DyM4PI/cBnsfvgg
ETQ3k5duT9kxWDJo3CewzqJqBbH5YNft78HJIEfXnyvYFFcDLo9pypAXPvFCuHLSdxj3YRSfpmQO
ItO6ChP48UVtgDG2sAU+duGxNei6frHpdwwrkG1w8MuXka5qa2nLRT7N8IYE7YHxqFreeTjlJrVr
Go9HnWNWjZpp0ADrmVcbadbh13EMvLogONc0Vb+xJnKSlrGXMFut/z0M8zVwrccyaNp206hSO9n1
3oM+pQMVeU9QHVXva4IPoFfB9dxiUPNTb7fWfWn2xkP1J5v0DIRGffwdKUKihx/NPOFybKtja+p5
1TRP0oQDTwEeDFqT4ZSzRwQ39azYK6yUCTviLGrVbOWVqxxJymaPU+HATRJ6wf2soNa2UsqbQV+g
S9DynxsP8p4fPfb8tfO7CFCd7r2YuzMBPc8eI40Rcn3rO3fvm52cA7h7Jdfk57AyN/6V6d8nIKg1
BV584SufN0bHtkBNbHFZH+ieoW1I/GoGufP0uPXnV8vmkrmHVPRzwNe3czpziMlLCszdpNu+FW7K
/DF+4PtyogQ1ajIFdhNxYy2IrG53YrEbMXpj5z+Zhs/KCvLHUaqeXWh7RIa39lSTJN7e4iqA6FSm
MA3MvjXc1QDO6wg1JB3Es6/K7Yfiv3D81pNqDEGazxS6h8ETDzOj5hk913qE6FjxsIc/TzVn3Bgm
HqTcf8HjOrMOIhipwM8XhqDLA6FkjRQuE3vIyeD1Vmd47T365eh5lblBCTNd8K2vpTki5YZv/zGb
GyDvEqpSu7Nqh084sIgGzWI7484cuzLm5Zrk1yEbQQ10EiLA8xBliq+LnfkVvStK4vftA95sXg0+
dqRCVu0NYm0jSMmWazQl8Y7g7AjyzTkGyaLMg8oHhXnbZ1xeoSYTemjAfdqirHnXehcJjq0XVFem
5rtJJ9X8eHGOJ+SPGMuPqfeAsOiXz01mS0LzWw5XBZfArPIyfulvkPfE0nRtIhpn/zG+xv0tzHdW
TMD4LLAjb4gJs+FthMq6sPDOBswDlZ+yWZgFSm9cP1cWOitEiOyI7nDPfgRg9bS7ABOHGtnQZUxD
eHPm1DD01w//Z1Slykm1PnyuF4zBQ6qtYr/0yN4syAWifS67UGmrcncJ5YnVL9NOTFDywqnddSc2
bhrPgxxErYQpjk07O//hQdysG2ynRBjyLyUvNbxI67I2osPE4Rrzy9usoh//sPniQju5O3yEIIZq
rB4rRKqd2j8PS0oqA+do/sjzlcv/g2IOPHtSjK7p3gIMgGYD4UcvEDYJPEIuq6NFkrs4di+QIve8
Agal9NLQnkBrwR0PFnXKpc8iiqtGR1tLG/N2RqJU7eABAI+xwhkJaVjdeLPrNHUvI96h9dR/J5Bv
R20ePtuwO/SMWyn4la/H+W5IitCKW3WHvXdj6TUXz7humGRopDKuEs93mhnuYMpdpGMBDTD13lTE
nFufcsn0Q7eBFleqlm30mUp6vovl3px7p/yg1lfJhpluTD++Izhi9G5of5taMxINRuXdL6eq2qaW
Mip91nnJD3UYfXZ8lZFLs3AeDBCo7FP/FeQverMUOk4DEyq5qKkZ6O8kueTTGp86GjnxEAkVw5XE
9M42wdkVwyM6voGmEbe90MZFCfZqK50XEB6pKiSMAmm3ZJhANHWRveJ6S1FP5F8rVCkYvIw/1hVD
3PcR0h88FreN9zxlhYJyW3u9FqGNJGcoWW3cMitMVoeDay5G4yS5sLdipyhSEuO8S2CMylKHqrPd
vCQLuRme+5kTP6Ceh7GbMder39MhAQLE6elskCjltn62K99yHDKkgHU2d3mA/SYWc1Ttyz62SZBJ
fteHlGEgRKQ1fDGKzwGRNaC5zAHjTsnfKKr47TYHXLtHXIuv/yjWsZf2hOF4wz3Qh9msxumDH49A
KU1mgZptJc9wgUFUr34eDFx9PaW83X4tiUMie1RNhMI+aTAcAqU9+cHZTEWv3Hh5gGC0hQHH4VtK
jA6fExICPT79nlMM2AwXRel8FL/PmwW24JgwTknTs407hwX76kLVzlBxDzHmqxISqE3BEpYe9AIt
FiBh3rXD2aizEKtutWU6mSSnrMn5P+DjQn4RVAoU7RVI+obQwnDJEiLfLb0zw2hxCBpTGRF3n8O2
roe4uRqPJ7RjBNHSXeuoTpvRa22Fm2z3oQgu4v0RVwQgjGQMm0EKk3ZsoDU4jsRfCK1jK/z0WXdc
huBaAUkACMI/ZZycKBJa1gbJ3lXuhA9pschSsakLXtfPVD/CsUtJW4xfrzTrasCyIYF4Kv9PVZvC
bXKt+jvjlSNWpsKvqy/xGhUOrbW97T+EGJPq9rd/7JNBA8M1PuZ++truYFJHJ5wDyCDFC5rq6cBX
2CWRrtXiycSzNfJdFJTUkqHBEfb1m3+yApGRhzxNyUb9XNgJ2VzjbcgbQbbqzULUuZODcF+wtQgD
Ytrgj2ebc0kHeeLEcKRlDJimDyzYwj4+aGB42w0z/Oxui2rp+ykf8VxOfM9qzhSvD/Oxnb1ahKBm
dT6G81m3pm6wYJRRUzKTjW24mdmavv5sL8D27aqiSNmstZ8tQtazKCQqItbP2l+55n2XlpUcYykd
CeDP5I4Ta4AnNZz6Yjf/kXg1h3iQyLifRKCmgeuNFhECAk3YRBIwXqbH4lTHPskxtqWcwuK8AymA
vNw682PGQuhwT5683ErzFiuE3ESMYaLqM/x0F+IELP3xIGS3OgSOfgrXVYF11HbHAvrczIvCqPAl
uo60NuiuoQEzb5FRCB25ShR055jiKQK0FcKfFMH7eFxqdkpO04PFmIQzYMOWX8+56kYtIOhZ5R8g
EamKKqLlhmIBqU/EQeGdMp/aNATVkgBRNYiU1Tu24QcegC0TXS/wxyPrnJVJJ+h1G/QImZPB4as8
5wyOqRjyWXbmDJuXoGlhrdHOR+QGJiRO6fsXRK/qDszOqVqKKb8vBVkb8D6PM/WzBTE138Y9EJV6
7yKaZxyRp8o5/Qvswi/gpWR1HBCbzjZIbcGd+6AqOCfxrIVsq/KJvyohHz3W5JZbnCD8ZFsLip9N
ACeUWjW+M1lt2ZXfvO55ojeFR+aoXVS2vNk0W8+hUo2YNsf9uUClLjBrg/+MOUixJBdouaJasWjE
9e+8O1Y1ir1MSxDg4uUWzyipXb2Ms+0h0ZIB64u9D/vhFKEr2AvZ7fZrh5PwmLYGtVuUouDfTjku
1hbmLvmR6j3XHbpFNrew3KhlJnNG04PORfiiMfvU6ouYggYpPG4zotbbNgV9oGRuDV/BwIBrw7qm
+WbzhzqWy/Jc6KQ7OmaM6TFNFvQB8c5OsR3VaQfsVBplR3OIki7B+Kuc7AOl4RUcausO/yhGl580
4sJInn/Ur0sUcFUHabNy9tVTbNu9n8gLAGyHXkdy23wcfG2W7D3GWiI4aPKxdSSSZ2DgMYJm/Bwy
LmVInsLTmQtMrKHWhbrCoaPXq3jhLxXHNIrEQuH98JAqArcY7t1pEYcYfOUvV1CR2cw9Twm5/sCB
buWXLQW8bb0l1O1sIOKo+SrZpw0GYNZUW6IBzYvyO9FIxCIfxoNmQBt3OGeMlgCJnw7WNARO70TG
FLoCrcqcikb7DKim3inMY2O/TnBnWN4xUDt7dLP96GnXqx/YQMikaN03xnUWe8vdyuEsiSJM8Czw
Op8XUd+K7Xn22MvtU92o+Qmqel/R9eni1/QyeYng9XzkXvTAX7jGpQ8+eczmmj1p+l+Q/ql5SOcJ
MvDXWPCHYAHsDGtXXGOlVptjvOMsQ8j7fdK3rBVj3oeMXnCGMdRZO6Q2KhuFpHZerbaliIn1dKTu
IojR/OQcCEN+A995bD+Iu8tESrbTChF5P4jnY6/oXL/5U9vaMXuSViiIjMzwBMA2cmS0qMgzt2S4
b5iX3LzXFKWeNW9TwtNC1rpz4w1q7308CV3B13VDYotNhgFy02UK9ZJTyNLVV+APUE+aqC8JnBiY
XG5Cagzi2ySm5eTpWBGW+LuxlILuNJx3buX7ey39Szhu9A8yHiGIr0TKjU0tcIcmfZJzV+rJHBGc
t9oUIo5bDPCgY0tKarWGZFyaKy+4lMCT255b3sUtypPIrgh13bli4eSMiYG2nK6+XgwbSOJ92dAW
mHC0NCfpomcKWzdPvD/oiyubyLbwX6qe1UhPrr2sCFzElHDhAVjM2+28YubxdGhsGhQete3VuoFB
q1PSXQY8PJnroMlFAfo2ni4Q4dezJXNiiwXcLaRisoTzLtsVHE+SPl+EHfhbeAcDpYIyFvjf0j/E
qhUl4f3owqTNC/A2u1FqWJAsGVSCNyClDuPXDKimp95OW8Tz4KZ26ZkgFNL8W+jGVGMrc6Gkj1Kk
Wp2syuTEwb3q4I9waFztE6bmlUixWuaZbduwv2F6coQB/0JF6qY56BX/c+u0e/15ik44LhO4sF4M
62JpkKnUXJTnepKMFzNz6f0CgYejUSOjivwURiRdj+FgNaLWzvhjhTVqKcLXNCp23FCN0/d4Z0gS
J77Ips8CDmcE771u0dv1VbRF30VryEzt4+UlVPwXM0E91NFETwpNlErH/fBV/gc3HhWoK3oKq0HX
4OFB8y0N4lCHN6mQo8LcLmN0XeBuNHame65sO0ORdiI0TsXP2fkT5vPPImrMxEmM5HR6JPRF/P02
NPZR/Gbm9zDezLi7WAuocR/HUw9rCHaTZTwOkm3gVJct+PkXBrVLzaY3rPCHIaRnxLwl0z3yWzKV
kLdvrhCzHsuqJSot5F+2wDSWIfNd34aNCAfLUuhLGighe1wleMI7tfvg9h/l826VkIty/CDjoJND
0cc4M3Jt050clxUfGPEqiOwiNTvzPXTETGjeCHDStYc6N8bFvbB+9v5mhzspXpxzKdHcdnL78M7S
OaArsc42T+wdYdfGtbeZUBcs0I7jgba9mfXQmFbRe4tpLyOnp8PSUg4BflgKtFtSuywPQQ/go8Pq
TLyGwCs4CV1k0z3LRnCfr+u/n1+Lm6LXLgAdxgew/r0RzRVONSeOAQ4NPlwKhu1Gt8q3oSI0aU07
lBC60qAlknR+4aLzGKAVDzHM8kPWBZNwVSEDPqB9TOjuRBk4yWCTBgbj4/wXeeMeNOSGy59lfodU
8i5m3tPMfNqM27eX8rTMdL4LEoIME6dTvQ8cffjelgM+AScMB3QQkwvyokFmfxzrbTd7w4Zx6hQs
1f6X64I/1SV+jTsU76ZcFbgPOcXjfMbbp4rsfG7g/oV+0bdO6cgSReZ41l+5UWoRvcPOXgfGlm0W
Z7K1AD1Y+RsWmZ/J4GHw0C8GMYYokKwWjuLPc9Bub3A02nzTgd1NRcvdB6hzWADPVpQnlHMvksWV
1zZP1LHT9SVbQToScTDxqtQJoTxGm6NhHbX50UWC+M5pBQ7m520RL/hK76eL+f9qoftEKD6MSxf7
YzQs55c/GcyLYTAwC0gm789VEeCinIAR9Fv/yEUOU2N5uX3OlcjrROcNYNiAtvyjGwTm+KgzEnSR
oFlNjMAO2O8jfu68sdy+ezG857mvY9Uw8yBe6xyaxRKwALmRYMhT+zz+XuBnrTeLEzSl1sexSWRt
akp5eGr+h37+KbxXXuGbcwqLq2RFleccNE34Yqy68aWERm73YS9nsTvHK5pE4eqULeQvH037CyWY
P+GCsCF3fa/HfivZJb9LpD8JnC+nO5ps2ontQecU3Bwyjvr0c5gADFI1x/BPAqG6M5C1kugDMVBp
qXWUDdLpUt3akVM5oHTsciBUHveYklv14+Soqdgkb18aLrEsvh0bUsAUQNET3iURPOBoENskfGf6
198rjR5Q6UC8PFGV35MQNESGddrXc0FW+u5bNnJQ6glwmQF22lVmtN/gBi8VFmtmAj98UwPxXSOQ
8soBKlxVDwV2rPNfqye6ouUa26bO3kNo3ON8Zs8PJTybnlLZLKmTDOrudvKDtB1JQ3i4nES3iX39
TRZ0b3y8L3b9jhtSgQO+0CjGyFRwMwPzBD9rF4LLvLa9fo2U6SnyI/JSplXnbbDGC+Wp9D5pnz5Q
YzXaedXjMtpK9qSawKywTbgeVNqKwrgzvIwBuCSlgmi3jWbTE+VMsC9kK15HWl4ailzCcDfNqXMs
BGoYG91ypCvKVuQDZ6Q+r4FzjHqxPbf4CQ2HXIVD8+NIU9OHGNSNLGe4ccJW/Lq26ZW2FYTXHJ6o
DZofhLsjus1YR5gli7d2XVcn9fKvFmhLd8eGsH2d/2Kq5cI795K0pE/rYqntVXviVA25wQMQbxb8
XIqZZd4oAAy0KTFDande0IP54T0yxAXcqwnA68v/SYx0FO2KVLKW3vL+x4wnilmrede43Du8FSwV
fXOh/6fp6B4y0PKj2cPWNSMyP2RodNtFHve8iem9n7+MQ9UdXKmqBTwsWLaWhlhij88xyDy5Q8a4
ACLecFMW3s07XpjEDusb9nuzTrNqmUGMbMk03YrCJzD9SGe2EkYpI+FRw6v+LCIgrbtU9HW8lj1B
C2CAkoRla6lBhzkjEn3Khe/P6qfSNR42o8SEjJWG5ApCHsVMsvhpLbkIIUk6gOf2BMzQYBhXCRtB
5RyxCdNL7Q4sj57kIAV1ivK/c9iC+/9E79aHdYfQ6klDA0EHxMDIm0cXP8NnKjzxKz5wEuYdU8Te
C8nToKDY7WdAopak7kKfsULQ5a6y+nuql4fKBbOt21D/gY51/4wOO5wgD55LIVMixhO6cZGmlJXu
p8PMNtclD9aKMzrq1+jR2YByTX4wJ1SUovorhAeCjYEv11ORH0Sh6PCVRVowB6asX9KTvcKs/ZjZ
n+EY4Mn/pQIdMXeSa6hCCXWc9z4YFwOzzTGtezwQRrHkljplMy9kZbIf0BccTmKNPTQsjxoROX7j
08ppfeSwoxPXdgdPp8X1jXgUZsSUeJTAikrYaNTRMscCIXk/Fe6oVR19gnuqAhjtcMGvrFLTtpzZ
eQ2PrAK/53kqwe3fQghF3aksd3XKfFs11Q3HAP+7V0VBrIAZ12izdUBLsp3WXJd/UN9CNiAgd6WK
ygMpNjYRNFa9PBLFZiGCY02Ykk1irSfzOyyBMcln9xu/jc/CvvQ5y7WKLcASN/rSxUQQdW1I1cPC
GrWmfPKhIAx4Bxg0ZU0jyDpKj5KBa9RfVg2CCJ3CZN6cpPHJ6MWwGKQx8z2C1RqdfknRh5A/t/XX
PXvYeOrg74Y6xYMuro1UNMk0d3A3dnRrwYwzZAe5OLQVrF2zaEWho2tM3C9B4+p83dAikKM6a9pA
zRrPsbQ7ZXc65RjhuCI9s2wVdHu8tlVV9xqfit8VCttrNhB5Geht75L4cvg6QKqxLUE7T9/d6GIk
djC7zkVSndb3yuKxGEa5F43Zpdv0C/PvN4aW4yKbBMLFs+EUNki4Rg3tEpDFTs40fbsG0Yq/qdDc
Gm0XR6Y9Un+YrUUqypsYrnWXsADb1guMGCVixvvRxsaBaZzCR+A3tGKyuRGTRiLq9glQBPVT8834
7SmWYxT76fqiF3m5Stu1AqVWVT0It2JC09vSX75gksnIT1EAlko0Mr+5mpmSq1g1XVY3Wd1Y4HYR
1l5n6XmzbrrhpWE0HvhHClu2bQnnSBBymyD9zAqN31GH+C+EUecl7dOGDm2UZkTdwyNcfPrbkl2n
YRR4mNdJqmP44xBFkJkW6rpL8PqqX5oN0APsn+0kf2JG/H22wjMbPqiEW3PmIX4pCw/qqk7W1dCp
2GTC670LQNHHB5gEsqCXAFihth3JsHEcfVkd+0DsDl+8BVrYAGJFIhgpfppCfh/wcb/mi1ThuzbV
0sAd2idruFFhOV4gUOJyrL04T9/gZxYsLSkfbaDO2go5Xf+N/Du/HrVmLkOQltySlk/Fqusvv5cR
KVxcGPh1MjsywxJ8e9UOWT9vK+/fkIqrq7lHS/YM4CKcn3cS41AcloUE0XUwrQDOgTPlUW+YXujw
n9Dr5M7L44axrk3356E8ajp+DhS3Ip5yk33ofitZe/0qQ8Ay+Ekd1hLXC50rGtnCY4ffcSdaHQ7S
c1vSCO61UdvjDMJgSXQaSZv15PQfKl0Oo/DkVEH75DTLDkKtAZqJVkLNeRWWCc/zGWk0tcWOm+Eg
HXBq35nmiNxnD95h9ZSpcme8gvmzJ56OI9sQYrGN8gfIeBZWz0mGVBIrrOBUdJlBMcZlwJhIBBRp
OVh6Dmg15wYq8qPV4uWcjmujopb9RMlsl1OMAQxJCuSBfN9XYJN6JmIzA8hdIClmxou7EkCyy9AY
8kryWtpqBnBjieNFQq7e61KEdT1fK4j+O/AepIqEA4Ff9UE1besoj6wK/0VH1Y1IjI3uU0U6hBHg
Z5t4WMEpdpU7iDfYZPF94146GFlZRQYdF5ySqEW3T7EHE36RltQaVyzPEfWbIaNJp+bqxxBRKxps
M+DJtNuQlrHBZy7t3/pQyZvjZrthgd3Q0NiK8dJa8ug4qsG/MBc0jOQVaCx942f+XlpjjL3BpRQT
SKMVIdtGHad+TXCCEvYI/nmRH1venSzxffrsHu4Y+yMQF609Csxz3MPPyh41NEgwM+XA259PxQrD
MQhVjdOvrxFHYTC/Pm6oiDq/SxCqqNqzaT7VQNbTgTZG/kXLiMfmTHS6Qk6h0aZn1CvIK0pBjEvW
STBqQf+3x5i5A0CoDmSnHE+gy5bMeFvsks3OLHeyAagzHPMrhi5tVNC7CYkohzjguqv9nO+OtMJu
N0lkcFSgF+6QcL4e5r8282Jt1DXPNe1Ua1qOngouPdyuaRMoCBa4sf0RS+VckfhlKfiRRyu0IYLl
HIspizzRZi0SAF7yJjeRhvN8kgz3m+hctpDSeIPXowfTjfp2Ph5uqTYg8/F5PK/uzV4blgl4nXFR
90nEoBnJjHSQ33hHkleL9UD4Qbq17deoVK36mApBXBFk/As++giM90m20GsnV/KCL9BvtdpESR77
S5bWUIs4ociej5DHFurud0NJp4UAZi5zRopHLxYjdWEhr8bfQbhXP3v6BWBWi8ADfNavTATzeQ20
sfoXO5RyXH32dpDD7PLJP7atSwJYM7eVFE4gO1kt9UHJYGoZiVPexh/BvSP7uPAjwXvL7HdA2rPp
XdZrPwd6HMn54RWJD/PKte/u0+P4UmM1wqWQJTdP6bmr7dJ50P4ujMwPkwDkE3BUnpX49zN1grX8
4VhsWZgfjd9xiErk0s8fZpgrzo36fLWkynBTWcGFCJ2OUV/efUrShfj8HDNa+luu7RAxGrSsOr8u
rLah1x8G4DHra1TSuQM1CR1NHFheBecXK78VbKBm0NlZ0psGDYlAWtMeUOJOcyJHNZn/JfPIDrjl
7Iep2JLomqTR8bN4RA3yni85l1YE+dBUpZmovjZ5rV2Aa4hC+rMrVMTbNQlhS5h2ygh9OEDdPpBE
brBW9AnfyZp7XSaAWIRcPA96AFGlisJDzlPdbUQKmxed9PTOneT+blhbtFIwurjV9MTwyMf+hnAD
e9Xpa3Br6vxe0XDs2/BrM876JnhO/VaOn4p4eBjRdWtmlT3tA1/qu5taqz4t8ODr24wST1pyWvCM
2p3lqBUHaTof9mzdP5+mK0vWAk51MnyKo9s1lGQ26RjFC9SxNGK/q304ua3NvielwgPwr86naMc0
zAgfFvHd4yikKBgLPVehXHjJmLYZ8wnUmiTEUZ96QaKI/spt4mGXZwjfXenPYDAanln2V8Bossda
nOnTUPeY/cwFJsk8CsWQzAs6/yYBb4VuiIm+2MGr5WB7D7CdKdKc14m1PL03lzq1leuc+mnUjQiz
r9fnglDXHbWZ971rdlcLwHVTrJAE/zNTyBuRd18dEKZDs8/fGlFIK8ByKcSHMVmvePNhtyePMVJX
+wK75as2Uw7/f4G1/HaKtFaT5dShMFzpqdXsv9lnrjs1lF/EBl5BDM5N1phDpBdfAPgiETg12aKh
B5PM5Tgqcc2Z+sfa9A/r5Ko2vQ15nHlxdTyvdWBnGK8YpazlHFyhH4dYm9inhuVg70rfauW8kbk/
6Bgc+f2ydv0WIXO+k6fbbR0LOuDXRahLTohQQQ5VQsaCsDhaoOHSWD6g5C6UrSooNkR/4WDuOGx4
RuLhGyC+j8k85tz8ge3l644HOlm5pBnVQZEs7vvmXl0HDfyB1X9ZYDA3+Uy5b+t2dmQ0Htl2tRij
3LLBXp3DDaeJLjPn3NBqek6/HKq0H2O1PKLDdTEQf7c146e1Hxu8XdpoKnsnB5qPddM0g7YRByzB
qIp/Lj2v3bIGSua2ltnc1PxIKk3XX92f+xtUdjlmA62dqWdPkmRan+CWwt1pkUdMzHmGzJELg+LJ
QTi7n9b79C/R0qEIK+qbSjy1ibBIUMlqspMnFPEn2LK1tA16Cy09fi81wyB1jat017cK1gBYHlG6
wSYA/xzflo8XxoeDfR1+MCxsMhwx6k4NQeT0Pi03mQXTtF0/RRlFXfgZZd5omMTajWM7Xe/tJzz5
eS3JbHU8N8AJzS3YxbUp8kUdfuWvM2Q0JgKp7rZg42tu+Rd86AKQueZe5GtAdv9HQuvmpiuQ4DhA
qtFpHf1x7yuGm55qwNqe02AxzfXtg+GWC5jsPPOVk7CJFQOJJ8yFY6ttVHUMSyUVoy1dtBocjrJa
UByiQnKgCzLxO+QT8wAinL06KzTjWmxj6pp5VJs9GNDg1MMCMFlYVmaaXSh3+DKFQZTJtW9tIcxQ
FaBmzGDqyFAH1CFZaEaQFROAwAs4eveCcyF5F4oYb5GpnB3FsEd8TWiLJmqHu4XSXEbuSjVMDia4
dHVXdOy55+EFNz8kKAhuSFG2wjCueAC2vAUkCJn3DaZ2IuT7rp9QL27D/J6RbMg3q1NqUUx+nutc
GpjRApwyp32w0882wDIWOd6js4H2vkbVp/Owl1XYHm0Ewitm6ydgMdyl/NhOGgslLm3xmfnhevUR
9qoFH30pRzmve6JcaafLEsquPkNKLucSFvez93xITWa/u5b5vDFNfBGVgIs55yzmCUCuOl7jZBdd
/VsRk4UjUAFrI0JiD4Ns7rhC/9DyTCzPmAHGUFHrL2hJ5Y57OrL9UGk8KeyXZMzb2bX04rCP11gQ
o/VaVimt/c2eH9v1XaRxZTsh8bao62z7ynTQ015bXcgspyIca5ivLY86S+VYvNMiRxJ0Ytr7Nken
P30uGpRIgizdTVxZnXnrBd61h2LR54TslBbsFo5BGgc4nRsqCbLn9LaTowUlEhnMzuNiXZApDJ5O
0OqGtxr6zDfx01ymh3OzoivDRtHzf59nFahBcTzKhSs+7B+34zaQFEA4gZSU/tt3Fk3tAjgaTVh3
m15FONI1Jd1rEviuS2iYtp0dcU5aQLtAivz5gJqS6qXk2M/IN2DlElxH+2Zzok+zY8VQ6UmIhFyL
rJClCrjw7aVCDgNUS9VC5XjRlqrpmRoa0P5MDaOwIK4/cI3xtDN3WKE3qCFAe+QRX2SelNqElkwk
rRfLZP0VMWbKdZegNW8rWBdoQdDs+q6SV6reaVffuD0W3OudAqn8ObZUXI0Ocd+0rj14YdekCjEr
mH+vrM4I2xPv4NlFQoRPwLdrSjj+47BZRdWxbmT5rQKbKYe8eVuKAO75PN68HGgCF4p4cIcJ5Lo9
E23srY/cxyU+TIJYnCE3s+KR1s3vS82I3afy74gcaL4V2WJOshEoe7Vj8RoRD1SfyF5Zcn5/4RKo
gjpfomDK7d0genKlZTiN/8kaRK885IPlg8KhLY7LIfszr4WWbiuwE5Xs/AFmONQBfOl5gI2emdKU
j1QiQzH2vhFGu3IisJ3o+NZzdaqfuZy7mnYl2SVpVNeCL7ee8fBPiFynm+Gp3Dzmb/SkHpN7Wwpq
0420JdzFBtezH6xUxa0V4bCvkKUnkRHCzWFw314TLyzcH57N3Uzb37H8Uslh/JrBIcoF4XGJGEi2
rppfEbUQCh7KhPxmnTOAIpQZMnif+su0+aZ1/z9qag+SqekcAdVvffqpW5I2qNLb2GDfqeSjlHCh
q1EmidGCuxvYJzvZuQPJoECTl5QkrrTkX3w9sEfOQCfYvu8jowmIA1AIXUur0wgdLt2QS//QpcL9
BiL9B5TAwCG82Acz0rVqjHf0QkCWTVkGtypYrvk1SPUvyNaenxsnKMexK8XBIgrVw3y8EWARB+ED
9dvK01+i5aERtZi76bskdOnVz82Smc6IRVvmQ1QRFDfmUE8hXrsHQiJtbS+Wg/4V1vdfk+QIWT+r
dOP/Verj4eaZUZ07WETADIXF0dqeiPUQ/OOj6ZxZeHZ/2Rwmn4spgfORm9fnJcvS1Ztfdk5Y6MJM
eHacc8htaohOndNHsSwxeZQ/cAasv6wX2XqD9JKu37CJnfOgfLCEMAmaAgdpstEF9EniRkcRWlnk
055xobkzFWaGMULWRfLx5Y4RmXHKjKvOwhmhEGc/T38jOA9A1AeVAlATw3C2iV3YHo8WNzAaKhkr
h50wfzDv5CYFFHDR0nISflCvt41PURDPUVtqKLrigdUm9yZOJj00JWo1YrEq3VzMKtsYK9W7vxM5
5Aur95pQ+FH7OHtBRIRvFwAhukj9XBjgQBaQzMAybjAjCc8XpUMy8GdoTiRuTwn55Ka6wK2bBuWg
YY1VD/QiNFD0Cov26AKSygKbBdIzwNBZjK/7gRuy3KkkLQdtrq9jigkcdLadobUyvMcsX+FrcKx+
56MHaAhvwuw7LpPFeYgEkW8Vxk2eyi9EHBg3pdzAnMqUgOzv+/EE5d/KDon/QvqEc+sLUMnor39z
aNJMxMur7cDSZ2hBNFr0oCPcJVjWGmkB6+g1dPDcpRaFf+e6XxMpzI3Ou+m10PbDIdXxDPlloK0Z
dHSrDTusmUV9R+llMF5W5xeHqAyk9Zouq2zhbtyAlVe2Mh0VGtAAoqHQBXKbMdlmAnnRtxhq4sro
b7TsBiLrYQ5QtH2rtghLe7xum01tp2krs8a77OVDmPbaqhWtcUnJkd0ZOUY2c+aXbT+FCx6SCGGa
pPreivOEEq+drMNgeWaoXtlO+TsSOrH2nJq2lZiuKjc3lF1etmR5tIfKLGiXUJhpsym2Z24t1OLa
uIB4zLP9VvqSl+jwig5Q66yE5Z5rHI0CQcZnhzy2rHRvhCWVcqffCoLl1dk4Qvb1XUKGBpQoYxTG
DxunsZYfwSc3sWuEzxlFTC9WIs91bHlATgsZt9m3ItSRyCCjGagaDogp6P/T4SMYH9uNylfecm2H
rfBgSLe4x1tugKbTSPVvgOmgGedz5Xr6X/32PAsBF0/jgEz87lBL4HcDSy+pcP3o4tE+yJsvPGFK
SKsicbiW26VY9ukEN3J93ZMm/aqeGQ9WaJPDenVDnxUyCgCCYap0K+G/j4tXkpr/6i88sVsbvCFd
xNnukO31Z57nRfEue1qfBRA9f6bMdiuN67QeGUEbuBpTmLfXnO0GS7T0qMwiJmfofWqR2iFkG6lv
EpcUn3vLwCihNG0igotH6ap+MSS4Tin+JAriSc9pJy8ZikCgu5353R3pDTe+GMwkJkc4g/JXVYxc
FR6t93Y729Bg+VOyowM98nYNakD9qusnfFrJMf5SQliuETpDWoZ6rHOoubC1dbKN/xoCiN8SF7j2
O5TJLk8Z0ioencQqDs6NBy1ob6He3z49gY43nUjkC7H+wjJs4snA3yDs0mWfGeJNiNJoqcMkeuRa
U/bt8Nso4mW6xgVW8sOPUMLSTEtf3FD6/GGVWY+hHo6kHVW2xzw2RjlwWLnKh2sHu9qXQnQoZmlo
1AYSuiYwn7KzytDy7ONChk14oeLIW7B+vVHZgixNbdhvGrl8iLCbRgl3Qeo1JXqvilg3KwZ1xk1E
xaXR/1BHPphUBg8SL49ttBSWsbkBwx9JbXt+2R45KS6jy4TuW9TCMXX3S7QazUtv0QyAh7qperMU
qbgetGUr7xuzSTtDu/TH3S/uoNONupS+OvDoiO5EO6MqwEcnGvaZiwpRGuzkKN+OKPCIiFIDNPcR
/iERiIQ3ujFyzm6ChZ58jMGdG0KdT29N7aoHE2Zzt5ctFmLxHXehHesGvwBEYmEu9PbHymvnFUJK
ZGJ1h/m8bmo7L95l/RX+Zyux1DUZym5mvEeVMAKLgQLHesRY9xJQElTr48XkbJSCuOJxM2xDRI2B
H9x0t5WU3zPW58UCEEXpXozWpeWnqeZx5nog8EBojQNhUlWqsD+TNk+80D3fjM1qbqnzwJSGUgC5
x7jZSKHHkJ142Uzh8KOaYh6zL+8nZBQb7YhgMLzSyyFcQmEPNacvjD3tlJ72OHyLR0qV/lMkSRR1
tB+g3zG0NjvNrOXzFkoaOWlBPvomjnrseZnssglQd6noLNw1txNUCfpVyOUkDK/KYrsOSIimqjXK
WrO+q4BDVhr0v6wTPD4gVFywEceH7c/1RYqX0HD3rgqGyVRN5sX8Yv3vBksf7rMZ6kncnEOCGL1h
iXqE8uwPVVSlli6f6yXk4Cb6tGVA8QA8FXtsUxp4KRmXgeCLYd/ywkB+MIWGb+ZyYifuha+36qyq
Lt3czgnaDE16FmphZsbFt4ij//GOf3s8ZhqHeJKtyHfsiibN8xa3lUZtfenix62W02xYp28nWzo8
anpFJt9Vb81i0kc9oTmiQrPgqIOwT2iNVU7hqgDQf65gbU3euFEfavhMExy/Kyd23lSw+nKeUdFL
L7ZuCc772pL7KPCSz0WEdSxXTnx3xyColqNQ0//jUGoeAbpKgQuFcGHnuUe50xuADoQjs4xetAro
/T5xat48Z+/rQ2y/vouOalOOhFAZtnl0XzqPgbodHwYAEbhAs846babc3cX++9rYHiSyo/eNGc8M
dIeeP8HzI4eli2JhxgOe4o6PJOTodX74nQnoIOpETT4GJvZhMu6fggS6eOJekCmLFXFKJVQP1zyb
QmNN2Va/TVye+6G0c4whWnT5QsAVdXQUFoM6SUfxwNjATPrg2nIizWpZCaMXJE+Q2NAwch9Gg+7m
fajSY4I9JrDLHeCGR9ArfsrkGaoyxoreju9NbNxwG9/ckTTO2AVbbRQLRPs3I7hu8WDP7fA3h7yO
+cnln3C/3O1xrETTAj7IVAOF/xYSIS2/H3Wsem3sQva3PvJqw03ByIInlem7tsb3Zh/irAn2lqYE
SsYOBR/UTvFTRw1E2pUChzViI4cDbdArccO8ExZj7sPj+uUnPGRTy+2DG00HmWDwFq9wmNY7FVPU
VZekMrw+lsPr44RIX2FFLtqb46dbv3dxtSnb5FZlT8EQGSJ8ST2GbZm41WqeSe4p0dmp2XVBjIRF
y/bLhkDsUxaVNNkJRGNplAdoS4gmOc8uOeYbPudFbMKcmXjiwfx4Ef2NhRCjWHKOu3LcBQwxkudy
0PCxE1jvYyoTxdFLkZf/SVyVLChZo4TyKPvpe9q2qi3CpUrOk93FNtP4QhPi73Emuq2D2toOTIqq
0mWUe8rHKrnieYMVkcYTumj7VtyxO4u3M90FwmNMGYG4bEFNvOWU0yjJ+boPubuF5E2ScbonHjoE
xtWFjvU+KlTdNLYPOaKiL6SCtxFILkHIrd8FanPLf8kNwGFqd81LXPTUirGfGJp+F3vFCz2COXb/
jLhw8nHeu+E5NJS/TOMFoUE6TVXiEKj6cmZcGGSrazihYjAdwmb51J9we+nBfvc1KG4aPOzf5DkK
GiNu2bjJEAYZd224tPxG17W+IetTYKM63PJhyxzwxTma8tpZJMyOtJOJDjmPPHDgy0LlsIQEoVYm
ISOIIFfuRaJ7u9hmpfHhC95u2CraEzX7MRZLkSUDKwvRm3/P6Nf5elgAr7+Yc9c6+5/M8bPgOZ8p
jOay20qzR3gcmHDv/3vM+8vyN2Mc179X7h8C8joJBpD/NUEby28JmaB01FhpwUV3TbBx2Dq+0clx
krd3f3K9LHuSsheLmGeos/n/XYr2xZt+AY/RnzqpRwUoerl/3g2gRXgfU5ZKcnYc0KMiDIjdU0lf
AynVrStjIokW2kxVZpcqOVOgoCGYWA2nUNIaOyo8SPCyZiaWSbF1H/GoIJK0DYF5HoBdLzYVu+TC
eVv1xInqW6fDBgup7wmz2TSDVUiCBbgYI185yVfb6G6TOSh9Y8q3GVKMx8/DI6ihRzaMk5pZG62j
I4DM380RpMvolRpOsFOpV8ra31n9vWpwuW+Wx3zMV13drlYhSsziCz4SNXilTfJFBHg25/MO7EGP
T0eTJZT+kxAD7dIkcQpskJCceclG2cWqn7ae9TSegENuwiTseIDJ5z1iXeQTdmnCLANzi0fopzXS
nUVRWCFsibnWw9CPXYkM+2/LkbdNSCJSw29QSPqld4g1rpensM085vDWwZSyntzCyVZvcF6uDvg8
T6vBunZfGmvGBiP3PazZaKpX9gS1sDG13E4+wHZ7l/it84ei+KPeypSDDNTyH6+C8KjpMBt85BfM
rP5jZyFuGnJVPHKVPc8GNpQNZ4ufoILDd/tzGSzhR+3WAe2BuYEVvD1S19ofPH75tz2qBWLX7Mi8
sJcia9Zr9zpu/ph6ZM+fx4LKvzYRjdYUez/YzcVpyYpCsgr5PkM08XXUJN8seEzd95L+YR7Pa+Zc
gJby2n01L7F4VMVayE3fdlB5+Y61GsSpa6D/hZZB045sXKKYCgstM4AdvvDmuSTkvgiSrMZfL7Nh
Gr9cMoyMBqLi6yPNoZ7CA8JRjsRt5jxmopi0m+9FmQMd57DsI572q54dWP6+POUFIXY3yqGK12/7
DWxCdnuqLan/TI/+udRauWC3iSYpFklkZHO3L+N/Yp9UWVih6FRZUH/KbKdcZW0k+GaXsOVxB6UJ
M1g+51EmpO3byrxD7JWEFYaP86SbWyzVc0ftIWyChT69DceTah6azIUPnSVAVod3MWxlU/yQFV7C
QhRX7RlYAOSKmKPqacbA3XqupIO8ZNOC51bxIVIl+8X2CwuJfFvQb6Y5G4yQX55xj/itNrK6DSu1
OyOQQ2MRsLeoUifEAjLdXu85hNQRH+I9X3+G5FZlEIVrpKJU7525zh9yIo3MPTZMiQesBxdyqM4I
yCHIkkoHjwjm/e4gCV2z+zSa5DfZsdLYMEaoJMcuEboXBqmAp/dDHWdismFZbVFrURD8T13aPc8K
Ktz65F72iIWBcnQ11cJBcapQqNSTkQ62pELiEeiQRBicNESEtQ1Bl9XCFIhha55W0hKsYJKmPhyz
YsrpOnYPL64ujUsF0wmv7v6a1b7Cz9jAMncQ+3iB5jMsthG3Kgs20FkJ3ybQIVjEChZ2T9oI8XOE
7qlH3v3rCAUpGFub0jDtOifj1RluJXDtzVXXfLqpkt2yn4MBltSxBWxCx1YFcsSTmE305zSmTOul
jsO+3oPnRtzAxVXyzd8wm5S9H4B/7bD2i9seexZWsHF6CVj5hwe6f1gf3ro6g/faQVyDO8i0SgHB
tyJbH7mx96vkHP9UU3Kp3o8v5JnuZpyAoOBoWgMOr8Nq/rlhG9a4/VhKhe2N0tdYQ+OgY8od1/iq
sgX00jd5ykkvTkFR0Uj1QfkrU/8nu+JdoPbTIL0pBwZoRKYUedibOgPA2sN9x+Yv6W8bgS8fgGy1
H3b9gzRmlgi6CZLOiLsYEu/Bw6+jMScGG4QbaZKG8jflg1k/Zjvc2vQacrszqTrLA0Kn/FUbcwkV
xgYXtI+PteDldYCpRjoDOWMwRLdOvDyxbJOIPcQjNHrb/2d8VZPgbSqynf2fbN+KbtpZ7sT1ZCST
ILnkYEAvPqJwCiBiDODlAMfFF2jeCF2XxnIvFkn/tgrlJzqCky/KfKkLv2aTPE1dBGZbJKvU9WbD
1JydqT7dfB3XqXdJOvrNkvQgLEQCyLee2gyOTV/bP5q0MvbgUTQVUszvBlk4hy5Z75uAAM4enHoT
gI/HpzGsqhxcHcggGMI/sNjWzU82xgm9vXYZI3XAp51sFzUdRqgLj+ccfJY07z/eZszRyPLGot1a
zzAfTOQ1JoUss2csxCjrY8M7ZZ55BtErz25BSC/eYc3no0rjUZF2Gh9nUHbXRiN7+yKeXTXR9jKd
lpqVMxDJuMroZbuCsZreED7GIuL6bMs2HCloUrud5HvOObFIf1CVTxWPZswxKpkn3/JIMe0Ptwgu
uJrT0j+ztZDEf/qZtiJNW5TQQ0QDiO2Hyr643Mw4vE340FWNHCIyx64o5ksrj3ENJspvQiWxPi3S
0JHkQBUYcViL+rXoPvRKLgQVxFKjhk8BQsyi35QcRVmUxWXsI/Adys+IxC9hJ2DMqQVHFLkwGWxi
WR0uues6HYlU+SFo2OaGmKT9syNatDJmGMpiGSs0mfRlavFO8OLH9jdjejrEY7HIWIdODk4hUT1P
po+xTAUThN933QIsgs52+u0tSHE31n2FvcAaYo3/+rnGGjC5t4f6mYIR98mBUA8zQhHXkZNNiSHz
lhXz4IL9zBYqt09VzeuBLktGpKJJ9qRUn4rZe7cQkaKZBkpl8eK3cTQW+2fuPC1iBRbbweqZwSPv
cnO/F8saodJd+S0OaRKq33k+og6gWnTEMdtZjhr5t3PFDm4lxC/Xp2lnZ30D8wRe1+mAwIW4KTqw
ey2lYlkt7F6Pof9kkmyQRUiZZVcy+4KBO9Q+xAQu81SkOfB7rU80CPtYg6q06KHp1C1gDBAmEYbW
WSfY8caIYcFL+3RIQR3X/J02OZJC2ERnOzUaGgrLEO6Ah4Bhdz6B/2ZKX0sKdQcRjPxTC1MlMWfB
t7VwbfeVZhcSHcD/csbPanuputYWD0h+rR3MPARQ3/2oFe3s19GOJl9FKYCpbutFDfTCGij0VpFy
IwWLuHbw7G94ENaoJp3tIHZznxPnDF2ZEr47hrsrjSUbJC2156DiSe+jJLUp0LqBDfMief1Vpwgh
F0Tdr9+tzV1yzPoKV6BYSJ5rj6E2/bVzmxUbePFAlDZ4VWM6BqIdBf2j3d4Zg1y7wQUYyczMICEd
FVcQnIBimShLPpzaqX9t0S7CjLjeYtqhlQi6k7lrnJLiZaKpholn4Z+0vtJpaO3VWGTGNvI+ESCl
rIwWzFEX/zMPAZW2YybnmGAH/z8K5lDIwjxhosv4Rk9tasldLcbAItIRb1ympC7KGSOEgsyM3NwN
tyddxjttnvYGUVfPbWzeRQpVwiMdY6lb2CXT4pVD88uywVoRbzC29NjQUk+jniCYfa8n9Nh9j9vg
q1ngxXefJ1BkUw8eG3HkCarpK8YSJml/Bc6SNRI0nu5JiEx8KB+nO/jBKSS9ay0BVoJVwABiUyWC
cUC2bfOn1xanCAULt8NNTJGc3VFQDnBw58QKm1M+CVz/6FMcAHFkliMNE/BRG6jzxN3LE110eLhr
yf4pCgIfAAmcIZD7sxWZAxo6DmkFSrc4QVYbUV5UtjKik5uT3A6oLHKm/q5d5O0qdDQ1XVmW3HxG
2BXmZCcuM9xxwBWo2nZSyqAJ+Lvg5/8Q7q3xwTgJvyLbIwpf0w7pXMWIXljLrRAua32ZqmWTC4K+
YMLWc1a4Qrvp+YF+BRjmkXUb/2NbWEYBO80gSQyrVx8L68W5rFY+pZ9gwVV948rsS43QVm7HZrxQ
ppWpFTMUfNu/D34Y+vhjDTCnoM47DRmaE2c3L8kqgdmhFESz9pmIVIMGnQedLNFNrricpp+Qai9K
YJmtZSQuToS6k+REfVIf34fzosbyAzSuBx6H/A+ydOXZKYM6H5BYnGcG8X8Dq+4fva6brh/luEfN
ipSdO6Cdeavudo+YjrSliq+Z+fEfyj/dS4XUjaQn2RtnLmQUJIrexBCW1ewRAjZi4HcqgXhgrKJv
S82La9Px/sGZOdEHDGxTHh2/EZbdh1N6L86yMX5J6XW7tDbvNNDBfsz+B8fUAvVaYJRgEIpHeNAc
LdyikNEMLAYBJdgvWRpVv3pimhNC21Ppo0x6UKX+qtRbSnWGuQhyPDR5zW3F6Gn3MtWdfmD+PmbH
6EXWtT845p7mnFUWd8hAppab9b0dv/pm3kBLkms/hg+h8AJGuv5vA7PvgtM5EjCL59EKkxLMOt1K
3Y34N+NPUL0iK/VZmaG6wq2eaWnuatTeUd2dXvBNmEqbGKq7+vcFNmwriaCW4wFtr6iLcSAYu33p
hsD1DuktDWDnRIBEnSSfZTjlK4dZFR6Iek6zF1WXjvbKKO/huQGz5qGIYAeZu5ZbSNNeVnoY+sZP
og1/M57RfTcRv+vkmCkagWcWWAJFTWvNn6kVZtnzEp/Tqh9oVnqpeOU7Px676rn10mgxKRfuYqCR
Tv4ZuXGtc8bamlJUslvHiPRUtB01ZZi85VtvYHN4oZ4EnoulRgOlYTfqyik/sM7HPxPnJpo2GtOb
3hmps+p6d1+fwQROdyOL3RIsY/QezBRWEk6CxFoPrNGcdqn4kuAy7iQhZdedzDjAGbx3TUDEiAcB
0ibGjYC+KQqOwyPCBn2ieLUAoslw+V0GDhvoLfIpV4RmmRWgyf0x1vq1lIKKHrXuIac1/gtKpkdr
D1Pn2Ip2RBqlfMQyyMA3gW8oCerXU6OI8K8Ph72lXk+SlACLNJPDGrkOSEzTOdXuQ2LHopsFquHj
K2WUI/WwlYPolPzh/hHdxbfBqdwWAocqkdJdsLc52IckxENfP+tgqzrZM+IoCqxau4MLZY18kx+8
tZx83/wsakL1yYir1kAWCmO9JeXqgfGar5do6g+qaC8yrfpsn8lsrEqvOuSRG7GRtTyfs+CmKcaE
QtPsJflwBAscNihVl1bcxW7IKfL3Y/MYxpKCc1zEAOFrRXks4lhK3X5naEzQatqxI6EbzthiaWB/
wvQ+PS1EeYd8viBQ8zGNuanaMMddLphu6Ip6SJgEb5PM/eLPFVX+8bx54GesBS/kM+nHwx3a+/ss
gTFpTRVYpZymcUY2ei4KHxz5OwmQieDCntb1prG8ciyC8Ta4fywNnMpfeNbu0JxUT0tSxIrtDLgf
h9SNQhUPTXjzASDOGhmRievSLG5mm+NtOK7SdGvj1b1QRPW+Ve2BwLUWLxs3L5aVO6Uaa0ruDoYE
V1dn8f49rl+c5faY6dkoimv2VzZggtITY3zxp7RfPmaAcZeQsD3NH0GNt5aHiscIwWI8S99SJkdd
yBAAJkdiuZvGO6+JW1eSo96a2BlPXYNeh5lZ0TkKp1Zmr2Od6gatd65fJsy/s1RUOKIvFPDGdFb7
y+Xc+x7G/MpMOqdUEjvHwlwFAxOIBNurk8+ZNRyfuV0JzhQFbsUwDo7yQN8z4Npri6aA5kLceD1S
OE+PTIPXV59smSN7/mzKbZLw0b/Nmu7WA/6vVhZiwf1gMnT1relqIIKpvRo8RyN1zbeVnvUPAUqP
k7D0W9nOn/gc6SfZTfcUzizuJLNoAyWWD5WCASZfUIKkYS7oCQCzTKwJ/Uhr7fmpGb9an+428KA5
X4X/+gIB3+H2N4j3uUVzi4A0FMJZQhD4Rmz05QX1TXtEclvKiFhg4GZ1+DoRtRUbiKgMLjQz5sgj
wdWR+so4tdbnJfRKhU/BDriGVOanhRtFFf/pBrjUJwTAhxRJxy4zX+tuHPqLGR5MA9EQkkelDTjj
puGcHINR5p7tkhDGT87ijvtq4dHYZ2a9MR5B+bylEgTMenBhm7whaaIR5mUYDlIDQ3KTTR/Kshe1
11YF0hyNAg32OJ5iYWe/OplhnpkwiO3d/Oma408C9IGG4ZtraIGXSc9ocq0A7OMm12fw+F7liqRd
gNPYxXzxxoAnRUtCM1plJjPd9Sy8m2n6z5tQyIp6MTCPDwPUU5BVzIyxj5p6qaeGQ9viM0exbUlD
UFlgCuSM9OQ5NgAkhoPosbfVZ9z9lus4U+vUmfbFhvPz4/PmDHAL7iBzY7dbd3adOEdnq/dRNt78
0vBo8dUHaRdp+NXKgN3rqyTPZKWefWvg3I3eab6NkAx7/m6ej2q2NzYhc5OGsB/NFfUWqXZBR4Rk
g3kv1Xmlrc50jjf12mRKVSguBKisqBdoZNMYUmtqBvueMWVXpkmriUtb0dTnvpcxWNU4Bgn/k/bD
7MsITrImCB0C2+SUHFu2WrqVNGXWLLL2IM/WeCgJLPC1HOY+3tIFnZUHjjGrtxwQvF1M3nEcSHf0
M7uVVLEDWg7XKmRU5MIZaF3LPIriIexOeihUJdwyioB9DuJTfQfckv6BY/67dBL5BLuceh90ps8w
HUZMvmACbCA/nq+SEcJUqpKCe3sVLVAt+bPGdcdhRUKBltS4Ra2WkaqY5v59Y/v2MH5mTVwgRtkv
k6IICrpsVtcQapJxDzy2/6BTLhqNJUxD4pTnDA/HmH+ko0Le8QOmdaHZkQSDx5xBkvdzUklkmC/H
SEI1IgnlkNutFWW3tMKYqrtm+iupVyJ7z06ln3jMCwfrVlkcgxQJjLvk/JOApE3VTKtlJT49dp+p
qqV2kBt7aKASBeZtIF7cCfQDbwYZ1cyoEiBDD7dWQ2n93EgbcPG2rp04clB02Pb+aRqSl4trAAMD
Cif4U2Dk/oe9dv5X+Ecw5NWrE6iO+GIegfbid8Cqt253+7w8vOFoFsc2/7CxspcHcNG6MN98ZeR9
+HBc7t8VeK3vRUFA++GyeChOrkg/2VIlO2tXb/53xbNsJaDo26NnvM6dxCsl+3Ql5A+B5XjEp9yF
3zQJAUMDCpV1ZMBK38mnEVuVRBKSm+6KAW/WpUf0wP86pSP4CaVs8kuFEoPiRC5+F2bPEM9yPpVB
mocxC/B3FSrzaLVWW0arOOoyQtTTttFp5Hi1TR36DTABTWvLGOdf7jIP4bwko6Kypy++ihFI3qUb
i3qQoLAjv0vWle0XgWxnwChZ+rMDBxuumgtr5ywzr41jC/uALkmoxnADu7tPqoV5iK/2oxpu89pC
YUseoOASorklECdi4u1uJ07mGexMVcrL0um/H3RESQAnNKCiRSnMBHXTiyC/M5OYDKhJzLe9CgnI
HaTP9VY0P+1xUrYgkQd3yCpMHtscQhxc/dv0mvnuI0D+kuPs8Kaotd/x385XERhtXR46HMy5yI6/
wwMKIZHq04UW8RjwSY9XmgmGd0M1tXVHjVAAGPX9A6FPdGeU++DpIvn0Qx5EvHvVYSau4y5nDCr0
dwwR6m230KEaMIr/xS3zyh+zkttvy3iB9eMjKeV4rm9lDQsmK+batV2VCzB6olj4htU3E1LMqvwU
yoaxapR7HxNt8g3W8FuvJSs11n5g4j9n/V7BxDhmjZMt6GIQc70jj2oRK99+Pun1EBBWY1fqjS41
yf8TIkmUFLMroJOb3MepZlDBuJ1c+qFsAVrXN79e7ypRZ4s2SUJ5b1fNJmBDsAZ0SoSOlcjbzhV9
U054V8m4/qE/haOzZnsFmMwxxTfn7mzi4KjWh7FT7o1FCXon9M1lpiVTehJXhF5Yvev1812x6kNc
RGQDce3JnLcnfkc0CnpZBqPRXJ+w6TMFhIGquB677nITa7xHG4bjQavbqSBH/qnS6+nMY2JrXK06
RwX7jICAlmSe/akmEEcX//FG7FcB9lBAEHWif2Ixwqaw7hXwOutGbhO9kyjDv1IfyE5jRcXa7IZ/
q8OLdGq55Flzc/TS+onv2K/olbeCwspbl2LLl/9h7xmqVVvgaoNbC3b/s1IFHl4PzYED+qkcNFns
4BN21QTLxMMsjpVWz3mKtiMVQ/W9B0mc9Bc9Ns1UTVgnF9wiNgDOXn8VbEmdMfCRedJQTgMLSNbi
QeG6SxbPRrQmki5zrguQ3Mc7j6FbLcRATStGue37bjF/qDn0wqAQnIQBg/42uydPkxIC2GCAybhH
AuvlEb8vu6btraPxVAZ4BSlnW7BJcpQvJHD6B25d+bFKKfB1ergn0HyoItC92+N5Z5wlFvjb0tjr
5YMaV65ynvn83RYBwlaDIo/yQrWtB7zNmh+U+tVyeq9dpYd0eh7cIWoZPkCb8R/N7UDWLPeiTyKX
rgk7PhjNSYg2hrdVkjAck8IdhYb0qsKSUEp5wkdc7gyPK5o8xyAX6A1ZAqsUa65p3xwCgIRVQNxH
l/JaZXAb/TBnk8Mfo+Oub9cwirjL1fycrPHsJVspAm8LHspJuXxsrDXhfQTcdyv3VwJmeM6qtnMK
NyvutLQRYr/cgpsyd0McKaIxlhz5CtSljVAOkGp/I0WZZK4gTd26mUFxaKBK8/76N8aDzHyJ77E0
ekAcri8dxVnuXekx86XyqKIF2mXFjHGXEnWIYSiu5V7GZfFqlouvurblmo2hHxyUYD85O3S3XZgH
iIh6B/x+eGFWK4PEeiBlmDTfMsT1eogbfMaj2fm1nmWQpQQZrJkpTVLQ597IRb+NpYUXtA1muwde
bwBVyg4KKtdOagAQaheKHDrq4UMa85fEutR4deNhrLyeUcrlbnh1dRS0y9oHsyeBDLu4E3Dp8r0Q
kdKa9Cm830r3kOM8VlEQwdOrogvtMNkf9UA0QoJtUya7oZih90EjjMhQukTYG3o8YGpwflr89wNe
czffYOX72qHoJs4Kv2+5GF/QQkNFQosOA29SDicqvkxI0PAPmUIjK77dO4I7PdZcds1feY88sxV+
d0Gt24jtRNegqr0F+EJE7+B35EvwsW0NxSB1uoYiPENz8glKuyAfqPP7WNQ5Aa2c8PSoLEF16SqS
GTRcqyUohQUjeWO7DvM1Lsd8jS0/VOoKoGYbSufagtBnyNHOai+CK9BGhVb8aNL/TMni4ejbZBNY
FmRYttrvYpTdwQC43ZRG9Evg75s/dqz+1aVrJvR7QPYc59WnMHtEfzOnMN3fxYi235DSjz5KHUIz
y4WwYqaV0eQtVGgULMtcc24lyDkFdKkan+SIMHgnV63+E36QaVc3JUlQh8NGLqnHuSNKXkiPgY/T
VTJOXpxkflEF0RlcdPIfeYZQZqqEvo1+qGBGxlraq+3Lxu7gEVak+RrRP5MLaDk2fdO4m3VFYGYP
i9wpfRasvBNxlgHuifX6ciB4AT/WumxNxve6HBbwdJcSZxiKQjEsuqAn3LsbwiIIP236vPmE5Zm4
QHNWSNqStTm8RA5m1vGiLzLXcHG0MFjWxooVhKOMlDlgkwTwDPBD1qvU44I2/sIQDBeZs5ueTer7
9m8ziAJ7dXZzpfC8v25d7Dn6cqgmcprDItQqGjq6KA55HRy2DgR6PBW7b/ucgHDX/bBOFapT+t3Z
M/xaA4ImaV89rgQ2+VeC8vtKYlynMazi8utQMhmTmGvCXJjW5PVvMBP9WNVMXD2XWm9iksihE2Fd
Z153xtHmNHeTCL2tP0BX6QbrBt2FfMAMhwlgJhbvPQRCCM5hfaiUH5+kTqK3e/0joU9g1qExNylD
WQ8Vu046v0G47IMNijHwMP16lTicvihiv8sxNpKjUiufRKpso1faRZy1O1b/M457dXulvI9VnHx0
tT4YSCHK/bq+j8MIcJ55HkFRnncbhaCi/JEP3IQLkN6cW2YLc1Q8dgregwEOLoMDZyswVDCKxQJC
w0EDQdO3ACkOx/I3wMw2mqt1g9WeoYQfX4i2gQQgp32UslFkejN7Ml61NhhXmS+BE9A0eaaMkAh3
s1/MxJm1sXPmiXHaa45Mw9n8U5Gfx9vNn3pgvE2YAYXEk6DbbpnIwCy96wFvhzBACHiFEJtC67qH
LXmC9xsdjqFjgVlAi5IVIsCJX4WDpxT/0NkH34A/tOrZuWjYKwqa46r1JGhSw7hgMmvXNOSGW6sR
fvx8JwICbtq0wPXvNnHmuN02uLe2/xzF3mQhEtCdkeKKcZMVxNH2yWrbVqBMjHRepC2d8ztl9Mi2
JUwL5I6RKMElqaDrMxZEAM3eKFTzm4VGae8GApaSgt5xxHZn4s8o/US4mfulHBG8pfAFRu1Dlk7R
167q0vQg9dLQwGO6Jt5xZCX1k5/iy3gAAFZTNm1m59k6Gy5GMetM43mGoZuKE212wwV0M1aPiZ7W
kdX5HkpbJPSk9MZAXXS+iv5CSZZ1ItBuf/8ywVuRV8iHq6f0YkrBHmN2UGq9gkTEFnbDef7k0eWJ
YydsrjBo74nZdS2T2lNCGqlICLk64ZYSeAISv4KiSZhA9cmf/VIaDm+BfQWDE49FzYliZYvGesGc
i6/OB/pmhTwXqRXKyUncDNGeUyG/BAI6Vs9mTEjBji21ZNTry197ykJ0HiPWRW490SKRnQOt9+/j
LLt3I4ncmNsPBM2Qd2siD/hJQFeq2fbl7/px5Z/MnVQ+P+dc7byvyn068MdgSA+B6Ve5rDpZROZz
mlTr6GF53r1Jnr5WNEnTO01n7U0KkT1S9oHpkFvJdMS4qs35ilLj619pjwMIEvLBZfia/AcRgz6N
tDjW1aXFeSI5i0UzY3WrO//GV/sX4Ytk7ITyy4OXg1PrCqDa4HhaECPjXx4Ll8a5hSb8lm6KEgvn
WY9e1J3l0CH1grN6gpH6zX00SVN0tv8tovbhAw+B1ncWVDOBqIVsKgWR8nN2U94JuE7RqTF4FYoZ
xXik6MEHm+603GPQadQYS0fHMo7h2cC5GG4QuCiER/OmXsoWRZNR5Fk2cmFhd7dWNX3EHdZY6NSQ
KqZ2unigYaxXZdVHnq5V4yUc677EogkiGXxTgZYWD7O+DMrqQH+bF0ho9HgzdnJyApIqx/w74kGL
ByWhV+oTLxAc2kZuLGKi3ENMu4+KZF5h5qDkTy2HZvEZfmxtYjAbi+0lYz+r+vy+48yGOvyLpZF7
FrgcVIE9QUSoxs1eMZ6muOdVNb5XtTQio/NR/0n9hX/0sGPFv8rknfNYZCZcPBFwHAMADCtqMvEP
9xzrXatqZ4wmyY2HPcIYX6Q1sx0CKO2KqjzcZpo+R+pfT0xKMa59rvZe+cZjFx6fbhk9/pbNrLSR
3ymUASckG5vWuNzUPKdamyRZK6oinlhAY9svauv5TxkNxvKY80rvzcoY5H1SxeJjtRG++hFc2VY4
ybT0H8CTipj987JZHmFVf4iWxzIJmt5Hm/D2wXUygfYP1PSs7e9k9Q1tkcF6ct4f8fVFbq7NwNjS
2dHiVX2uXM/ashLX1PswXFX831fyvSkeoxMnV9pCiE3veySfPlfD7nu4Ux1j9FyicuaHtf6j4aIi
2pfbAOx3DVJEwAnJrgN8U2wqf/k/zsAl0vqZFot78WbBoD61ICNfZzA7kCCQQ2G8iXjk8ui6ga60
22zUVLCeHDkmzxlG5n9Ks+ZjnCMoAwv4Mmb8DuQ0bjb3Pi2pLvfYTloh0ihcpAWHvobv0I3e5wkz
iQXhs7SyaLTiKwqCNqnYYcB7JFL7NHhbiEQF2c+5/X/bqFZfsJ6vdslBrErdUz9oMPXP5NcJQTPF
rsjsVJw2I1I+MG2OvMn9QUmnDxXvgYXysFU1yMNm6qRjbhWliDgrrzGhR1kqsavWLXZreWMsc2IK
EksRkfv3BmPV326R/GNmzB+6ItY/8bT9WxaM+qnxPH+xjPpoaUvrgNAljGsQZgMEWgtrmMZ8FT79
NvhqO7zZjchjJMu5BIjYEL1t4osPDdfD/8aNg2FocL2WXX72UcCIN5WJlpzXXbBnfJldLNtNX/Kf
iCBBBZcvfgBFuG1BRNH6mic+jn0eFM2i+ic6LEXgPivi4DFpqYQoP7sZqBuiRyLyG/KGel+r30kd
OGxWe7iq4fyJ9OE7ym60JhqUJG3IRRdn9pYyxaY+/FUnUukOG24DfbaBKZQcAiWvS0aQDRf4MhGb
ghJ0kfT0gHD+RgXIaZ9R/I+qgG0U5eP0AGPcAi+NRbidnupFsdKg4XRPS3LF5Z5dPZ2MhnRa09g8
Xxhfwm+qQ+b8jCcunWCOw1OaqjjFdpnpPHN7eFPuGzJSCPAAgCZ+FPgtgYkCT/zZzkrCg54iDyR6
ph63084lXWv46z8jpF0LOnn+ty2tzStBK+HXuoVs8XpCkyAdN9gStXqSw49hRQdZ70OfynryJcoP
6hyyMduBLHXA/dePPHLmGq7utxgX1Wp+YO3O31P4IjxqzoIXzVN+XRKF2C2taGU7rcXbLZyc7fZo
gdWAp+2Pju3seJGV+Mv10aWo/QzN1li+IkWkKpNFFcIP4U/mh8RXiRfyK9tv57/KICUfFWRikLty
wqi66gnkjNOr3msMtoVNUXUf5UDQp+2MjsMOgsDmxeUvcSLbmINbjqHmrUNYQ7bdPEO5cWZ71/+O
2pEIw2OcVk+Vy5eAB++Aradq2Q3GBdHIoNCVXkAaypd9X7HejiA5qJ75UnnL4UNxLCEN313wq7Lc
1xOWHzBeGLkeINOyBgImOKbNdjNTAhhYnDQjE55IihCvvcBSa7/niaIhfiUx/mDkUMLPUiXWc4kr
1PQ/YUYwGVa6cKC2Wiv+81S+e1cM8MpOh0a1yfC5+cnlmU4cfTpfyshp1HFbzbBySnqOcK7o+6Mr
UWkYSL+838Ez1ROCH9LXmJ/DWwv5ZneYAQYPd6z6haBUywH7KDC1JhDg+yESSfXghh85kQf/sTqC
ZAFwVaiHZU8qH9Km4UxdGMBXnF8YIeIXc2jKwCeMdsG77X4xu9BRni8LPJhzujozDsijTR1dGXnT
6DC6lmKiPurrqgJKJfY8TN3+AziXJyAvquchowRMF4hT4UbpQu/XbKcENFFbyZll46nBJGiZS5Mg
C5FVXZvxjI4kozxxW2akVlDirfk0KgOfEmRAE5MMH9yRGxgEmDVra8PFQ8O6wsDJz0zp1oaYU6I3
1NPWoRreWSaqiCB1wmj8XVnIvlNx1nzG5u8zZavP4nWfUssizW6HWVyOWfdvCSGhQQyCO0MVlCkz
TCY+Ehz9Fel7QdBd+J9EVO41zUuzufBIO0O+tL92yfbM1+7DhgAPnb2tEdv7VlbThzYG7xTDCbQS
euGOHRTP63vcIwJ4et/MuC0BMkGv/6HczWJfJfRI405VkLsCH0qPZNM4ozdPiLJOcmAw/n34Y/oc
2NQ6MZy9F2PRAEn1dJa4nngP63UN3Q/IQELPDO2NgMPvvpRKy2yVx35nIilHc8MCk4s+r/H7mKxn
GN9A2yPZu4c246eKyQyceoEsVUS+HN7gmYInzWpecAB5Ds3HAWXGpvTHbaJ0povz4D7yA3HuE4oI
JstlBICO8H+CKGLanPkPLfcMKZi6mf7HQTDmAVPdOvvDuAZoIBVjNrFYvrMokURi/ZRdLlOgnOH1
sSL6tidbYxIwmSNasYHyt7qqeyvoaqSzkxGBxG++KnBJsom6d+rfZgRT+2RkJTddMv6Gh38ELiiL
7ezp2nK2dpbKWXzTMc+j5qEoSK0tbe/tMxdrKgbkIa57GACye3a3JzDFSRrXYVGqt/8M53AT8Hoy
EJ9mjGhb4i12kZsobal/bjD19bmUUWSaZCae6VYYA2YWEVRbNFCHTeAL0Zsj1l+X2od0KWrWit1V
KwxlUmOtLzt/cI943NelkdvVpX2UqKF6Wq3Olj0oeauhw63CcNG0Rbp7P+Svnq1Gda2Z4Oo9t4oz
hTbSQuNvLZUG+V72JqoIc31hxgAzh0DEZQ6/Km3GQfYQ3YGkFdzAnhNW/RkWSZPK4SkxmOD3gmOY
L+7JRMBJiZZ3zGcxZsG3BfIxWDqLeNujaCAyeqK+hRXlYBN8wHg/FfOMBXWxN1sPe6btif6ztysu
Fq4PruN+tY/OOXVUEq7+z07gna1UE59F2APe3e3unT4plelDSnMbjcWozyk5OhScEDPJnKqxrBWl
Ys/kYcTyoF7Omq6WmL72fWGQreO8o/U+R0mw5lS/8ft4Qi1EWOtOZpSPl6fqrGM3YQPfNPcxWUaq
ATUg+YgkG1SgRqxxa+zEq0vkVaPfy/7ASoas02W/sab94qVqHz8mQLavX9RTi+SpXKEiuIgwI4AN
PxtG5m6V7kXkMTtqqx1LXVuWoHihd6aR76wIZSPjTSCyRZzPMiXh9rpe1voc7vwmoSbFZjTQRm6D
NDCBEIOsFXnd713gkECjr6N2+PX4vkLEAZSXeO8Yk3vKFgjeIRDw19mRRa4nVh+UCQfaS9KCFeY3
CmDYmtz3bxAsXxcvvpNF+5HMlhHqKDRIHQAjoX4lDVaPZMIWqOtsK2Fz8lLc9NGZ4m70F3GcCQNF
nx0OGjJIYJsxPlDeXJzKNhNy9a3tzKUbGUBKTUqKTYwvRLo6CnFKsTma1nNiJbMYp9u9tpg4uoMv
Gz7EgLft5i802ZWwB0aZcX5N5FrfsdvJ7/+F1zhgN00s0kVfROhlL9UvXclOvCpUafl247DjgX1T
QJJ77JWm6DwYZ/eKTHaDaebifWWUG2AgkxGGHzZY+uM7/T3Dd+4dKPtS5tQLMJled66JhkzZpuXu
p5fIXBVaEVWmcfAZd+c/2TCI1xFzaEmOX7YunxmYABChV3QBvqr94dKIzMVu1Ry/tCDb6a/WQX1C
kwHpqcH/FOQoe4jUxYCvnUo8KP/Ya0AdqqNwL2ENSBpkg8gpKiDl30zB6ltsNyvcEqEMXBgCcgGb
G6vQ30tP1x7iCphR5WXwjdpe60GjFtFcRYB2gexcajfE0stWMYwEO6/8v6rndqucPoPAk0t9meBL
4zexHu9C3RFVgt7rnpVTZDEJ/OI909+b9w7d3uYSlSOaKXo9KNthTNzKkriAaKGP2eAc1GvJJFbu
c8rm8tCaOmbe8LuxyQNlBvdHyVZ4ChOY5DXGE4wvQvBtyRGSECDmqW9utUAmjz+iEZg8ABI9oHzA
f3DTBTAbfInHol188DYFIs7PXY6falaUUZiZY4WsudIc/Xk10KmjqAZVVlL0ZTM+e1AUH2tzMQk/
9ABkVTst3KCRvHHfA16TToLSjY2xdGi9DRr8BdBQIMA8p4Xq3qA9/ByDAn24PnummP6gS54GFAEJ
Sr+yYu9IWqyJRGFMVOIEkoYDekhWutw2mvSdtlltwqEHgSEByV1r9DkijuFQwn/puMCl+Fr4f0zo
qovlTutRL7OELBJiSb/t4n4gcMSEblghemQt4U1PT2Vca4jBIwUuRHauHw+qcngHXtsVyE0+4ask
smw1qqMCUs4jIEwoefU11ftrX/yzdRqktElAuE5BQpVrRjwaR24phkv8KZBJmBDjSkhtfupZcilV
wMiBKazU/0NcLPOttI8s5RVFWm0SVSJCqTfz4n6NSD8L/lib9e5eU+H9qa+t2u3yRlsRn9EEdAnK
YLTNCiJa8S13uhl1GrSP/AoOtfOPbgXxhiD+30HMihm1fiu04inrC1kIMP0sFrM2rV7a6+uLpgWA
ZNlI8Mauj2bYwDVO6iUSmbWvFlYpO8FzNBLcWq1oi0Ecwk5fcPivkjmCwTH89E3+sKZQHVMowPPc
i8Zq378hmbD8E1WGDo6K4Vmb7WA2RQtFm5+I1UHNIRz7csobJthFO8wGd7dXYQwxfhIQwowNmznd
1yMg0OsstNjGBdJh2wm6sQHz3ZQ6tBMYFx6sWjJuCg8FwZqc7/9nM/9ljchb+K0CmVpu4eCM1vhJ
GJjsdwkewuvbg9MSwRe0oDQdT6YaXOXBB8GIzPDk8Jzc1PXb+xp3bprFrU1AZg5xu+qn75H5YAcZ
w+G3DTxm8n2fS9Putcv3rPP1d+Sye/eVpXzYvZ2xUSph+bVn8Ez5B8YAUVfXS1mz/qoviVbN0fUf
rwaT3YCgWVPOtKCP6zY2tBXGx8AaefVju7XxW7UhAT3sf+En0kn4Z/zC8rW87IDizQxtlJW7tAMN
C+QoMVSKQSLjmY90nIWkrl+H+TVarR1MVlf5hgonl0gUWQ0smBV0HjChPucW+OT4u53BNjJXw54/
AD/l+l/m1nAHGGKtFnGyjHSW+AWi5uZ66NcEmXNb1orc9++lTA2v3fVAh+W0FLSaQmpnFeUlUYdM
+YVEwY4aRwn4hT0dpMFbWVkP7RZvyS7VCKUQSLTertjK/TWtmSlhlasms68NvnC20H0FqwM3xz00
mO/COCLFosPE7qWAMiA29GyoIH6G2nFwRTitgKh52gFtD/ZUXc1s0yZ06TdYC2mVYN/eo+1gAbKS
eygLICtkAvBOwuXMWE6kBwqc6aK4yu1CZ2n41GH9ejg3TVuSxfX0BGO54CnrS/mKcN8gY/U5LKmr
c/vbuMfNwhiqajdxNrXdXhcDc924mEZGnLoyGXkXC6Ayk14VdGbgjGcnZxc3Uci0U5we3h7FTLA7
CvY1OA8CYCmhb1ZuU5P4Mr/W+am7kcHJj8KkGlCCVvTpCP3eDXa5c/wb0NFJa+9xIZQENZJ1NtVG
iVIn7w50YmsDW8VvyX1ylSdsKBYHbUzXE7jwNe9YeBmq7hJGOy8cKH7k/5uEmCV1QW2vt9rhl65X
auDZXCSUqTLQiaZku9iS8jLTUrC9k+uFgrK0cCvMC4II96PPm1xJMkGzTivIop1SCoIUqd6aglzo
XlKOxN+jSY2sOesAFTAdTGaPA+pFw5oOG3mYuPec0bN7ecPM8lkc6n+EPs/6FrF1gyfjHZRO/0La
4T3UkAUgunmxRUOrCVQ5tr6ljQu8fRMKEz2Sa03lTqRLgmNc6LiFu2GQ3dI6HDDIBIEOWvVtDmja
dQl1tsoH6GZ8ID0sDjhTdbJFFsX+TNJasCBN3TCSAoBFErx8YlgsHcjD03VsPMXLmcWr7RbzdwnW
yxKCgr4V3V/5ZgNtHkKInlXMFz98briCy9V4grO0wJHODfC6Yt4rLa9zZkaIfZhu9xN2C3DVpTdU
9I0a1ynmykt1iGZT18yVq8cGgRBocvBMAOpEt61WuthbUvwqbgBn4J8h+Ei6fNQQEcr3Cc8fUG2+
+vdOCAPFrNGGUeGzhCgJ7M2kI39FrWcSCF5o2VPu/TLd6rXz1CQRxudlk51ybq6fvHb2t4aqYhFZ
6tNLFnK+9wazCNVdb2PigfhT4soUMGP0/FAWKcW4iL/sjiDO+nMV3HMroHN2ElB3L9o0P72v3CQq
oK6+ZVrZT1yrkcTm5qmzJCV3+RQzBAeCfHWzM030kNkU/+XWb9cH29lH9x1EZYiD6FRrT2IG+9IG
iTtddmlzHC+NRU+auv722KJqs+a0XgeF/fUB8FJP1cAKiInWw2HcV4+nzH4soUtBr0+ASzKGl+Kt
MKSJkXod/bsqVUgQNbz4GRInF8h7O+mu68S/pNnQMLeKa+7WncPea1HdVAvhuMwIy+NEwj9AgZns
6Nw0tDhZJHXt0RQI2fuQfwFlg5kL+9kuF6ey10fZ9pID3IU5IpGWU/rOzLJKvjE3ApFC6JZUQU/k
CybYWGikPDiQnwqvNqwB9OcApaTUQ6aq9ODvrO+M6n7FFHKVqh+VbkS66L1NEbg2wrjUESaA1lbG
+DkuepNZmgyMCwguJt5dd0d7poL7d7mww0dbYV1kRM0DjwYuOD9SOyrtwfP8mopAnIqFTHfjHMSX
9LFzAmR18t9Sg2egEBGWBWApl+pQ6FbgsaYbtxsZ4F60MZYn/kp5eoE2fBn93x7CvnYi/1bizf/h
JcX9q/8He5FSrqwLMuk49MPvWoVoFzX/OHDjshexgbqlSTUXjWKxsvugonElAl0fzPS0RLZcK81q
MxFU97SCtq1APc3/6IL2WQZRvdGIZvOoY/XXb2xNZgwyD703eoI+6y29NJ5Dch9zrKbXCFsrZaFO
T9IoXeMuEk4jxvG/IElt3FixbniZOiGYOUFH/dz9OoWaMhngvt+tfKDnDXugGSW0hUNTLFsCne5Y
7jxpU/dsXAlt6XJtfKz+x1eSSVkw9vNh0E9rHA61k8w8p1+tZnGBEjoap7TKihLme8RzrujpYBCh
vpd5TRvMWKwlWySJq9pPuhX1XEnwdgCYHm3vYrXT5PRLoYBit+4VQqQP6oCKOSlYfkQuleZ+2kaO
JQcdALljUiMFwsu3p9bvyL1x/feb/HZG4eHxNqGO7RZ87/Wk2mupwPlx0HYsWeg6bXrPfr/I+Ev+
Z7Yecjye3pcuoQaiu3DXy07mN073P0wTyR+YXVQuL//vHXBBLJ7M/ShvEPe9+UPPoP8mVAqcQR5C
eIHm/FPbZUYjvBinIUXTr//wIEmO946l5TPZ3l8UbPZgkEypymN7w4lYGXFvMjaFx5Fn2gWmhhzd
/O9CxBpqLx0ZbJREnGOmIjxD+NVFJ/4qB39/637RbKdae5cPFiKEuSJm447dn4As8QRAvRBSNHEp
UGEqCgc9szinYHkmu17Y4u2Kqn+qbnNouNSdXlrJyS+/oRgEmusuQTQD7Urkb2F/Xuk0qtYrEuPs
cpw+bSkG0XxsCZdDYX4DpE2pPEM8n4XanqaGiw/2aLuJERLZzXncgOY2yOA6pIEgZJEj2k7vRuBx
F5b6QU196G7FShezVM8j9pMwBcc4HZRFmXMyNU2L/GG7hURNSGhcPG1xQbdTN3osZKKyIF9r08T/
GIxS+t2OcTuv7BSWCP/WA94yg1DDvPbt9oPpf0PM0MlWWd36wHG565fDv1MbQESN5YSFkQP3drh7
N65Tw19oS/2TB2NYmBC2n4XEvJFQHIjb6N91WUnQ43HaK04REkduhWeg8JDRRgzAJZj7qAJ42AZ9
RkXrT22umhToY3jDEYbCTOdI7bF9wvw9QQ91XiBrTgl3hO78+B+87sF8JN0f32ML9+rqXZvOUMKh
HSnU9fUxJJqRHbNtW0VQmfjbjS9HO2rFcjhbfCJ4toTqPkgfV8HX5MAouyaOrD86zihgN0Kybklq
b9mJeJD8poBQLUgECxTFt2dOHYDt5VHPQq8QyisFh/LROra9GXEXBl/mlZeE3ojODez+fV2maVLd
Dw8tKOwgHYo0THN8Tp9+JD90WBZYmfDt4/PyNTT6QTX8s35Aux/qG+oNY0Om2aO9qKUoL4HjmgYg
qZNrsFQbHaXOVnT4eyQtkNSUZpcoJRYxWF0W88wSLZQbJjq12DVffV4kK/RfJBCpsrAJS0PHTF/V
LIVBFlGh0IvCMZQhHbfLZEsTdRMnRreRgfDOFecvvHFnyO/bakFPZRZQ7Ai/qrAHwposHrr310Kn
unqoInYFIxdrc0eHyw7rZdXuVS5mk6mvmPC/W36WNrK0Kt1m0131jrMcodqBmPRhgTp+SGmSo44H
rv85KnMuTXmAHaUvnhH53DQZqEv62/v1laCFu498sbz0vNrMeDJG7YZ75cphjqOlC2LicOLHQK2o
L4tc+F94mipgNcpiG8rG1+iyFih47vmKAqTz/Nx+c9kBn8LSI064h3MO4lep6ojdRVIkcdWReoUT
lfK44gWXt+MrVAay3C/LHSooMI2vsw+f/G2+rotsPOIGJBbA92v/4keE1pd60pzr0V3lCM9X7HUn
vMhE5I0ZblgpXTQ3gPpcTrJVKBLr1j4CrSleIhVGTHL88FltOAsxgR+MrfTlTI2bHkf4QrD999Sq
F0VI+tdjipUMCm8+w0DokBCpJ2UmcJFy8kP1UHswDjeOJAX4IgyM74MPmSu57sXbIFZaQJb1kCzT
oEM+NyW5V2oRpnoiDKCXcResvRWV0Rhz6C60ngo6dNMHrO4pNVNwDaSK6FbzgA3jo7Mndv227nOs
sVOFv2ZxeLHGH0xbXTKmtuw8DHwZTVh4QZuD5dvb68MQPBdd2ijVOlKBfO7Mda+EEeT+HDVtSVaw
xhPQyzPov5lvLuu5w+POQzEiFGyIpGNC6kkzkJ8Mya3WwHRNPOXFv9OeIm+3nk9W9M3+o1MY6aps
UiuDaBX/7lYgMFfBUe3vFrUkZ8rs5kxLy0kIUz4VAuZDTFuS4Gk47X+63F8qkuGSpd1JqC6PN5ac
Tmasm9mSztqXV/tVtyaUB+n3+spOTQjvDX2kYH34YOaHZGUhTjdplDJuU7rR+EwLswonQW/totTJ
x9/FKLpDHW5ZyVAoWK0oewI1x+TVhy6tIXJgOY+bbnb6g69u2PZ8KMwb84kMftDu6odAMc/VIL2f
gP83EtfvKS/9wmjpDsrAfV6YRqRpAdOnaitk8QuHQcyoXmSfcZGt6T0YrOxHSwu8DtU0OeMBgPL5
FePQpqjeib//oo7Vnqqq6WnyJtm+7JpGpjhj8C22WHAVZWgd5kp0VEGlq1Hc18IgxjS+7uRKVMep
HMSqJVJeNRdwY+nOwIdokNpnZ1neViuG9tYooUnrUjMpelf0MVXIuw1NreFqzY1LpijKac27laT+
OHXa/L5WuaWfOArT8kvRU9QtmCxHFencutyA2arrlP08aTDmbkZyeIMUtTaYPEuPcgOju71u7zqH
lZIowwbGPwXRDNzqLzPb7b/QLatBeaSIbz5ISVB7hSThCwu0bkfVr216W4LuJa6esfwfrBfYMiJx
E0L5b6qLUY7Qn/veYYnR7izXgwf6UdI6Uz57AM+Z/cVQUel8TiAQscjxp6oN2nzAh8SoXDOWXKlc
fSA9zX9YAn0YWbOn6e8gP1RQDYIa6l7EUIHlI9JA+MNyUtDKeXpMVB095HUnyvLCua56lbhEMV/1
4z89OYN9yKRq6NRZ4ae9WrfE8XHi36M382HMUXoYhAYbG1jeIHrgSrcYM6T9EQYiLfVl/gWXAYgh
4/gtQM8Fqd/BOQW252TtTxYRmX+ctzeFrv1swFyV94pmCBAEACcBy+IF5KmrlzE+IN0h4gaPbdSs
WaDv01+7rOEDeQ+jDw9FjVN2BXANztZjgJLktTqoRPOlYvPkw59PEMB/rFkku8nCikx9l62LZhTD
cmEUoa4GayENIsFAJ1iAa/3GGEz2OzcyyVIBfnfj3debgMF2lcA4wzSb6BqlvTLFWOavEzdKIH9R
eDCG/EfzUSKbMSYseQ3Aj6w2AyEdfC7kvJq/Jfs9KJCVzQBU3HYO2VDcx4N8sT9r89orH8LWrADa
t2jS8JRuAKYfgMSAiihnUEw5sNkP8Syd4msoR4PZany8IDISUkGGfbEw9QXhpbJu5H+GaGt+bRVi
41J/11DPtYPS8rpkdMrPEC5G7PMLhXsP18674z6QyQac2Jd1rSWOWqlPDAlMqGbC7NkC5pGghRyl
VQ1zBBtXbrGaB+l2A5Uhjc8feC0m4T+a16jsMVLmv0e2bH13zQgOai9Khx7kgZvFWYer4mKBs4de
8V5ECJr1qf/fUUmAX5hj2PwKNgNWT1bFzSetgYYvroAF9KVx5drOPAzragHlM24QbGiWq+4vwKC5
m22Oq4QU8+ALgQfZx/92gGOoU9s48ry8e/dTjkcQKX4/e/0opD7U98Q5TwJ7RIZ2qHJrRJOyTkD+
YUjG6IkXh8avWZiUDL+kAlAuodoXAQCOfgicY+JEIT4faRgGT//DHDX6DOWomhgxg+oGkzQi5VtO
Ba9q60MRQzBoLhNzsMZaELACaZw0HfjU9ocVqC9v2zLMsID92T3HwiWvxxCyw0L8mWH58ClHl/u1
IBr6sSyCF8rpx5x/duTONGgYHxWQr4OawdcOObpvdWzDxJ0mG4LtWMuh3tDGGlSuJynCiyG6rq3A
qnXeI3+I4Sg2sMR2OGzCUoCFF78mqwmVvbbsM/xP3DphleznGoKOn/XdG+8N3yTe+bPh3s0vZ9uX
oYb/k2iV7qasd8ie6olHregGwUVhPaHN2U1vMLuV2vqIU8aAF4nktLg79VSO6K2nOrEXWOPQyGfN
GbBJK/bsARl0z58HNTy3P7b+Zagphn9C/NcWac3LSaX3vA1mkIzLQFnTIgi6IefCDjCZ74md8Rm+
VmTDk+Pb7xz/WyRJrqWSX8QtwpqvSZ2nS4Q/IJErWFLdToFZgDoR5Rc26toy9Rk1dyDSNmr6DKP8
M4KfM/JY5m/Gi9P9JlXF5fyIivegXZzW5/3m1LC+VvSH8DVcQzvrDj0LNz1ftdl09GXFfReGCL6v
9MUCh3LSjaxW76GXdaku6juzvPQHMopayZBPgafA3hZec+ZD0XbSK0bSozqWJ49UzE3pBD/9bT6S
Ku/f4boArRg46kUvHgBNd/ZEqbxj1CpSRL/2zt2NdoTKa+edcD/pQIybQAcNR7c+FqTl4GQ0xARi
hBdQMxMX2ll7kenohEZ07T52nhX5w1w4kaj/YFUI7q/pN5LTXUZ2s+Hure/DLnJocBR3L4+ME4nf
o8F1zNWhlnwQSfrA5XJSmCOtjYvj6XOG0GkxVD3n0p5mdL5fq2uYfBhjst7+7VEskBD358Pu4X/1
Nh2CSEQD4JzTnRqN1krqMb35g0URilwigEwoK/b0xLxaR0GwgAhouaP2XHFT47aKmlD8TKqIMIrM
uiRSCxGW+sbTAHC/g63pJsXhycozyhBGizEeFp3kn10bi3G7gMSoskvJfMdkpgUyRB4J9hHtjKEk
uIEwQ0V0RoXcrDfxoM5r1KwBTs4PsGWfyd/1omJ+hiCzArms3fg81oYXj3mCCLtpVR+K8lM1Wymj
ORFb0qbUWA9G7WMnCMIwjcLX3jajiim8UALNzk+Hz+4NqvpZR1V1RcMidbvIEWHLwb+UhRFiliiD
FdfORrBpFIs+RDZzOWhS0zMio/jtcbfcAl7z7wqrcfcJXkF8qeskGgMa9yjaWD9fEA1pEQDnOSDP
aYc4zVItQsH5bM2f77h7qTXkDGvzdJcOG53p7DPTmOSql96rOyFI5DYPYh1eIZH6gF2THGSpr8di
HdokhUXS2nHwHDXnql7zO3YlceQlYkcK/Y6D6AquAo2GduwyeL3yn5tYgKK2lKjbcpyMwvptw84u
gEgGDsJCWkEP4m52itte+1Ji6G2eWJo0bzn5cpTN+NZ+Llgbbfsc7Kf7VBaomMlIOFbV42b1ZO5F
9SwDY6RD8vK405xY4gHdsxcKRWz7zk7V2FYgCxlHKaQBZnakgqaPR/jONzxdHBFWQLjPPv4SXHnd
U9gomYW8X4UQmOO5Y3kfj7llvaS2YoaHXtQTdqrMJDicgd4f6fZMfeto5+Xm9z4VUHCnIpOuBO2Z
pwMJozyfxV9+iqsmY0lGxVEwF1FoNz/Jk3kV6vLXq7XVl0TtztwslNPwBsk23rSgja/vlCXFysz4
acflO1bEHX37l2lI9fndSAyU+VuHE9xtQp6FF3eDKFuDbgzNxVv7WCu5fTnqLAh0jKDXTB279BxM
FKn9+cmfG03T10BgJs4AITjF+GBKzycV7mNdMff0TwqjGOFbSwlC4JOddQglWompkKdLLhzoJBER
ab5CR+6vk1PMBxU9MrZmjGcHqxaI5DekhS0sCf9qckHXPK1aqdTCUJnmJEldNgV0QKbVIEc5j/QU
e5ywC/Bp6d85aKqNxD41HXdnCOjMMhF2naTlMY7gomSxlOSzGxgGBywXvdy/mnEHM/PU1C5CJdgw
/b7ok3U/PA5eYtR1v0rGb2XQRwv/7SUGDKNmk6ILaoSnpis+O+IjH1Aqr7KOOCd+kAfGW8yz6CDW
HJZI80GLJ5bbNZ57bG30vmbrcLplV5TE41FHCXmmmQBhrpDatETzlOiCv1t/w2aDU7/wfHRKNWNb
G8atER5TeDAtok+pU9P1AhDKMy4a0Jf6AWWIWbOTAwCsamJXO56t2/TRmRIFchG+AUFMfEHV+4r6
v8UVYnhYIwyZmfnmqgPhsIUZkXgXhf0aKf++WUcnXp/J66e1nb0ZOTUD3hyB54gUMW7AXS92SKNT
+hVNSvvR7uIEUxyS/Xy3fpiP9CCYXMBkIezp/7TiCwCa9ZtBAJ5eOKX8nlPpolPuOr3NfYZ/LNHv
97BDTAkJcAqmAtL6i9DSTdEbjIsfby2i4wOZMfFnsrh59YZPkM421kKn1lKX2HklZZ8qtnXSsJ3L
dPYXlDuGUpNsP05xjBMLD9aTLeDpx2PBwpq6sHhJfCMKAnY3jPmGbRz3ww+O1VikGnfYbxnAlgFb
QuBLQ0SPtaIJul/FSJfW7ilHyLUN/cb0MC+Yn/YnvNhQgPw+gqqPN+F0mQziaaAccw7Ae9Gfp845
eimgQS2A76vEnVq85eWsk/8u5vMR2v7LZJ56VOwpWynE77ZZ8798APMY9M6xBRry8fcKRWna5JhT
a1w9yjJKKdOHRQ78Sfh+ggyT/HRj5CLCvyV1YHf8tzgR1CiG2a2R+iLi5kni5r6YbryCsVd78s3X
Y2qLiLczSWSvalwe1Y0WRbKIgHeOeXEoYkzJoBaXd3uuV/30KkKa7rxILk8+VhJ7Gz5MoxPBDE+r
aKa+fbV8eXkl+UFVXwamGuYZ2SnEDI5w5igOnUbTWxPg08QjEFzb1sGbS1OcDvXfeDDvxoXpcvNT
EQl9jfCkfXRS0DWC9zRiwRI4E9uhlCyj4LrxN2VQNXWaEp2w/pONKKTBFc4obj2OBBGqeva4jMpr
qmk2rRjjWPEPy0R+mWbmBMmDm7czSSJLJfS1VWpJvNuu3rEitJnyohPamyQ0+GW7FcbyeOlD2M6H
enuQV6faDl1peXUcCuGcrSvn+hyX9puHE3/dz+dAUHRFeIS+WI3hdy5Yka8WJhQHnlelVM667PMF
4h8fJNcCP9DDfzD2agJRG6mat6TvDY7Ziekvw+FhiHRy41jVXa+iWY4utVS6/wdexcuBMTEMwJsi
XOO4/NjzjNKVA9j7LHb42WRyPCHEXkMj9jupFi+uabNenJmQ0/Piw8jTwDa3cHN5jcktav6Ek/Xp
ZEDbNE7nD4+XtMQyH117DkLb92oB3APwwm+HCs39P58gZtatBjGFNLZcjXXMlt40O9VcrGzTu4Il
ihfK7p/qWUCdlszgqRRtebRvO3YTJkMPBcjny5+f1d4R4hCEGUZs1fQ1KbvqOABIiN4uOXVxuiMK
iG4qgK0rLwqtj0fS/W3MlZ303sf0OfSgj3kzALGW08S5THpteJv36peo56OT+o1Lqf1sxRE9Z/k2
oQfV0TlT6ysYHLKNexf5GJjyMdPvBwO4bUl0qAWtIY19yrC4BSGy5brI5whUrYncyCbjmadLeI+Y
3AL02cnPOC1wx2xzCswENlcRFvhW9iXA6QhV2YcIx2+pv/nFovw42SjgmrVv42SZuIZeuu1yOI7y
4hrKkiKqfmRDqbe9tcqDO9vga12bJ+Q66BKvFAK70qkRJ0/TjEneptHyH1NxvneBIwmqtbqc9YW+
vfOnN1hP06bM2U7/wD9NHRnlv3OuD6vGXNJ84YQqEFKg7zIbFqkv35pv0jezc8EtJo+q/1PVcBTU
0V2SA2plbtWuFenvf3AraNENiMWFeJuU4guTvOoTYS+EB5HIg+8uflKeYHqQlOJ30uBt7OADLs3r
hvVSbcHy7KjyhtQtLcSTjVGC6P2wuL4J6fn51gTcCCgeEkljPXCPtI4CuxOYiKtsNPYXLZUiQHki
v96KkeVyQruZr0tq4rRn9NMJfwPEnhWsZhguVJr9UCk8LG7796VXGWribjcJes7Shv/RILF7FnKH
EV8QVQ+LBLY+PhE330313hMEbSrKXe5U8m+Y7b87TcU8YAOvGmq/ufGNNcZdWzmmWRDUpXR4YkEX
wU1oIhjpA7/gHun/uqRYfK0ehXPLETyiiz7OWz8EfFiEb8J5rrZ/19rfn7MYHrmbrW9TuBA95EOq
KlAkKzZ7CmUutGPjmjudBELwuYY7+OhJl19Txp8sMkzySpi+G6Bluq54mAW5C2AvGFSbX0yS1r6t
haHt9II8jtrExevVbAO/fRbFD3ofkiGMPdcG2XgKeANIWZkHqLf7v895plbYZHWSzylcmYQyyKVE
SoLDqwQMrLjow6iscsRXY9+hNdMKA79+iFD2NJlCKURg7OJpZKmP4ewhPTm5EJqwLlqrMDO4TcsJ
ALuhCQejTrS/TTOlYffGB88ipy1rAuJl4p5pRB7g8M0mtiI/LuiTU8quyioqifpwBBnQut4KnTFw
/xOYNMXQHJiE0MvQQ0hB18aqB/6l19ftljdTBbiPxl/mvOTsIUYLtVMncSzZxYzldFKHiqafNp6D
jopN9JVVtlXQxsvcaehYoRIedhXFGngPHpXdGH6zutW9s1FW0gLj8KRbRjzG8x1Fvhafiy8CfMSs
ucItQUG4EFxEJWrYk/Eb2tgxlNABjzFCfrhE+1pnckXyhi7n1t7V0O13m8AO8HvFg1/C4hSNt5CJ
Su9WKdXaFi6SAYGrXqJteozDznB9mWIlc9oYdma3Ul6baQelwXLHtoZrWWE6e5Ol6iyD0+iVQESC
0CghBMu2+sPn5tj9VsgbmoEtwkS0xR3iHCyDNqFfVNWQ2OVaA6DtLmXBHu/TNKQeDkyiSZUi7Owe
Cl96GmSJszSjAeU9e/mgWpGLhwACR8QJjWUU9zcEYUq9nqbrINKlSXImEdnTe3nHK+g0AkPneEdU
86g2iuDJhxu72UiE4Mv+I8wFkLDLr+VfOtsWXNlk5+lWwv5o7ENhLhZ14QcG1yHPqyXopE3lRq42
PdZfFfuTvTYGDzQCkpILsN55yvqJK0+mW6sV+Vq6BWJyd5tvG1nD6GLW9SkFPN1yc0JpROfFJURM
u0sbbh81CIOiV1EBKfBclb6CuhuHDZFNy27bc2urAv4uPcrhHFajiw4D+pKTAsEbpk1ruFM9dYFM
713ukJHOUAB2mPq7TiCzjq6xPABuj1JolDwyykcvUMCsH8k3D6w7lDMmMIyJQI1hHOh+0CINUw52
QIJC5SLjt/CD9Pl7botmxDh6BAfjdy8DHlMuJMzdDG9w+NVzKqInpw9I7pKAJyrSH6m8nPyECrgO
f9tlLnrkPJd+i40ksjOmVRmDGqbBh/W8UtmHiR7HrqOOIoAADQRIaG3x7O+6DYAkXdZaQ1iku8DV
X1fPaOfoC5fOyfUU4bgaRFIUx8i2PNniBT7+JeQTdjkr/akNqDWyR8rR7KqkZZN5AzpfgNRp7C7n
CDez4hq4zieN2MtM/tZqk+2LqBlUwCZIPk2R6cmV5l9nJ2a8gZEgLk752sU/ttWomUTeziisvdWg
i6tkFBP0DU7rOPIXdSBbn553mcaSYGFDI/Jd36NHqR2TAr6tpnUnUABYxE4r5xN4sj/sDp7KUOIA
Vawu7ERPsKf/YRelQduCUXqG5q0l5n0PA3rdoEqT1zVyD05BRatI6+lCYR0rBncPADf81MWzp2bz
jSuVLMXdrT0l5Vk4YofwGLttKFs5RjJVq3WRxgeNg1KiD/yHCPBhojD7U+7XNl0CDthdTrhyL0bb
cCSYRFaxtBxteTI10RKiJI4+on9WufdPG6QwSCExE5ci/NRaFny1p2QeVmiug1yVO6KT3H3DxBrW
6Jtsm6k3M+BoywY0zsVPnlkRUWA1ijnc8xEZiX2JHK5PI1I1dENpPz5Ki9lfoUj/V8RuOpS/8kDD
m4FomIvuoZBsvrpO3KqKzwyMSRbGEmnhIMMZbcYebB1RAyyPgspJcBQFU04dIm7vsspqByLH75BV
wfUxBpP6gsevZcT5BZoGAJ2yrVp4N0oASl9vze+YE7n9Bx2e0v04qJh1txuzhOF5+eZSUKrljUBI
g2oiGhmKZD+Hi8CkUmeprnEL6gUenh17lFRSMUuE6y34Fz8OUAaTOlvLr3AIlhqbf8+pm70cnFdO
4E03Qnyny09C8DtdIh8X2S8vzjJFAcudyL3LG5+3ivEcnXM6ageUo2o0ZxcEnQiMGMBDs6IYMFd+
sKDa75sSXaTYuYEaxe51HeISNgkBVADp8CLr/OMU6gl/wf354vQQgYGlf7IKl8SyMSWorkh7huGX
AN+0Uu5rA35tTHHvQrT0DYW+Gz7SNzuNY5+gWcyDcb74rF4JUqfCfaanvLUNo9jSliN6x0X4dckR
wdCws/P9jUFawjlXARKCGyuMd3mKV6iBtZ8YUSZQRKPU7atgujY+/tCRwVmhTNCsnt9uLDoF+ThO
fEdyJ2jQmkZM8zJPzuxNTu9BM7AWzdoIGBAyZrsXXtMyWxyjA7CaLI5OOIi3ZfPoy/TSA1eiaoOP
JFT6/DNfuG+ITr9CjgC3ntHlPyYooWHqL0kRw+Afi2LMDgeEiUBRgKc6hzN3s/ml4gYyy7Nu+wsw
llspB6+O9mtcG/mfM33O59rxdxvk0gwfgsQV3fwADPF4BHIr/KjCL6rTHQiWLp3wf2lhOxv4Py/7
nMILTf989gRh2DVRftE4RhxrQfQQFG79JSrQ71bvUlMMoNMVb+40FnB31dicW6WMML6OLx0ar9XC
jN3pCmxerKY47UZuW2t6sYrGRlCHBnexXmkUI7AWDQBa6r+J7DYoeN/nqoqaQdnTV5vZUTvNlorn
HZJSR/0lv++XwW/cZ9qS0UaSxJ4/gzqCOwBVH4Vz96ni7BSRm1LwZxM4icV0g7W4AmU4fuCj04Op
uJarEQ0vNnuHJhneY7YrY5ooM8gdNqZUPZq6H7EBLBgcoOJvCBB/zdkiGWmCJKVQRZfGwLgQbjho
p9gO+jHUciutYrpOKPab3EQNOb6krXvOOlxljd3KOruUOh0bIkTKIcoxp3PeZDaZcwOopUdSZ5Hz
5C8e5Q43oknKZa1JuLx7swzJP2TNU/CTPjSTfwGrQqjQo19jPLEo98AP/DcXFa1ri6K4EA5aiSTu
+CjbcSPPNbaFkn3CVefy3CaAqTHIv2DXZOruMNyCBkV4gH4cliEa2q4UW1Me/zAoxm/3UFT/IqFV
GBYPdhRqRbPNJCVZUpeFp8Oa+WMXKhOF2Oaz8dDgITexfgpjwEvjXQVVo54qUQ5zmE5IPu4tDjJB
XD6JcSlxmjgzMoJzj7rrX0xAyulyd/D6Lg+6NL3daWPJd28L8SxZzkLf8HlEMo8QpC1s5gDBqSq5
PdnjJVXu5bvJu7+Qwztww7c6NTw12oJf3rWJRSm76S+gZlehRnp2pCU/9xdMBQd0IEHnfmBO/Jbf
JGDi7CrMLp3wbjgyVssgDhwF6crt4yzffZAd00Ss6+eQ1V4YQEyGVr4Tcotp8kHAKASmFCsStJMF
GaF4NWPohh3I1xwfj5MyJVTdhZKuZ9Sm2/L5mZ+g657Ah9XDG0WIiY8Y85BUNx5ujhEeubU33jDJ
/9MURBwFWanB0hsf6eAoEHkP6jV5NXiComML7wY2Q//nODQFVuxfHe8z8o0zwNGyFEu/9NsUegM5
uVqzK3L8rP4daKje/+HRY2hd7UrP1dreBAS5ikltpLRhXqNMEXHmfRdoadeBzVLk/WQIB7aWyad1
5OLOnRxS0379gfqAFVAeiezpajt39GF20Mo8QfgkV0TyNwUsaYonxAUBqgHbOey8xc3RaWO1XoaZ
nat0Nu2hmvQOLtP+dVFiAvbf+OovwjlFxXXXAqBBY2vZCBmZA/zsdWNNJPm+ffglv0XXQ47uZuDc
OAKXNpIF7ibQikshv4lPplXfJPje7qczcy4ev2HlMSZGaAanKK8UAvfr8m8u7fmPjJLjAzZDRXyv
1h22YaslAPJozUb5jMjbQi/7RWsrKLoDkCSsid6fVtna6h+fP9fOkKXYYeyeZer38p7WgKm/sgXY
hDe90Q0XjslRqh+dOYg91zVjW96FR5SlfnIXhSqVqgf61/8BnsLETZ1yW9hn2kmmB4bgrfYtlb4H
vHkNEdtF41td8K3a6ofU6Ig0UC04kTY6bGdgu0NYHHf1VAOdXKr23TmfrbGRZs+xU+8IXJhFxvtL
tjWYF0xR3lcN0jT5KNgTIP4X3Faq8uC0D1hbAudfiPiCQc8SPc9MSLe5VrKJAyjJRZJkcIDWb9AG
/R0Y+dMZ4gKRBlYvGr/daXbRhDOu6XMvq8T4tDslzDXlKVBhK6AwCOSG0UJYk/FXTSLvkmVwlOzb
GA8zPCQsq1NYyekHFOLT4EjsA/OSa46und57BptR8yuZPaDp5hKa3Tc5o0sH9xpf6WLVhE7z18C/
I6Jtv8PC1uXrxMqj99aZHTGKdhvMh8+FuPKVkIwQB49TLnsmSbS9EJoATJPXlVQPFSBLdfCtc49m
Em0BuRGU8a63EwajWdz5h7ZA+4m+nCKi6scA19Y908s86CiAkuBCymIKsaCNcXyOCzF3G5vXgKsg
NKWMXDFkL7K4qQ+cckC+VKNgZBIydZtuQd+/VlRlryd2cbJOltsmWR28i4xDSQWOlDhJeWDA2sNm
oVFu5BZFX3nql29vOSmwcjlQQhf7Du3W+QBFjFsVbkMuknDV27Fv0HHqKIMKGuYfpLZRUetd3V76
qHwYg0ZwxUNKtqj2xCtU3N/DIRw02cJDV9hq4NskcKiAA5IeC0PgyQ8mi8IimnB7BHLochTa324s
st0MgJ49HVDtYnZEdKu4vMX1taPnp3Z71B3+NLAVCLwSx/A5YoXDGrdOqIbC/b2Lz/Osg16w6IF9
iX0OkW9szH+2wZijVm0cPQHn8RvUWv3aTU4dbhgzukjThy7Z+1AEjQ6ye96bhagSqOtue/kVu7e5
TkVGRCywT3Yh6+UFEzqOBnSwdchsgXa+i2DKAsxTpioYg1F+c36WsrOeC1iwftv/3tCHcuNaZ8Mz
a9Gnud54Y/ySv8n4K1nEVDVihmZkKru2+w+2+oud55wa46STt+mY/crp3xv4Yr7MK+6yB8RUiSKY
X6kVMMj03cI/F2bYL5yI8X7DMFOZ120pOB6ZFKygT+XXhh7LSubSAFEx2TF6h+Fls5brUV21B+6A
SJVD4vWgFy9AhtcIRzKZuS8KyTg0LxrHhHFmac4W+uPCTeIsoICdC3MMNwrAnRGJ/dpuqZqCOqiG
XHEjGrK3hdDynR2mR8QS+s9aK6sxUuwZkYa0aZKAlfsDmZG+i3pC+/DPtS+ALNSmaf5Uz056fVEi
5yR+hwvYLrpMSoUZ1YIfOsM9dBKRhsgxE4YSAJf3q8x/FzU0LSr0Z2kTnDwnRu3MTI8ayZM2vhhW
hv3dI6IWVJ6hyRtftiH55BgGSIYqbphFeJNc8k3siSK0MljyuBUCoC0Uw5k134xJAz8Ajbb8syCM
XH7PKwyZx1snwvK6zrJsLtjoXGptsyECHnHSN2qQ6E31Ijfyy6yvblcnKsOtFt7ZtSM1FQYd7jdy
nJCO2Vvf4qP1T1H+mUA3TcEqmmpa6Sv76Lcy2bVT7cgMdLjz4U0x1g2Ic7S6H0lX/e5u0tccKUL8
4LOXtNw5fxXaKONqhoCYcF4sCYE5z/Ep9ZhxXBaOGYF/M721EcXysJd5mebrJzhl4sa78IOkOKDy
CjzgG9YgarrbLBsz9K0lye92WeYnxpbiQ1nzcVgWX30YNYcwh6CEF+wpKIoa1JxBR4iw48LTqb22
2okZJ+/cq/5cj+xjYkZDm9d/H/uhuDvDjoOLGzgFTlDQzo+06wIkXAqszxOzNnTKnQaByX3dClHw
TyWDg0YLCHSybXwUHHuyd0kVNKtf6zsxv7KGWDBNLvQADeRGYwRBZNDhmUjQzCv0nvy6PGPoSHj3
mXt6i/vHc6SUtApz19A8lLBKt0UGLgYRn7ERLVzi5IXujt+kVfRmgW3QmQsWQ0NpePaUK93WTvu5
17ZJSWZ4r81vYJIUVOOSLp9OqekRE4rXxfYUdDDCuupvWplQdmcybyZY+mDYee+FI/mecnVh+c5B
Abfvjma/nvG7y5x3vGSEeuUW9HVihWri+hRCC4F4qeAwyac/cKBIgeWYwfoFrldPbtkVPD8+kW2e
STsuyvpwemNiuwHgk7iFOvnq1DFiuBTPgA0ec9prW2RjBusHTQMy4apj4vzVw1q4DK3GzF2mcsaT
QooxygwW91X/zGteHsx6cRPXe//o4yX+CZrScqr7v4DGqoKvstxIDStVQGKQG8wW25Y381Pj4o8b
a/oSvisrB6RQ+euBIMa0+DcTvmC4H2oiCs5PCjXntybPMK999vC2HmNnl5KEEDqWQuStnTOKBeaa
cre+CEmFzpjtTJ770X8P9rlzgCRP88KXqKJzkqVZMY3vIpvcwD+epQDxHN1DDtVpsJz4GawKFRSH
jExpu5Wwu6Id75zgRKQfHlsBiYKM89iecBI0tum2ojUwRjTV1z0mFnv9v0rDi30V1gBMfvg7U8YK
SCShIQjRDuQRgojqwhUg4e6izUUmptlRpRyTj1EXxEfSDN7MR4rSmOEA/Flua38B7Vjl5hd/+WCp
Uy+lSU8/pBMySWNpdY5poIoofBCWL3yC/qPbXbfABDgI5iG1yxNMqoI2YOb18u6lSDxn8szPEPMj
difm/3aNAlBRLrgfvawWaa5SwHS2tPbXFffAQjraRwXDuYveR5xS1kQ77HCMKPX4IKAYvYXrMWz0
s8wB3vqz6XDHnZKO4j9cZraGWsMe7T99FXXoc0fQBLYuTYMWK9tgVLByMcxX1aESS08ti2PTruzq
b2HWnFmOftSm5fcLd4KWit+HA/4glI2F3OLF3h08cvMFLx0XNzGNU7lcgX46suMdl0SNU1qhSWyy
eGY9Bq5wPBNZFMQPlJHdAjSrMCetilRziR3/Ii7SJnGNnztQYpQw46QZ4+nv9LzqnzQuGgrtGeNS
0y3fA+SyBlBjaJwmT1fYjItdkdozCb2uwE4nyqASRFUA1K8AXDvqDI6yZAUlePM3MyBibaY91z58
fpahYDyV6ICSTyED69BJJs4k8wNnmhzzn+k0g7R53ExxzkvWFQr21YpoYDDabAwTyt6Npd9ECukL
K1/h6wE4LJQZOW8HIB8zch0Ca+PxGnOyWzULaMsOaIvwKNFJgHtQ11cNbLyuloexCgV9VZ17nLig
olIBHP5vghpG3vAezjGqiF9aJfjmvAb3wkuHJdqHgbLY81QTH4ENPyeRg6IZrx5oeAVo2ikfmw4I
d87btn4og8alMcrhtGG9PdEXhbMJ/bd7q6uHuC61fmQyRJSa3m7mhJ3x/YYHxo5dnVaibaqhEniQ
/9RTf6CAfp7kW3q85HAxIFQf4R9ZagS4HFnQFHKAyrv7b2TVsVsrCvf5NCeTWgk2oJkbuAzarFYQ
NEnfFWuw6cc7TuS+50jXiJTt09pWhTUAM6p1DET7o0DUQFtxNOmW3Re1HFUE/55Xf5BPghPqeJmV
AIqdfKPjPD93C7Uy9vlNzzlU5TBTlTgUQ7p1EIAbgow2cZGwbIX0LzfflGZAF/ZUkViyT44eftM7
R4QzL6WBs7LSQGewF7KTOAdqAFGgC8oKVV9hyVFtD8prpaivB7fCcd3gU4XXA7MKJ97shE7ljyUn
4ZlSziTuzaXtxoHH55u295OFUQKIZYK0y7Bn9TmMy1/4t5obTyYsEvGT5RZUU0Gup7/WsJDxKY99
HHbs18gswOjjemCVrSHS6w43TUbQ1YBset6hyFTJwCNIARifvQDvB+vZmVC3YLQSAHGeH9J6yO6G
/H/2pXpO65wDrJrotmplCNnNqZfx4N5yFPDqMBE/JqVrDB3uyKI4ter4SEOJUIQ3kroYjFYUguhH
Tznhdz/w0bQzuYPZvk11kRVw8eBkEEBuYsIURg1WthkaPjtxkbRUdNN3Pk2nyPyHdcCAIiFDkcix
mTme18MQX5s9kxRtc7Ef5NM6F+QjYHrhKkwn4KH9Mld/sJhBDbR+Ztwj+Zqs4LBxufEbbBvTTegt
aKD94HZYMzCA+nP9HIB3H9WZdHv7+sTbhqumgGh85558Ds+0XS/w1EWaEJ5Fj2IHoUzi5o1M0i3z
54X0MzdxR8G5B1BYNxPKYq1pX9SlMk2NgaDlN3ISxM0qbPBLjzez8Ct2dpfe3QaQLfTXyt3iLdPo
FkBTwDDCkhP3l/7LIM2J1gC8VCFrdC3jbY/UOPv1rmXGUz/xnq6cBjqqPyI0By17NtkbPwQBWt7K
OnpXuP2LGRUKrQvNxiC2J5ahJosXmsm1K72eaUndNzccPFuCAtnIIof5FQtEfVwA+xorV4XSU3br
DAell9s+5QcVhf0sxLvJ049szzuGHYL9oAfulc7Kde47g53ZRYDY+YeuVt5+PaUwEWZV30G5sHLk
iyoldGnYS8WsYelodj6qLzh2MavagSle5G/ddW8mDKaUyeq0A/oRjhlNGDKRArTf6d2JFeJPRhAm
avDL4s1rZExRw8n905rDYFmCm0RKmZUBBlbwADSk3QccgAJjiE3A1qZ3U1Ueug9kdsa51n78QiC+
xcEV6qoe6WEVhsTDvFCsISJRPJhwSo0p7zEd/ud/OvBtmVzBsK2PbPQzYmLY0Mb5BkrQOkY7metp
0vzv+nDnfTtNZLvPZpen7ZL2WBkIjqut2yKV3cn8GEgiESL2B3atN4Alsy1LuT41sII7Z5PFCpkg
v22rf9oPpG7xBIhggfHoAQIJyuB2WZx1o+OHIXkCCohlXPIAoMAMPaWKi7My5Zd/DC658MlupPUl
kI5501QD4MfnoyaoiNSGCfHMPGB2wM1rzOkxmgt5KOKLeyDzOe2ftzwvNDkvKZAU/HAhajWkFimk
44liTZfkUfiQVhzqgaeTkMwOdMLP4z5WV78xsRChRm/8scq6GoagHp7o6AAbqtf/lTMKw6LILSuc
BUGYNDXpJc9/FhJXvzJ6JgVz3dF8hMwwcEHCfSAIOn6zHsn+nt9bR1iIziitE9iRwGLLCRBBuyfO
ZOAHOEZ5vdK2C/tb1JiYJT8q3poPGFwvH9bsrXSxjb7ocBYAA8jCm593E5h5y4h/DLq8YiMw7G4a
1wcYNFk/eqaVhUtTvYL6cRGuNy82g0c9A/6X8cYNsJY4xN82xbUgl569awKwbRq8CRn3ItNtdxSC
vprtrfHXGF5Qv7WnPwK3g1ueE/wzRWOyyThhuaduooT0HW9KP9bdHTPBf8V7rBBliHnGo4/+NyY5
yVmtF1CsGjMntiSRkztVLJ2dY6JC/JfdOqOlljjZwBg9TxBQJ3WLh9SBnBsvAekwfymlNu6Dw2tv
U58XoNluK1bRYM0WTG8ZhYtAIjJoEZOF8930uFvqdJcqTKPJAWy/Dz2pPJuLuPPLxG2xnpIAc7ge
32WVu+IAmnOYn80lIZoBtpcWBJrUwweueb4J4rI2QdruwBo3iuUqiMrE7nz08cKkcyisiHIBUha8
FNByNHejpKKTliDIjMQsiZyKsIsaCHWGM2yKM5x5AteES/fCFN5A452MVKkC44C4gDv+pgrQIhzo
Q26EZ4XEN/xvIevlvihJeQUMNOX2+4uwLJIJ4JJB8HSxnJIvm3OLX/jEcZBJ9I4phnuihU0icrH3
cZskoMYqyDHalGpVdwQMqETdtfB4Sjtc1mGGhBDLZjWNWN3Cwow2zqxFqHjnTvTujzPz19TBziow
nda1zC55KmTtIBuz5kHbtxfTj+Ao7TK4cZ0MF2jujM1pCTPGIIDAZGlrKZ7BJFB9xbYawjxFIYZj
eYSupG73sLFH+bpyO3IAcOpbiPj8c3RK12JU4WPaYK2xLzsB2AfhueFc+rLvSvYjtaIywmsyB5nL
qoh0bWLHh+sUbFd+zVfDdBnpMna5pLabfLshy2dm3hLtsBqtQNToNeGMoWTdHaHb4TM2feNa3CjB
U9Q/iU4LB03zJUpSCimKAeEUmP27Ar1fbgn/Tg/N11dqwIyikBJe/nUIFUAXcj7nueTutWRSQyvH
VsUiaEkG1Bz/+E4A1Vc2T/oVGH05XVpDxGb43fFtHFhL8YK5iVAX11WLrXt3Jwk1UcbHCpYtqtVt
xD6k9NLLFqfW8eBbJOYPw1ZRG98HX3jRDoq17pGNLOUl7okm880VRMLULbHFu48nRsKPlBbfET3Q
CAiUsfs3pjISRXgcdNh6qBFwZTcl6PuGeYPgdpS958ByqyIv5hu8XQfO72r/9ZFttheFxvJOyrTU
P5YqxXALtm31DcT1fne3SSPZt0aZxooBxOkdAyzMeEK18GEL5xHaSDC/T1PDWZ1LD+9ImcwUocW0
sKcWt8uxXAPaSqhpHib0t+WhULSJmtvVT+e9EbiQQb5LF9iteCHAz9k0flxcdOBRHyrq5tYCvcLY
R1jze9/PJzboyWvCiyPTVz5uPHjKQjnKJBE/YluaJfTp0btxppjjn+179y6x5zPvm2wacogBwt1D
vdWVBeiH7J6K8DobREqodqomEzj0Czpaik7YNbBP4EbeJgz3fiWrC7kkxTEwiHbxAMFSqL+8IQX0
tj1tefs7CXknrZv3bAGSJF85etsTGK3asLuvAaGNhk8qDf6b7K2MZGXXyd/5og0PNXCXBX+r0AJV
rQ2OX5pyEXNc4FVSyEH8kjqfQEiYLiQP3WP9BjNzCwkQBFewAsJHso1NonZGaJ0IXYW0lIvlzVCC
g0Xcfoc+EVqAwXTon/zkdhn8L5zujMH2VwuUDGrg8LTUUUmL0DKx2LagNYO1DL1XdGTb2oNXr/bM
gEGNURFo6sr/bZgZH0Yj7ShI/gglH9yPz3TuUhcEXXL2W/FJRV8fOQWqACeieugSC91HQPCPYbkK
IA1C1hO4q8vE3X2CwaxCsahfQYTt2T+ORCY17N7qPUgL6YhRLbogQAQpNCG1H9h7oHAorWJ8iOTr
WoXwwfm7qT71hY4s6p2eHDlYz0xiLEupNAB5ePri0fiEDbo7XdYaUPwyUlzJ2QcEHTHrYTRWdKTH
Yd+Wg6em7m/vPoO/OvXIZIwgHR8801VheZPjHw8oAuViasmS7FDMGWrFh8IwRPQXAM6/aDfk9oju
xpmYMrqx0tJLiFbgVG2R/pkTGBUeeF4Ylv0lMpEpm8PyLO+H9R85K6kyCcVtbD8CQEsmiD32RaAW
JyiZnLO4KEPOHlWZMiXbXMAr4hP4/Rr8oaW3n1Aw0eZw7QHJSYG9W2bZ84Yx+gGGlOezBKj/KE3b
ceVFQ7MohCkJyJsUQqAFr6n+7+7VtSgGL08ur4CfjDcwRVptDJAsZPgjaGFhgS/raNZF97b9VVLc
lHut0zebjiH1OVfCTwZLeH1Zq2K5j/m7FB+Rl8LoZXu+FiSsXj36tKh7CVojlksmSPsjenb8/boI
x7tvzDw4abmS8TfYd1l8ep+WOWhzStpVb+q0C40d8adeJUkdbctmWExYQY2OvlSb3Dtd/4fqHSxn
BlZ+mqVVCJ0uzvcStMLlsPAHX/PYjUtoGjgMrbqJ7qC0+MXnouyKSPs320MrLz7y1LyOmGI0WS/G
dPTskGm7YZitH+i6SGmfGYgejNaf23c+ScjivNC964iNB3vZYlKkj+bXO0fgAs7RNKeR9Vz2CtDd
ZO7Glqy2MlZWkv/RYgFgnu+2cylhjTAkRsERPKYFJGnIDtoCgPL6V2IzJXdbvtiaDbbx0/8C4U4G
ntM6AKDGYuykaZA1vZWXzWTdse+/KCJCnZlOnTigCcucixQWlZNJ181zDh9AzJm9YyKGLDUPZZKF
/AI6bQjSNizEhq/uP+fq5CD6edaiKKg0G2rwPvN7sWaPTtZwmvJfNPyK20t1qUDIE9BepS/F8mxW
DRbkfITh+bq5BQwrCVBnh20r0KTSBMs708XyVpfw/zE20KJ7nyiRJoUlFMTn6iTjiz0Vg+OPGZc8
TwBtyAnGAeWddl6Dw6FJo9x7SKIHyUG3Mhn3epLDkyKqjjS2c+5degne5/UmgE/7Xi1rzVTo7lnJ
BBVjRd8/E9HW6D9kCmJCVGdXGP+DoJ6QEFGVHfsrWkonls/NEO6ATJQerXyY5YV7CBV2y6uEdwGX
fd0+K99ptiogjdMzK3UADtwwEMl/mikReVN8XpHYf2vjn+5ssOC5DgwRmpZ9yW3mZ714Xi/G+kak
T07mxCOEFy4Ak0cSfMG4cCiY+y/FvF9EkrK706yxATQKMWWnfQJHP0B0fX3/8iseAoOLj9A/P+DU
D3ybhEzbHu/eqd0RmkAKIkOvIR5iisxolWPpo04tgotHpf6CzsO4w3zF4tQLHJaVIgPPXbc5df0P
iDurhYnaZ6b1bAAp/jDIeX6XkehunzY5h+CH6CtjOttm5v+GAPBiOUXnajX/lxUsQ54k4aTTFfc8
8hrNTopNWhlBA1qlBST3DU/UaxUoM5ErsizwUseczz5sdM98Jc9YFupmE1KD557JhUZbHw0oeA6e
wE+kmhQrNGLPBG3Zj/tIJV2AWPSl5KMQHmT7XViMGGHt0VpwJyhN+tdqCICXwlLvr80xIqbetJsw
isB+7U1xad5sOs1GOYW7Eil3WcJFGP9BNga5137FE2J8H/bH9xw6CuCWbaU25w6JA2JinBoVoHoR
oRCOkuzVC28ZpdB3RkZHGCviqxTwK15rCIfV8xSNPETsoKDEMDs3W8nKOvUlkFVYnVn9TtwtzZqo
dLOMbXbe2PBqJ7fn3rUOl4kg4cWCw2bg15aKwDjOsQTcZa2RPLqe8W3CPSDJXA4RDoYVmUFpKEP8
dUJiR9pASF7tPdCDo0WSw5M09XF3CUoLBwdL1EWfAncPDTbFCew0UZYsxo9QQvb0NB8qlFvTsHlB
q7D+T+ExL122X8sNXuyzJLQRu4+Vyp7FmfUarpwNcpxbJ1uMC+Wg/dncwGYNkY6cbAT2Dai+BJ1I
nL5QUtWlVL8EdkjWPsodJSa01cwPmpJD1K+0Afn/yX2NgI18QWlgEGiotkO7YVy9wz7wpYDAzznT
9I3k2/jwHvyXViCAzrDK5uJTDYzzmwzPiGK8FLM4J/qLNUdyhMSiMSfQnFmsL4oSBKKBO7Jhdgmw
hQaH0mvBL33o11CuW4LY5LYRkKVtQxTZfA+8kYOZjBnZwzP+shJ93jRZJvyB5V++buFgDpcrtHaO
7L606P7fQ4wR9cvjHoO6iK64Qy9TrW3Sez/vqiQAD5DZiS/d9maMSXNuG8KsVskPDBOBiC3Zm8KO
fYOrU3l0Tc4IPXGSQp5wq1GYIapuQ9s7MPRN8KrXqyY2BeEB1kE4e42mE9lk+VAWX66I2uTvtAHN
CVvmkBU797wG8c2lvIECK+gXZ5yGUO+tZuf5sAB3qVNjPOgFqpklC91NMSECljhGqGIWHTdyeh4c
2umnT4JCCUD7y4e3xzyDTQ6nMg0lXqcTiQ9rgQznd4D7XEQmK7FaJll9iLK1P3Qxjp1AFgB3x+LV
06M8REaVBax/g6vEGwCYJgRwBGRpHovhz9QXYwtdr0sBya8ol7sZswsniFmusMu5v6JpRbGWf5o4
bF7Y/3y/Pp22VbZ1jbzO0hhRnnY5KhNd0uefh12LhA+FOBjIknNPR1Ciu0cRndrHOVa8V+SBlAKs
yHfnFGG+sHIZLtSRFYVluW6vXcmClJ90YdiPGTdzyx4pcZ+jNnCPWf2dOgrfYitFLD5HoOJANJSS
piwUVH02x7njf/uFq/DrvZfhuBXTOztG1q++7E0dyhuJRjlrlQB+rW8L3B1GUVEYkQbiE/wH/bac
6xhXFbZ1WvkYE3LXiUDb/5fWGoTJb5QpuXY2WPiZ1/Y+cXfncwFun89fRZjOrZlGmTiBvEdIBFNV
sCgxSjMztIyHJUAcAVwRYlK5C4LvuZHMRlFu++8YjuVleLIXozG2nbj8MvUkZuEA3fXtXZvg3NFN
4UpY5K5tUbPhZTWvwV3VDFhKBsmA2rA0qHgELHzehJEZivCx/LzQYSOVL1NXnFP/LkXY/sKq0Th+
8z3JFmvD1+WitmudI/tmxL8VvPDVEJFac9FXUJbjXoNvjp9WBmJKnILprXOTFwxHbwtf/k05gMHn
1pdXvLp+RJTQE768w34T8jzxmg6crMqz3pjJDbgG0TMIQX2epaM7WC+sRoQHwdwYcEjTYTaLdH83
VBXsaUqHB88HbLYiov8G7Z5pCeAasvmXlS6azmI3Q0FszvYdTWC7dfzSvKGORCSorDdpNlHSYeQa
FfjhRvk13Relix5F1UkFAf6K0ZAU5vSuhlRGOPCDIk0cNpTFwj90Q0P+i6lBV52dSBaC4jmMaH+R
Ii9+faxhLV6iT90KpU7mX1rDpvgWxJYPqrmI8fhdIgCvw83KgfRPvr8rR9zDQ59IXpuwkOBJhTE5
+8pNbpdHoV0XDPnv4t7tLb72CP9cCsQhsB8pv9JyCnSbQNx/k/6dHgGTstO00hz+dyDtXj6jyoeN
fzwbH0SLIliigL64alXpKzXZ1jwY/9l7Vq8Krsu22d8AK9JDexEjo1XkEw1xDROXD5rPQBuvKFgg
qRWPOoOFyaIDbfuX+0NPX+lZ9WY9jSoqQoC1f29vM0BXziOiEJDNSL9Sck2XXKMdlk30xcHhoX+8
SmQ5XMZ/53rMZ4z8edVj6LzcWNKC2qJwRg4g4G3tzG1yo8LIz+A0oPiiuhhne/VjibEoWLxdQdMr
/bRItHqt/FN0O7zbsWC4IG6N1KK1nP3wSUyvFJDMA0XBJ3a40Pq9G6wcGzz6b0NLBVRmcVI9XxlE
mXwR4caLQ7CkeDrw1j54YjHuPpIMVi5zLqEMLcGofn+hXIZ4T+ywjlXXQHUs/QVLjGpIBxOokkLX
H4reO433T3txw+Qz8Xx6lGcD6Ch9MQQDAzwZkZT1gyroWOHyzbH2nzkaw/JzhvC03KDEOloItT6U
0+Fo/8Y8Sod2/D/e5hB4Np75x0U7hzJM7nwUZ4x9BIT2JIG7sosEyvD1+TtXB/IGUuC2wq+XKK0S
ewvwoEQFDAZ2wXFYsSgk4AzyPz76pKunrHQcJfue1BXyLFaLzLunjoStZwHGZMuni0xQUGhrw/4N
E2Jabczn4qlw8z2GSX8Pjyi7z0aUefMbtcIww0P+YcljiKeWerXJb/GDuTulKVDl3NIicde+qseE
Qa3CaTbOuTYwyX43rMYtRcEEQD9ExSuN8imX71Ax4Ai0APeAblj8YGlBn84KSQEwIkpMd4BJCjMc
0SfxFLGFS6v4U8nhsxv5WSnxoVtHELprRHSj95A5hKxKHCMFf/JN4zLt+PZ3M0n+PKN2nLU0RkvZ
HG7OcUnRKc5skhCwCcKlSV7omjhbIcdDOWndKKf6e0zLODEJZkD+pcRHu+4V46h2ZQan26QRLLmJ
AlUdAJoH7ICtMSPRn7RzB06zJZN5naFiFZrzaUlUwvD/MBfK1noB2F0qBiyfPDgLBKYV+IUNIele
2hciDprPZSprMt3h5ENLB8u3J+jbPzvPZ5EHxWFm8hhn5DMWrmVaphU89bDDibsCroTxhyqDfW+L
sG5aU3yjVedZLkSC0tLZMaTGbIHORB9eaxmXYlXMFtGgIUIIJufXYY3lXwXCRnVzdKMrZQb8hV0G
h8HZ1tRmuCyijr9TFl8gZr3YwWJYKpJrtvfB18uyz2lLz2mCYujpzD1SRUd5xoFnnbPR+ybCPs3F
+ZL19TZz1Xqai8D7CPX34F/J+ItbiEQzFOtICpnrhYsvQZOOl9p0hPo7tmgrIpRVI82gsaxRKLR1
LG6qj/swPR3qDkxd6CpCi5JG1OPQGJva4zW9INYFV4004fe7esLaovcNOJIKkgLA2yjRMvsr11BR
xrFRNtM4nHrYKo1N8w5CX5B148sZ92mWmDDQalMh0cwiL1jMD5BukZ3n9vCfQKALzi/4VtoF2h+a
i8mzXPWf6x3RhMSWvw8/qVM14dpQdqFyR+fLzg0qyECwhtVm+EuYdn/6RnrAUos5uVzc6lIdxqKa
/HZgZtLiMz1IiL5SrLuwZ2LOR8+iGrMfoYRBBuahR0SlEZbNKXgoJWNr1CINqGvTA8nupZ212RUy
anHfLO2GiWocViyt5GPCbysFQDbKydT2jLRdGIKH9P5VVtcCJLPUKNq5GIq0GWlGzCCKrzOvPS3H
VC6iWj3idD1gx+zkuU2tatu5PCJRrQYY0K0CdbMVb8njKO7WjX6Caw0xLBQoOT4B010PFSiXQlNo
XYY58Tc/7m1tLmFkBo/HuQkyBLJ+YZxq4UMXo624vuGW7ExPvouuO6HLLScr9IMM1L40vZPDbNfv
6BWQqukViIBjowCoADsIWmKWNPutwfrCmZl1N3Y71P2BLnCLStVyhfRSROb/roXwjZIu48cw98j+
TFnhPXh6bLNNYkppzyn47WwRgNH7BBoGMxZEsU6qLfiFrB/6jQmS9lhUKXilDIIGne0lpE2fMgtn
ALFgKPc+J1G41sImrCMmO4hQfoBCkmToYPARYl40ux3sWsrB5jIODdMhsr8Ao2yXN/It7wwVVHfn
ve53jIbArnutXRovOaGJjVyUpy39leEFKp1DdgjVI/CjhpIRhceIvc9DuKvfkcSXfxujSevRFff/
U5o8I3QEn4kQpMB4WbNR6yvt4tAom2ESYcSfx21fVoajo0XTx445dUwXv4etjYgEarkvaJ0kdrgU
MzNkVSa0I+WKhHyRRYSAImLSnivHF8CBLjDHHTtYphC2d5d4pymZ3tFhYsWCNXp4Y1ia962HHN12
F5T8R6ncxgBwlqtYWc52F5wgaunc1LfAk5DKZd/cu6eZd0qCTaGDYREs9b7CeYMEj9cnZPKPC8KG
Er8u79W8tM59z02XB0AfsetenqhnuOLY95dtZ38N1bLEj4/iYnGmeWawwXj/8lvxHCRWsWfwql32
hZkfdomBecEa9e8JHf5hTqtQJrj6wu5bihVmLHvqfrEjnUKwV15hc20aXLlmhUBT1MJ/lxyzvNcB
YYHNIGUjHAg5XgAS2h/pHdF1EKilQ8DohGaVRGZ1cOjG0Nrg/P0/B/2bjGSzI2EvOgJm/O05Z+lQ
UBVUfEq9GHMRhkFybW15O/c0gQM9SAGnXilK0eZUnMQrRSUJETOQ5/033TZXMZ2fXCfRHUyxWDM/
2cdw2gwrQH2g8nHMyl+akYDUBl4MmY/oLNcWYxVE1H5gV9HcZCQ48BrKrwy3q4Ebcjm+jYG4eqIR
ghEMfUGx4VNLQFVHGrHQsAyFlcuaSH0OQNsHwlKSE9AQrHG0/rXJ4pMixQq+8/9H0eChFP3EYvba
jp/+ajOg7wanIx0f0wLoloA8KWy7LUWKqC/1wCIaflM8zq/mDSghC160Xb5WICH1Btqw/hrZtcfE
NozJVzCwtPR0srGNuyXZjGyDeJGN3FZfGGmbFrKv/FkBK5zDv+7Y/YpP3pR7Fkh3mh8M5RQWbY10
52I0v8EhQJ3l9UsRyaLo7Wl5B1YGuitWHHorefD98I0hFxfu74oEaIXVKKAT1JhZZafkMQ0KEHdf
O7wUkvrIcgu1ddBV/z0IyDTzTgcjJ2Ujozk9uI2qh081425XmLTh7aMS4B37WgEi7uJIRTLIguVF
0CFTmQVMv50/La0wlkcd/idZBmYkEGd/L2iundZ3eB0hPiprBU0LJhOLEqY4qbmC7adIYCxKX+rG
UpndJnLoTJCDCWPSnVB/Gs6JtsVDHNEGbNSQ6CRZa7iwplUDnKUmBxG7hRRwmlmCQtLcxwEueuqH
usryOEAET/tylsLXRPn0xKW9qN/wxH204v4huA0CR3JrSNbZq0KtzAUx2rHf7jDfnFj9jFslLVmY
q+Bc5A4K+YavfxE7M+fcJL2iSonfhbSqGadiuN07yp8f/8uipbULNCvKxstyMj+wKazJBlC4o8dC
y0LcJWtCsEBPoONx7A1NQ1jCAUvA8WSURS6/t/rV+OoZVXn7I1ANPfQHeLXNrqtnRVSJpseSKik0
rCAtCBfJEqlSaCz/UHlfQOx950cuNVECHu0XtuXAFFZfCtaiDlyYmwi+60M8w1C/xA5ZjrO10XVw
6tufx+WZpcFF1ObzvFm9rifLIrmlRI6n6v2ISCgPhj9pzW83KA9QNQmAx7kQeHTOW8jM1onaCO6Q
4KPOuiVMEZ9IdxpEj7siRzQwmgpnYk+SxX2UfzL7ykRFfcR/jCQ3cEz3VhykzJ98FC9X7KySE9eB
wacRCkjPVUvvqE3ibZ98WLShzw0qRl7L3m6RseVIyxfhqmG1Z6HfPEBVPblh1DaFw7wGcKUWGH/a
s5Xf5BjCdlI07Trr92zlW/ZN+VFUHdYECc6Vu/PqutH97GQDgnbnlJ/u82Uj/blNikggcrbY54ju
S9ErmKoGwLwUh/0Cxsiju2eWqjTONWc1qtMq9AH9HE1vmDAhVfReXFsntOt/LoWWS4OeBEwmO8Dx
emgRkAT0Nr9WZZ7q+YfU2aQdqtLXvAg1HW4lqo0MxgR9jzAK8aD0HxePiI9ji4UfffPNJ5sHSt8/
Dwr9BNWyCN/bSJ2EkfAU0ouLub+lN4JkfkV9yXLyNheuwXE5TpNqjMKbxz52S3/dQSgZ/G01DDQb
gm3xGxAlQmW8mHaajmcdn1+vF8ceLLkFleb0AmjKpJEjzxboyDd0e30RIPFIKzqn3KTpGDuxCWnB
+avfjP1+XXCqbBr1Yi1ktd7tHhLud+YqMZ88r8Gfv4rAi2Tm/VRoAqJHYsXOatVhRhzE/jyn66RH
BmQyDOFuunETGp5J53fYwDbHyuKtXrCxrH9YPa3kAYv4/mMxHrTtMICyq1T78eIKL85JFHZRSuSf
4ihXYVky9blcWd8mhok7Vy3rr0BK7A4MyMQ0OmKnG9Al2sD2cl8Sl4ZgIH32FExUN9r/MNmNox3r
KCnrGeNrvqqgydTUCf68Kk3FK8YdKp2epe4qSXEJy9k035aU4jG5cQORpKah2mNqi9a9E+GVfnkL
lu/7SE47XNUMvqLu+qBlUKxfh+vQeVKz2tCEU7tC+msrH4YYD4nWNMfD6szzHhzHfdaLYH+5YIwP
1OvLRFh5eYPEHcpy5U4N7TOPRrwATMzzA9nGaVrTOcX9FpancZEqHU551gAaLufx2L46QJmLIby3
29LfpnNQ6v/kxgDoJxmoCeTRHBl9f/Y7kTYQFDIXWwaoeqUkzEy01MjRF7eQcVW57dx3pN3x6IAm
dUQVfrMaIskdOAISuVhyiTSkluVcyVtwZ/F8fYhKPU4DR4edYZWLS+Tg05gQF68+IiHLD5vGa6sE
1BcrLL/Rr2U1uCzt3qLBuXWT5dA2zDnm1Q8XHUe775Cr/YdqegQp4G1Ykker9gGxCSbYH5VsxbGa
2dOE53ySUl3YpShZXxfrCFytxrDd4WLjyUDa2p+mJReWWZi3kdS+LsXnXNrKamcjWm7JWv9/QypT
WxQV8fXp/q+PqiFmw6S4mNxrPVvuHnIiMz52c5bRZAtFXSHuV47xjJbuFY7mUVfMWYnmc4E3kFlq
LqDFEpK2d9E01zMsuw8WQ64SaxpCQfwJFp0QP+hTYNtAMyDgxYiLJhBIwzwy1Sw7D8AiiWgu9fXf
8c6PXU8MaqzMbmgkZhpcHn88XdyYmdmEsZqioWdlGuHaiBntqAFKRVyaHi8HRgZouEWrrQueh6tE
ipXhQ10XzxX/8teGYpCqNlD6L5omyaryjubRfWKY+dHyZnFPcDfuhp+KQ+dnPulul/VuW4sHDooB
aQig7HLpJDnksFopDU6pISQJr/MzD8l4DAVpNd6gAbSEDXs4aX7A/3kVOr+Jha+Whxiq+0NQ+abV
HEubRgVxKMRp0M8zmOIUfUrjzw0NZVSjWOo3yPHb+wcJWalS0sIRWLjl0Ml8In1RcZo2eHR8Xofb
Zw+eXqIE4uG/q5H8E2bt8Pem8q3IZy1Ed2Us2IkO1vFcmcfANdpKKgpdy4e075049UWkph9FpWYg
UwTCXsZLIqDQ4TI5NqiEuu1SsrmCtjAgNkjjvoli4NzuAk2/XK662cF29V4FgTreWc6iuKW+x11I
7DYIy59L1IPNeFGB3DJULMMR3WSZQV518w9b8y5IT/NzOjt1f72tgphXh97FlG3p0WFC7oAngkYv
ik4LXjdbFyY9Sg9KVg/FfmnV8yekUzhojX/qVk4FoU7rAjuZM/dXrhYEQbjWhniUh4gdZbSrKVet
poKlmQhdp+YaDLsJw0Ym7jBYZrJitkJihDBOQJSIWqX426wzXeUt9CbqT26nzJAqMCaiob36SJse
JgBBGQ1BW+QAnInnaN6OhFBEZKMpzLVPkecK8mJkZgv/63P5RCIp9LT6gpD6scMlLsVTMpnjcyDJ
Kvvv9dhBXIt9gbQnxuhCN9vnCbQfpejjfvHAvK5xMtAu+0sJIwcNaYo04x5IVZCLpyM3OlM969+b
E49PpSlTDPQj3qz+vqczhxVF+0qFtVLPMGiAMP4qKb2CLfV1eqqeuj+njLjV1u1qgUSPYi/16BMe
WL6rXJ9e5rTk1/kdyIif9TBLoaFcLbar1yOTNaeB+desdmNX0WG3RLGjOGcqRWA4pdpAk2cRJ7ij
6Dg6DxFIHHIvgJRwUxLu2ADW8rGX5IO+nzWTsYu8P5N39GaKh5di2yjCTXCg8IhhH/HDRefc+Er7
6xnJo+aFn9oUC6EnMBRagrOyvFp1WlbJL5FyTNxgX/wAGlxXyfXMDXmfY6PgKequQPYI823aguSh
VFbYsWTHxAX3y4omV03uvihwhiLEHJP/GELsDxGwCPIgGGTKVeUunBuyIQKTWnb1MSzS0ZPnjcrP
yytGtB8Chc7IrX3v43thSeLAxNOZVa3Ff/Lm0ra++DI8N/loI6GyZ4aMYDGDBUhOFPLfOj1aAfhY
PQuYZzFbwu6FNNGY4ZEBXLqPFCVjbWB0N5daqdFffxspH0vFD0dZuDQCxWBzAJwWwaEmzEVwNdtY
s+O5QFRkM5NnmqvRFssWI/VZCPEYMjtFi8jaNqP5d1HyaZY5kvy31yjpDhyyUXuw63781qTCzmwt
DuJisfUXTOTOq7nAomEOFtmSewHZMJWnpxs+Uo310SDV8xWnxBoXtkmgpwYETDIr96riGXQ/jNH2
gisb2iXZXwu0IhHCfcT65g7+8H9nI12m+i0R3eoMx3saqkeWsg/wMbbu2O86ScEyuAqK0/8Pa3hi
4bxeaEsP9k5FcYcNG04dLF6QOSc1EodNoaYVRl9IGX/rRjpkjhIIHPdPQgqh0M3Ip7BgkRiUuUrI
IO68LQD5AgnB0yaWs1CKf+MaMJSjpaAB0Yzsv/qtJqUjrtlbqheM0+9JDEWv13KoNLcTQUDROSAa
wkzMXw9WhqxhocbHEXISkmczO1CUusc3J2mwwUc6Fr4oiKxLGeIl8Yrt2Fki/fnog+m54k8Hp6Rc
qpZyJ88IL6Yf0iiv+gXYYmNq8Qj6DGbL2ChIFrFLKsunOEkJNU4RPGrXrxKrxb/CMXgmrbFVZoXR
R9kPRSykMPrGrtPfy4gcPX8zgTozzvAjwwfbwCWWXd+vhgHcKeo/gxTUzkEwoUUYNlQlZSnxeXTf
c66+RUkbLyxbbwMqoxLp/ljkrCGDAVX9Rim8esEgazrM8m40kpWlxsyZlFf7LX2MiC4po1r/8A60
w0KuSDssc8I8HsGqj832K5tuSNTyKKiuWiKa7F1SPt6LXmCgoUMdKmolkO99ZW9bEvijN07FXlfU
VoUSxUhSCNzscwARI+hoFtJkaVRGyrzYbPARdmH6Mr/wJ09uSkIJg9It/GSlqtDMalK79V/575rm
0xNgPhJawA4Vhqc+nRYv9chiCK/KbUVPzg3IVmJlCW+qZmLjEvC8Dn6nA5EDNQSZ8hCBaoOiHsl6
QZAMqynJts8rH6uZofpiowySI14bA4EsvYaYEZ0vc2wWnP/vhXgrxNXp7G2+VXp19zOeb8zp99RD
EuNvyPz78w4P1cVCA0+8w74L6CRKohv2cHYc+cXqYWn5E6g5Ac43BvNjwP1Ri5CbiOSP98Mx4HHf
9+xUz6b8m8Og4dug+BD4ZuW2QkGgEAL3aF+85+HgcA+zc+IB6ed5CV6kNzzmTNgP3wymO0pSM9Wq
zhF0dju3WhN0G4h88KsoQ+m8tJZNHNobuRKs3D1DrLJbRibL1l7sVTiDwPV1nztOx0uHnnZbBQgM
UTDj1WC0KOnftydm3BUZ+RBL+TA4WxUHP6F6KNyLj8OA/HaPevrsVrHDQw+S7j/xJY5ff0pfzGrv
3Hhm7p0396lyFaeaVH8KZhM28kQUUkTW0WAH07CtQDG7KibSWLf+1NaSRW/G0I4JJRSs3009HwSi
uHBfkbk+OXYoqh9uindzO1BnsXAAv0VUoT8D+a00Zo1MzCsEEsI5lIJ4mc8kDDJmezJ6eMKUiK8r
uLMEyxiW9LXlLZOL06G+ggMXiMgFGS3AKjEFvqwkTekamNM4kLasfD2iDTeHO4aCp2Km6CxyTQaQ
XedQyhsb77o7zwmn9aBD+YHFT5iOnXFFdKlOPB8dW1cG15R9kWqBKe+xLcOhk1a20gZ3yhp4S5pG
lM8+6BKOUoWv10jUcDB8YAd1XvdDCjbRaINdlkpmiUwIHuPks9WDat6vaqM/eO1oKzRN6w7dDW/o
CLRdfbOmNjpumVKkNOwUF+hRFSN3aEhSAvPQxAdEBQqOvRtUAJfqEN+2V7wS7YiVY2Jnzz4r6x6j
pgLpHHih6eOJApLWaUgb2qJuxHb49XFi9q3hc3frxxqxAP8eKh9KHGdD3ZJVvVCx91jUagHTRVco
MP8RMAZFxulAZnkN/Xv8TweTgWzchbF4XvuCzdKmqCijzcz03uRBtga/VFANoKQnMjBPqYKhdz4d
v+cbUARbQQtkkhmzfu7grNRV+dsqj8ihFlikKK+8Ee/wGAqU4elKy+6R5nTg8C5sZyCsuWfaVJ6O
fByHnZEofl1lhy0eLS+OZtDxUT9LpqCQvCsY22lfXJFoHz/z2JSpDzfQ8B2uqOqligXT7wYIJw6x
y6+neo9FWIzdOh0NzgXgP0h0zV9ydIearijwgm2IgEI3dJ7oY1v2BzR/RhUPo6JzAMHUnzE5i/ZS
VS43jsljj1k6sIOO4wg/bpcGFwExTmvgHPSj8cgZpiFYndukVT+VgImYn2JWDcBNZlqMXaOq9BkB
br5A0MJVmmNT0WAMPT6dVTIok49pm/1PznjTOVHnxKqEEq7Lxc5MxC0Wz88NVthUZ15oSx4IvSRb
rDhnMZHM+sg1C5/ji5BcKoS+FdxXyCkIz60LsSdlVRlE3EAYY+x36pGU0+s83IfUp6sJj5hzPE2b
eWcRu8y0nwdByzt41whbcKyWWuaar2zFRifv2WwzXBsY5F64fMobeRD3zN0LJZRLrg4Fd2G7lofr
Ra0xmyanhkLBdZY5oexv51zXkwlb2A1ZvHXLCm6oZcevsNSdaJsLfPzurvuTkJQvA2qnT8v9+3d6
M/g4Y8nZmN0gq3I/o75QFrSC6ESc8ousqKpcD/MdGNR/QTtZu6yQZfd5WYLde6kE94WhW/YBj32x
+GR+zlgHcCPgYnyzAKgoeWFVHPeLFK4UT7iuPrTjzrIVMq7PpGNw+GByuM3sQkR4ixuUrVJWq19N
4nGz4tQDaRUEfO3hHMbdCRi91AORtIr95dU/OIJw483LD51mtyp9iLVb8ab4fHrzvN1H6NLpa691
dleB9azA4Kj4gH4qW4f9Dmo+T3Z1pGuMEdT1Qxu3f2tGZBsQstiyU+NtzYzglz/D6gKoBsZpV18B
+ko3LmM9j20qVTmfy0fKGpxp820NUzGZHajVAchyVCdCxKIdu9kMKrw1VbM+3+soGcC87LoQZWn8
ZVbhcpbPLV2KbdUagXHcfSzZ+Dx4Xb18nxQCeSKFUWW/3GsBxTYN3z4vq201lRVZrPESMVS/dLMP
OIQEmILKMbdS3RQBF/JTo5xXCGqbSlawqiv+IC/mC7+HoxavuLpyCl1rrbof9M8aixsnxchnTH1e
CP9n2fR9yx9upKMxwNHrvrJ9DPHWOYqh1wvTbreu3Zez8IzCiOE+Ar7+Dzw2H03uIG5QS/gUFkN2
guaioQ4XMxROA0t5ynjSFgKSkyGTuucLesNHTXJV0ENuDh7aMMy5INkSKeGkO/f6dBJqgz2tW73u
WCqFlPPUVtU8mNN6R54AiDkEa/LHyQK6i9UA7arVb8PMCvGeP9uTLHFRd3e8o7bUpZeWaGLUN7Fd
mIZiD2rhPRdmmbv+/jQr0MCy/MWJr5z0W2nkJzM8QlmpjjW4o3J3IpGc69ZhoY0Miy98toU4njnN
VtV6aIlEXzdhkVVLpL7LT8phb94kGl96/VvTq4Lesf2M25x6XSWyn8K+E3MDw2J9vSXmi0k+4+vr
ayjl8o4C6nT3BHZHqtJa8w8W/9w+Rrk6apDf3at+s5rmknV9SN8Uk1Tk0ZB1Z44dMSE0JiEhmdNa
aZfbEKTF51/7Z0XM5dh9XWIdpTuFQQXBk7l+DiIix3GEx5dGkqQqsBNLHDGKSs3jm/A5zofEvP/F
h5wjX8FZi5W4xzYIaaIBLX1X+hUo8n2fBvsMEYJ8dwh5lvby13LsZoCR6UwFXAzu95lLPshRjIrY
3Gh05LRV0SED8Ay8sdXchIiz7+O6frf1GqX1HxChRpk1fx93C/hfsF1TkorSVvVju7svbRY3ozRt
DpGeXHnLLZ89QjWoBRlwJrWeto8Kkr61QEfkw02Oy9k5h6eevgmWdQaB3eYfSLR0T3t/SDTN24py
pi8srCRnw/6ZVfftS2ZJGJl6YmrCAcFgp2PwxBg09TCglRsMxWAGuyNqEX1BQ4+dwkfEvPqPfFPv
7BGfh5994UNcTQUt/PMOtYp3NdaCYfABC8HEwQuwsn5XiRh3+ZFc7PK5YtteAZ5wAwpaEaSWA/PY
z4rmPKz9ZF1w8rfWNOgj46UchNoZlvv7zTKeA+RA1cX4F/+My73GmH0xMC0fuQErSFZdfWbUYSQr
oiCjhMpgrBdECNZT0gWsUoqbsc6rtjCsXKfkQaQ03+u3FWsYG0/A9ymMRrKFJGG37+aWtWFDjrfi
2k68TN7w5YWTjnF4w1qDyNoAE0YlBz4BqEKqTNazOykjHz+oZ13VIlMqVhQRR1wow1hlbcYccK6o
GJvaT0IsYdZ3Bsd/mXO4piwKy7obEkmIG/BMT3TFgCVpYXazeXPuR8dh+ghFKp6kHuWjcHlrJF/B
1wuVNQy9tfLdHJGsvXAwGkdp3Vxhlywn4Wa3y54HROl0awVPQgnPxg8Dj04PDnO/FraKDsoNQzwv
oOK2SAU1qs0RONienuwtQLFwTAdULDF3fhbFxmjfje1LNNT6N1+LIgtt8RPQK87ppjTFoWeNWlZj
4KsMniAKsaQvJEDkOg+2Stc6fx2O5yL9fe+7U0o0l1BmtW4vr0W7d75gjfT52Bj8EycTpih85lMp
2PjcRYCIBbT8My9lhML+Wb6G0XSuxfQWTPjDnfTEsiCuTHnP3bHTJYeracO6Ueug7pbsj5OzMubl
D5QASOOpX6v7Xau89lwZUn0oom8DUjgERPbGAyPWjUO4M9zz+ijBMVPrTRRFH5U3QwxK2LTdsUiM
P20/qrhNJ834pXfJKicheeYLw3gpVhkfFQ2sn7/L1JSZ6rHinld+8rf2vRW5qxn5ATUNYfd+jobj
tUDkJdR6tgn5ZSRy2U1KFb/oDxfuntk7t63N3hzGc1etmTXsn1OZgdbGruGQTch/25/IKv5gMvCq
lPvYoCq/ryg8odCsYk9jBdEFThTUSBheo/xE6YIM2kQrvptMSZ4kLZE5L5+5e7L2L+pxPmG85FEV
XJ5KKByRhVCUFAKEWlqLks7KYCgqgGMhQfK7i3EKJqN1Cx4KYfbyn1zNqL3UWXhKlL92xwe549cL
MpaMO2hg4S65tIkIXAVpKaQMkQSwNbaO3BhshRljv1pMsxw5B/bFah1Ncwv949k2g3dMsA2RRYCV
zCktmc+RPPHQ/E+04IC3tcK5X0fMFYFnk+e3ZaX2l2zc2J2Xhi5gH6TeATDaWXbAHrv5NyAQ2l4Q
cEGSLeMGsE+x5R31W0ygGKlLHO4LghHJ/8m55+r3rK0J3+AzdKMA6IM06lzahnTiK52CoArqq2fN
XXsCkH8BoD9ZAC/oK7gB0G5ZL7Y/4ZRogkgFnrgl2gxWtxKZW5fmwtRVayVNtHa0PgHBckFUDstb
XJdrZYGjbHXd6BN7E1orb8zoEW7PrklR+0rPblRavNQLTyewhaEtTV+Fc6N/WdtLxnVJlpwGlywa
4MbZhlh6h/JKhKF5fX0kCOA5Tkwqr9IDAPvLjrwXSC0YZk5wClAFDfLGXu6mxmKkVf6IIRFZaNkF
I7igddYfmPQpOQ+zIhFPRLHPzsWLWvF5Db5K2vDU5jXFiLh7FgrheXntsaVL9WyCYzAmdXydZm8b
VHV8Xkp3NrITk0l6qGCxdth6kzx/edgsQf8qRzgt8xN0ittAsEl2G9iHpVKc4j8/UUM+m9aKIuxF
wtU3FD+YJBG+CRrCeXgz7RRuUjLCgV3/0DzX0i1moiFs1HhcrSLTdpri0dwWWppxJyF8MYrYCvD6
RezI/m4Rmbf459sHUkvawRf4FIDJ9j65r1+2c5LXTQIJED0ATy4aGX01ySk0LSEJZ3KMthxjZwzx
18Lyz9P0i52c52ZCVh5jZREE5YG1vDmBKMxlEGuISNh2UZ2BToja1aX44oKlcg+RPX2DULwzWX2C
hSz45X2RHinWpnSiJqYIeNK1NxO002BgOaW5yplRxb/JBLQbqX+PGrJTp/ZwCAIUrOTa+PuLPWgM
KwsTCtpuw9FJdcuRGnc/shnEaBxA0TiLT+v8d1yTipfujoScfsy7pNgA219v9T+VD+4hGdDya9ws
Wn4sqDzxfh//H5tV1IYNqp9DsHXAjczzPoDwag9Slw5NdKcPvKszA9VQOtUJJrsWwyo6/Lt0XYfK
vy9ipfYLn6CC+GulpigsNDdQMnVwxUZlvQdQ8QTmiF6AYi0C5XQjXxseWWSm6RxZoCW6cWAYkkFE
fS6oaMyLtzmNGj1DpWb9zcVdCqdoPRbEKLgMa57SmPyrti9QkyGeYUQip54zNYmxO+vFGROCEp8U
Yh7kFEB3GBn3+o775euOf0IVGatIzrP9EbhCkkFloKv0c21wXf1ZE7PuLRONZLtbSFoDzXSMZNOo
RsGjlgqCDHysFbgZUmFQiQRJytEgV8UsoSoFbFg7VcFv7Qt5rsQ12WlYRJYgvgeo4TmM+ZQVw2iZ
vUYRC5/5A7WY9cJWTJrnnDWKQthCqTrJGZxt8iRwQvolM/L4fFzhRex7ZrPB3WBZsa4qqrFhAzrJ
ezg9+l78Pg58lM47UniqS6oyer9FWcDRK/gyHS9RitzfuY+1tdB522Y9Y2J9bUAa2kw5GuL9PqfA
Z9zO3WqZINIK16lvMetpkybqpwGvX9o/KSSG6zHLj+V4emFQ467frfmKZ9Ddmf2JQGZu19jVPKzz
uqCNM7S4W0P24VPXWziajlZmXz2aEpR/bpgPi/g+bFr82fVsBgaWEqLPk66rfccRyWennNqBhxfv
qAuBJy6//tLJGw1GxHWL2b89+VXY72B2YBC89NiCNcs72vrJYR1HNIOFlrhXMDUH/jf9bdo06JMp
vt8pElNlFYLU+06LpicOO8TMVIyXJyy+XKQ0C95/6wr96GDqIB4C0JV/UfV+Pvjml0Lc0Nb2gJ4P
mcO0JVgMKCSAG6s1IImpNPuweOiqP6Hf4BtK1o4tO9rg6Z5/unXgZo3qV6OLFgwp2cGgxq2qFUAj
2Ykui27/CNOtM1/sRKVLJku318VYf1lToVaqbk66iZgYmL02z2STB/vMw4NW/QgcvOOCdn+JBkM+
iHg+Qz9rEot71kY8WCctL2+NBQhu2ffhlRABkpOSfc/b1+5s0f3Df9Mw/qn9+XHOSInBhF3TEBCg
GhVuu2vxUNKvs8H24daIpmMRZVCZtjyj8GPjJxIgTtWoeBYg2WXM1+HSkDMCzzEhRT/+l8Prrsk3
99CoYDucJgnpe+sksoRVd7+K22KoGT3lYQslDcqO/z+npCBlRF8Pi9ZWXCtOKLGDHyINjT35ZQ4h
en/DxOpK/tKCY3h/blSpyXk0oE3fY/X1JFnK1WkSCDXWuEj5ZKHRp/+PleaahsXiqQdRDmOOT5Us
lvJ+Qo1i7s3fW4/RP5vimQllZPz/IpbsvE7Nk4fk4jLa43+Tco9WXJsurCHo8xVZiH76LGGKz8gH
v9wiVt0xlFJseVcrPzZi7J4JL5j0aHn0nFlmehkHq+hwAzQmW81suoAzgXTkXmwj39JYSXKSZSUh
wMilv0PzzFEW7kHkfSUGy5NXUOOgZ4rt/DPRGojRC9H9SLKDzFD+d0bBVluMDGyDmwv2KD2BsSaI
1lQ5F3ylKBZS6f7fentvLdJuWFqku/qLp3OwNkB5kVGlPyA0kpPvZAgKOL20lReJQrvgO5+zvcPb
h2Q7G9SVKDeKqPcfXVu7r9dGhnbFPyTINHI6fg4MwJiwKrND2Bf3qapec0hixQ6jk/VS6B+EvsYB
j7Kyl9ubvwGXj5YhfepwfM6V0N2Fd2rqWTwLG6LaxOiJDVInCvzBhDLGziy81wK7E6E+jGFasiFp
8u1aQK3HxN8clex3UjJKC8TCQe2+H4jjTK9qC98kU250RFIOeEB0a/R7bQOG0djX9Xhsrt+UwJf/
UE9CvnP6niJEjB/zi0i6n+HmozpAQKc7S4r+e32TmvyzhzM8nJ11iNoe+gpgzzl+6th3ZZA9LE1k
WaZDeBc11oMqIgB/qHcc7LlguCz7PMWQTBUDdZ13p6+xywQrkuDOPmdwY3UIcXXTwHh9W8XKkoov
rdKxT8QtZMh9Y5UUZP8UQEa0YoGvNQzdxOyl2jTUlCXBAy8P/F96NaDimtN/OGviRToPmAJT4m/B
Uk75xZ+FlWTCv193QxpaHoY7b8+T+q2GaK5DdZDfTjJie3cKcgEDyIVgpN4nQhnrbZPlfCBdhu/H
PDfrnsDdQRpO4lKdCaROq89ydfU1666Ww6wVVM+DAC/Zv78iAtIsx3wEUsq2MAJDiS5GPo4JJFtu
GEh6HIyZKx80ooCd/RWenrRYaDR/uB1SeLCHH5AoPL3rZjNciY+IFChg6SG47qVGlIPJjHzvqUHp
VyUJ5kFp9Q6xx3z1AAbCHNW4tsgOPIMcWGIaBOxafoefn+fLsHu7k8xjfQw6PIUrchQ+NakjaKqg
7vfgIjOHy20bQ6ywLebD6BQRMGKIaLi4/BSVZlunO688ZUvMc+QyqidIkOI3BOjTrBD0JGTqVBkQ
idDENXYr0KdN7nW5JGDeKQODcI2gU+NLwA+iOvUFAOAQs1VHuw8yCLcNjHyRnhURbzoymcb/EJhh
gPlNnGy69Bon/aR0d3UYSVWrjjeeQMmbVQnT+ZJkP8e4O+8EAqwG+0PVoR1gwFRXQJsO+4GGM2Iq
OAYhJFBJ+yPJdcEEmWCU/em0A9OWWBE34ka8BkLGTxcrLlKKX4H9VaSaqx2tzVqVteW+Y8Uj6N5C
/rBsn4lkDx+c39+dWLBbBwm1OHJPqD/27xHOtVYFe3ijGADzNm4KDg6iBu2EEhjbHtyHX+zJnpCQ
jLOL58lonIQVKtc8OWOJUSng7UTbvDlo6WhYXPXDwCthO3R+UT9+eSq82ubmqHBVUqoYDrd1yeRL
UeW/SSVYlDOZvTUBL7LpzUNFsh1po/muK7c1PmChw3e11atS912aLSkHu1sr1I2jVdG8uLha8jKV
gGSr68VRGN1jDNoraK6p0RN+QEBdX7SmRyJx5xdsdVKwy6De5u8feQqWHLD0m6Yq+pyS9fQuq/er
2ozH1ZVJPFvWtgKiEn+HPvM9rO+zXjKk1/BxBaKWCLAe+1p7zF+gnJ6yLuibl3MlwxZxkXk/VmLA
/+OCCsih5bTwW+cGcoTqRCyCAsfkmbrD5mwIfqfSg+PCZVd3ZWTQpV2fCEpZG51cTLKHDx4GyZGM
Czy7/wsiA1UybspS/JlDeO0bLZR9BA/OiSLsKvQFMgStIqWRxIeml8TZNoqkJeOlYjBe0pIS54cn
Feg1HdTXbk3o3y/gHXXqrcfY+O3SUkfW4EiaOAzCboQTM4B8cUBb4TzE9OO9vDeUBnw+qIt2EKWo
XGhBo/m6pz2cdkrk9GBn1AJLj0HijBVZgtc1MZoFMWWw52l3j75JgKtYYl1WCxyNxij3Xv7OvzRJ
hIE/x4EdS72RwnyBGo80JP9QW3MRDS21p7AswQCdLIHL7zjh+g2FXTcR5wyxAjfPqod82t96ZOOJ
U009pkpj5/v/4/+7Ep2K7K8d5Ttnntd2lS5Ud/MFyEEhX4SE4XnspTV8mK/jJ4zd/DGyWlPK1Idh
9eXY3cSwXhkrmIrKgrho5A++JbalTBzpWojCBLKZ3entRCj9kAMWcz+nCP6w39yMElRx8kDkvrM8
fAdAo9U37pbx9o/4ojZ4EkiKASItu4UqQxWGDZtC8W8cfItsG9cK6NWcmQmSloEmt5wLJYtZs6Lv
4UxkAVkMMClhy8bT+p9cbb0qr3exu+kNUXcvWDeoSlw3NbVVPl6WXTR7EklWPf7yPKPUQw2UEdBA
Vsb4NHsRCby0KKbaELBd/eClODO2yptwU1I2fRGqHurEQmU2s8ku4QzxUpM/Mw+mdKDQNhquavYO
6aV5PeQWYlgCaRMS/CmSw1jO3+AJW3JnNN0GCYoIAi1OG5Pi70efox1lG79uxgSUIK891lo1Rvws
itAutLNvi6hlFsFGB3iJv3tc89OFAmRKc9Ia/RzWFgLoPcDFd5IQgIvBeFCVIkSEe1oqf1ATQDgf
FLPrztbWlaSlbuW94Sb60QtmLnB6fY8dUsZqVW9AJ6wrTZusiVkSfdz7k8yLlQ5KyAk6BzSEgro5
66/fMIwAniYZd7ykFOdbY5/BXMZ7uayxA55EyhGPNO6nTzyEp/F2AlPZNh/xdPRhHyEOMnS2BZ6G
zuB6DKwW1yWoO+IB8ejFxu+pK8kj3G1eO2JEA1AfcXDhSKJNkZ8UgrPGtWvvRvD4L5y8mYEbblUe
v3V2SPdnrGMLUp3SUkeLReGtF9Z8KOTnXDvdJA+R9mAiHr4KQ8vk/KOqC6Jlo8y1AOZRso34OVFK
yiZgXTNfFSe+jW4CZnop50lB0y4KurIpbDJgXMm3+uO2lbJAUOJnT9/aFOWO/u0e14eUixSPSnUt
c8dTqy7SpuN/MFKHzhGTZkWIY6uie+X9wi4CyJ3ScczTEAoc5vEBN/rzBFL43qoTQWfcHJI/dOH9
pyMPi5oeny3xlkXt/3Cn9710jh70kB45waEof1FfeRbBpSzb3Nw6soui+6FeVlrHfl3nkppa3Jm5
LM9QGYJewiksEuA/iIfh1BnlBTV1tm+wVOXuwOhGo6bjpG8SoGSnr4RFnzni1yDFuT2qPlW/cc+7
T8jOMKd65TDtrmXJNXCH9hML+0kiSpk+SKSs8xvrfWkhjxWTUDTdSZw4s0o9kqVulfhc/uUh1SJF
7e0NpBPtvK1OO+F2puZbYCS6iJsmauPgqF/PHUXXlWtvKIXIc70J9RL1klq8MjEZhKyjCj4sTaYk
NWS2O2EafdR5dftgmpTvsDqSErQPPurtabpyr09pVtOY2/03tBCsf5AQPNeGpDSRbMkBegVs7mjX
a7trbLJ3BNzOjrP2VraIKkeCkfAn64/gizrukpwv3vZt3Hbwa8+jsNFXfmFKtQZBj1UBxFl1HUdW
p8tZjOJw/LO4UHzgThR2+seMbiiFdnS7nKVwfXVk7hhSj/W1NuS5/aZ3uVLQNy/tp+e4pjydfQh8
xO8OpEk4R2BqdBmpgDq/sJOlk5BeTm4umy9+k7XKQOlx/kcUM02Sexiu6gPpxiP55Iz2h9LNeTLr
VjS9WBBCWbvf7stuzsQW7m4MTz5Y/vEY5Ev20Lgbt9vW8wHzvCU7eA0lm6j1m0ZgL8rTSScVhSGI
XyZNZrwHz2jtU3CTGFCDh+2rwyQ+QH50CrS2kZbiN21U9/5eYyndj9TCeIH7X67pdyHwmDs62VTD
cZV29t4KpH1cGtRJ6tjGRt8e0M3WvatDeqA5ZA8r9WcH/5NeyN/ce3ygiq1QzWEUXyTW32psFF5C
ApDC008lvqty5r5TlmHFpdILVwhAg/Ju0WF0538dqRRb3PeJRwBlBcv7apZ0f3kihOmhjSrCkwzK
xGGckBZ5p/R79463kOjQ8ZH6x+hCywZN7oWEFpDya/q34YJczjfoUWic+tbXOuAC8FtK7fLCBv52
pCAmDo6MAzK4ilRGmVRuZabrkRVhMqcQvwaQMa3gd00HtDhz+ZJ18JZmg1nSEr8MqqwkNNySehwb
YuOXkwY/OT8c8r/7YfTFJO1lX2dU0ZMvqTd6KaousaoLHvAmJDmErUHTNsRgNMxrb8IqF8KwTpIv
PjauYHVDfSimgim4yPLA/mxXDRXAZiJE9E/RuT4xv9k6vlWFe5qfMzO9IbO1ps/2dmKzULS5uCsK
y00ViHoJIOItQh4SFvO+FBAPjPB/nwYlj9JpqjjdEdDiHCTrqqwZnEKVycA8NaawgWKfhJNy6NL2
AIBXTQdEA83aens8j67MJBsoyupuooZYmpyIVTxcJfj/12EgLWTAdCWmEz0E1KPchFobtQx+JpEZ
ThlSSy2qjb96IsqLH78xzxHEIaDae/LPxRLE+PAz5DXQ4BPT7dTHOuwa1md4Fzz5Uj2HmROsNuI9
2OhJGqYb/e2gedDdtUzdGqzwS2pn7uKXX6h7ikb+KvjKUVZssnxhrjxMrcDXV6f3lk7ocod7RyU+
OKll9Xr4dOe38UKpQHYQLQjHmnMwIgQ1JKbrnRjPQG5C3RnpwMZHtKdbuFu1rumGDE3nr0bou5NK
N+geEtjsXlbTokThdZ9/DFG0TOjWlWd77PJtIynOeet2NRYcV09GfnXgsgKLvu5NUXzsNBDE0mTg
yE8zvAMAd7r05F57sa/lUvoU7bN1E14P9ielqAKRE/TaxAit47lI75iU9sl7q7XuC7+SUd2RU2EB
NuHaoAb5t7doKrsohbU9HnMkLndV8fT/RLA3vOpIFlecoqayAw9adjfBxNG/IK4J7w6bZg58CVih
+MqrclhjebTTy3/ka2KNl8907JJ7o8bvpvOo04N16bcKXM9VEC7InDyjEebbgVtcVVxIjBWNU8Ma
eC8ZGYbMNfBFUt7l9pDVO3uK7d4Etnc8W5T+7i3I0YxP+b3dataIahYjHB6OAiphGLp/Z0OGdmSI
SpI76ajVpERM7tlX/hHXrY/RRaAJFe58YZybejD3tMZ0KX44dmow7SmjX67+y1KGUXwsbC+epf47
c1kn+e3p9WVNHnTTf0IdrfOFJEx/bomQixe+otq1kKig8cqd8p0wUIK+zYBlfanTQWuKtSt7cS4w
Ze4QJxQ1JSIJhVM8LNjvOLXyJDWReTi/YFHhw3BXQA4C6C/6xPbgEKu7n/YDJpiYiaCngjMCj2/y
tOPae5/CK11sRlNBywF+r7fWSbTFv+NQglKdDJrETrJX4QlaFc+RT48XYDfByYL5XEolHTGKh4QV
9/IXbuaYhQCxxZ15FmPSxsRg2C6NxhUmSfLZSB1iUYOHjet4qxI/DND1uzceBAPc7XnY4OBehNhX
Ikb6UHxFrWj0I+hvjVeGkquL7ivQflP6UGcReZ+JmlPAXnNvZOZWv0DGTQMWYLbk/AiXNhHY8dqo
gzNwVyxfExzu7cHbh0BlMYtoCRDMiv+UBjXabF7IvamfN6EDf0zWGw8qdHOdo0H+kjhg5dfAOWgg
pFs39wzUXKV41VaRW3WNLZ5oY7OcFiiGk2eG5dAy3nmskj/aXK3y0CTp33R5vRo78QZX8xhO8nDY
aBMVSeFLwtxf7ByYAaean5/47cb5bDoMXmkzgjtOaeGk0l7sfXNKnDIX7ymZpwGtB1bvcsyQ3y5u
FGMHc7UEg3Z7vcMvbG0rjF/9eSTmoNXau4w2DPka3lJDi39t8rRuvYpD+m4DWQjVqfgKx0vpvhje
yps+Kttuxskwd/J6HqJiYRJGu2JEXCRLWvpy6Fcrvf2LljkzQnhj2vA1JLDkS0aHeTOPF9bp0zSX
LkSjKNojVZ95320pWjQsfEQCnmMiLzcznlWJJij8mmF5rNdiUbkawljSg2cgo/aX28IlLjM96x5N
AQsx4CLHRU4B7LwrKBvIfTgeciOEvDrIOEAJpMoC+V/7U+5zOjrxXDJ6vlQFX2YfVvmA0XUUv1Vu
qW96r4/MqTc4UrtJodTGn+rJJhjBUZ9Z8FcqxSDQI4XRifBGfa2StH/piBJ0MKPAuW2jfOS2H08z
yl1zsKucwV2kKFz2ajtVRkm7BjQ9Q3PFvQzxZyoH5Gvw9JM1lQW2PSCrWUUI9PxPGtLZOHX5AEMk
veBSj13sFxLmvdQQAIOwglKtA0SG3rvWTu6eggUDOLcnFwaU1EByQqN9lRbLx2/Vd4UrCEGxadQg
af72s0j3TtI7yLaCoDdOg0+EHorrV6B6wgFNo36vewdrxjo6XK3abcpoQcB/XLuO2aLzQk7EEnL0
Wtfwyo7e5Wj1bplr/JRhWgU4b4CdmyGa9j4GsgjUduwbEVKFUDT/aZ0rU5vhwSqAtIgY1KviFfIo
B5tYrMWBs4qFWHEZQ1LrYGx8oCXkKQKKRV4IrIC+heQWbfEgjPkJeVwxsawOf6LmQsy0ElTwQ9v+
Cx0HMXXjfXoyNPRm8F55Wdymb0aSkLDtIcTeP3gcyox0L3kXwcMER92iyfqX6BVVv9/xEHcTzPYg
4XixdYQsUrhzhKgo+KHSJ2YigOJSjbGxTMsAS81l/Wu39tO8pWfNwp58eS+Pi2cbWnEHrx3vc/6a
kfbbjO/F6qerQtaTaNyYgmE+QMFetEgifm32rLX0STBHUjXqA83pPOIDHAIcDxkoRUam3sezClQF
UyUP8WcPXBtFl4L6mBD4wb5TDbT2axpIX/Ly3RKd6+4JCeyx88ta4NuM6O++2rWQSwS5TGPu4dX9
PACVej/hFd+WNrytT5d1/YTmhY9u3ws/FFtIQ4njlEP/oYolM+GVCM39VryqEDb6xvAlt9Q2h3m2
w2yGlXI47DzucqMHjGy/Obj2g7R0nne3EKk49TbG1swJvAdPFgZT4MxWPN274X6QtTZdNjpKw/Rc
Xmqiy0OG8VsDQmG3+OCPosqWVjsxsy8DGskkcgsqKPnJ9kJ7OHK3II48WWzSnH0ycTXpBDKxt8UA
lXp5BIIwYBCH0p8acs2Rw5BRF6u8DDLpVBGQN9RUxrimPvNVcdiURwoMTUn5P08XdIX6dngICBGL
Kkb83NIXtX9pdpG/VOvO3L5hhUGGNKkNex40dSTZAmajwjEGAIHc/Rd89bHLhzbppSl9Wzsd4ltb
goOTGlq/GmOasbwhZm7N+E6T5Q0Ja3vsuptOfcwhnKrEhHa0Fs0lhHKHJpBRUj6U3RF8f6ytg69S
f7ofgem15IWVjc02YSEwM/xILuUOY6dzrHVCGFM4AnBI0DDcywiYVYxRVnXnvrGh5aTkuMZO9wyc
kDHprI7H3873BQ2aVBgEi3RJEQqIqQXWI/8iVFmsW+N0dBQWcVOLjRty0x7IHtGQ9lmS9tUrdCZg
B/XhPysBHzuDbRSInPVQyfQV03jMVy789jeKkDXKyAtnHOUcgJzxL7yoC3PDf3nwdLB36VgMEiPl
upcwTdDRbyVbAh6e+HESsUeWSPL2sPLzSfafKMhHNTRfh7vELY9Z8P78QjtKf8UP3V6McIHQ0bYN
Bpbj2TlDHOfnFSR4sJPtWzPwZOcPck5+WMSGr4aGYCWyMpp3J/g/Ts6vpXwg8VIQuM8UBMqGxsBT
mcvX8deFe1DF+0sivq1glfTIvduEV3U9J+QG4pycY/BIsEllyjNf09WGvjUOQcxTx8Y5TVbo4dxX
dLcWI/ouPC6a1jOBkXUQx/9BGMEY4I+TAJd51sEWGpZ9ekJAOAgp3qDoDtsRRQtjAfc1MhIriu80
Vk3/w6rY4xSNaR/v9YGDL2Lha7arVEkDHMc2ryZVFuSztRrLd4Wq7BJe1xoxyDC2tcSy/XcE9Txg
h2kdyy6CAeZDRBKF+Xo4meMuwpitQ1E5MY/sPNkrIwe+O8XgADBfgZKs5+QIQWOuTFsQnN9FXaWb
qd1sn8w9p0ucJ/GZ6aa1p7dpiGdWKv9/pqUdvf+h915J8udXNK06/tqlDepZmI9/zI22wutmx2xG
A9RtJensvy32I9OCAWHbUF8yPdOqn/BPYgifeRN6LdlKJqvBadp8NuXafl/OCRcU5fHAdlMBmEyM
olNmVyr0zD3kWU89hk5SchchySw0MZRyPbE+ygzYikaM04A8Jzvr8dm7dTxPYGZeuoY6wVBcAdrL
SqkwMYBJ0r2jRUzn4TyZLlNYlzJlsbHNpYUQJQuOaf+mF51ag/kNpERg8ZwVhFJ06VFfkhT41jp4
50YiXddoKS5D04oYd601ZbF3QjWiM8uUQ1qHqaVCDKdIUTx1nGYVOSjnL3PsdMyY4XdgNstAiUIM
oVWMEA2DwtQhKc6z8FW0gkK1sVarb7IgO10+4B2LvNb1BgYCbTLlSc/jzgsZ/RDG8eQiZksm3tcd
Rw2tOV7Z5Y137QvwxBoHhfCTOrS/KN8peFMKX3qNNy3MJ7AOIZRuJ52e5laR0YzpPKEuUlWBhy5H
7RiOebDnZP4X24AvS2SAkNWx8p1zIaNXxv9AjM4DwP9yltFHipLWLywx0MdcEnYWbHOkYkjGQ6kO
irE2jAGzNYGWPAAGZQlEDB70LxuvoDYqCHDP6QVqbinONBkIN58hrtB16JmWdlj3avrHm7JkmYZ5
EjOZFFzEOrqNeAOM2XfYcENFGr3apBlFiUsYRPelE7gd3YVUCU9yETKFL0D0nRDJN42G8yvhBNn4
Som3riIktbGb8WqshkJ08f9iO+J7g39gmrPjefqr9NgTAInq3JfGjBiwOxI5GYa3GoV76cGgjR1f
LNPOQ1TIUrJHxR4Vb3S4c65Cp9QtKHMdjHCINkg+BvtTpvMc4uYXL8NEmgPzK2en937zk39+l0h7
LbqPlImo+GNw1L5Rhyq0TF1kLhaK720zQPE8V11/1pcNi+Vt6XikV6ZC/z0sievA+MFR79+WSzNJ
g8HuXSDPgV4HUu9owis5fVC3utFAfsRJjUASa+r1yNGQjhXtVjyvdk8sD/DChd5nn5oRE72GRmFG
sobb5Lm+dOfB3xjvjXu+r2v12VTP+m0yCO5NjxE/wYErNO/ZaM4qEpd0+4bypNWQFs5mFcs8PFp6
yOvpIhXXv5xM/LMrctU7eLIq56GRWzFb4BZoua5Md6RuPA0BKEWBN5hcBxuMdbtqoOSPTK1Z+SD0
vpakfDjSpvNNle+ofDmjwQvC/ffakymMLgjTtvvPPOIhE5aFBB1Wc4vss07SpkKsn9sSR35VTzFT
QIENe1LMV6T1zNKcAhDCEMUOcrwJOUGTzvYX2nN9b7xA0HRkuLIaH4Zy+h0JKZ+3SC58oq8T8atJ
flF594A+bAgawZRf3tDEpubtaI+B/Y3IYrpG8svXg2nb94wZFcFVD+YSZMxBj4eNO4/yP/pOb6Pi
d9UYrHdQtALgXedXM10X03Kkh9lHaMUlb+5dj0bQnVgvyUtVafCbCItylSUcYlcFtpi83VFZFlHn
xgMNhGT6VeLcLMk4kyVwGE7By0DNUJRSIwA4PIT/eguuQqwFW8x93dC0e+4toSgyqewOlmCoTdQR
J8MAsI7SSJDUW+IE67+v8jkKKDnfJtyubUsb7gYdtMHtJvMiMHzxFvl4yoeOBoOyxWAYN4fh+Kfy
ugBrtFg4ko/i0SijqqWf9s+pJ4i7EuaUJtYw8KlSu0rC+Z2ZkbzacvEs7doJUfn8SS54Bmr8RgDO
1xP7VXtTf9UmPPBXRDc4nv3klkSNMD3XSF0fUo6JabxcwS5bOfjLN5d7/BK0ECD75Ud++pLEw5Yg
HmWpFYEyoubIE6pczR1bj+l7aBE3ephKB40VNf0jTqZp0O9EkNKRAr2ZBZ/2nadSH+/LvZ9FBDUN
UR9wZQcarz8mn5OP/xMJV7H0YaucUlrp+kxv4SuxdIibf3V6lzuA9WsVKl/28ilrhKO7t7FSoW6/
lyx+3+usC/6xZLd9XE6mz1BYqrLxv2+mQqDZejnb3MhIKLpapbDS0bWmw1Q2veDFzHi0xu15szza
ImSo0bvuekgIEgRScyT09AWUYN1/67LYMzwBDWV2FgwkNDp120d5fzlXI4AuHAUokJzcU1EAxQ66
jwYytIlZCLkkiG/XOG5z8EQ5Rlm7FF5RXJAXkMMi2Qc3/STIcRJwsb1AWh7npz55pmPj3uvIjNFq
M3LMt0F5MjZrSenNmJ/4LM4YvNtXuBA23bf/cJ4BZDiafp+vpm6Bh37SOvjmhtXaPGLlrnHwQR+q
FB1eXVX9IiUkZqILBkw7P3QHf3EecJ2LNn2qssPVYvQTAEV2YQS7Xtc9nRhZKuvsQ49cCjp7sVGw
8pLhI0Tc0BdSOQVH2A0kEwD+J/b21qZEPIK0kyTrS/ktzJIFzcgXbq1DKqYTBgfA+xCsncJXuKyd
7mXS6ZycekFD+VdTo/uZyvZplfepwfc+UKqDEEjPFM9HsofbZ9AOmlHEdIrMpORQ2RKaMBt/FqKf
6jqgVYH/XWoLAMhZAJ/yMUg1gBosj24z9UlSm7qJK/cHq62xaBvzmm+LZaCR/vdvSzhELvsvSAyS
FisWmVYsX9vw585akg5OqbvAQyI8tgdn2Q//HesOI2cjLhgSxoiT/WO12vhFSq1jXVKr8N1MxMQY
GTn6DGFofrQXhcLNznd+2Jnnzy75TRmagxnb1WutW0pXuwBh4PSwmgcAExVQurTybdyaKkR2yWpV
VqzESDN1+CZJ6/YL2fxdcx6tguNptgREtuHq1Uhvb6+DeQZrYA39EDZ4IUB/IepQGahOA+jG8N3P
avo7S9em1X/oW+W/jF4inTohSsa0Da2hIdo8n7Lq/qXgVWw0hTR85ewbr0kbtSlP1ow06uN7Uln+
Drp/2o1J3orh9NF/T6qR5SM5UMgcNaoR3HsUl/OLgH/UeHgDyp+7UhQVFNEaDXX1qF5kN83KsKBP
W6T3uhcQBvXHu53ig7HJCisV8K4PIgP0QM7HDbtRWX11/U5m4R/CYUqTY5BiiVd3/lpqErbPTNqY
+N8QeH67t0RTlo2nXx0h2JmE8Ec3lL9yD6XeNa6Ed8ck2IfRlyLoHe33ZAn63sVwJt0gxJE8pcdg
ccAJI+WUC5TrxRfawzt8XcLiDotGLRG8KT0Ms5RU2DDDprHqh8ysQu8Y26l3KtmXYulsRKgMm1Jo
Wyumd1e9xGJeC/B27bxH55HmRSVVfsptWfULTNpnrpprJwOnStMkvBHKFNuAqjKB9jiuckrMi/xA
ftbTfCNHag6Seq33xycXcsFPV5XC8z3iGLvVc+nLTJWkzBIUnQGOJqlhIEnHLfjQ/VfCyGORtjIq
LsrlTdO0N1eYdNSNUkOpNWPvF3eJhicZr19W0lBVLC1QTFpc0wzDJjyf73cgSG286aHzCiWCtdSq
urF61+J8KU8I3Wev93UHKlwhNVsE4OfSQf5gHbFITJrZeyvOipavbGZ7JBeubhhmDJUf2z86q3SW
a6XTG17uQGVCYYV0dKZn2uKI/ncCtSEFns6tJa98uIuQC5MVEqB65/JApkHud5WVKziJq6BsNg34
vKPnwT3IM9vj2d++tPpmZ84X0gLUQWxeRGkcr4KI/4/RQIZxbdavkRQiGA7SIznNAOjEIf5GlkSa
8Q5GdcU2Sz5AnSP6eW+X4IiliPYtVHaL0mg7lqOe7xwQ4Dreufie27P4B00W9eHvcjA0cS/50FTA
CFLXV8qciHb1fay4F/G9RPIz/271cgbTCaXO1jG04yue3pghEOG9UKj0k8vfwkQVyA2fAM0+kDbR
JMLoBhfO98WKCXdyhMoot7ehsktA+x57zKAgQco03uS/LpJS2pfvLRaqxlhq7CJKFSiOKKp0EJiH
o3uoS4WYAzy1IFlM//PpAfKoVCExMHjlPO6ZgxUklJzSqFZbJkE+miADc99ulq7q6hz6q+UmxM/H
Yfn+wg5AD70j/jpzoHJzOLGwpG79E9fOmx0oeYJLrjbcCzmrSl8eRzJKRWI5hAGyrqa8YNLk+irF
r9/Xq5a6KUw/O/WlxlgYp4u3RVkTpep3sPzSeYJH7QYoy6CoFq3MjSAwmmqCITH0k8rZaPGSDFnR
vAbNpZlt7gRJDkWuHDDpMRKJ3XtfOr1VcXO1tKq23qDyVAVW0QAbfW6KIYEvHfoN8c1ZaCH+5U9U
TbwiOswS6I65Zl8fAhOOkMFO0RuaTgKZunbrflVkPONP7CtdkLjO5r5XjrASJt183HFYpabGOJ/h
abwD6LD3ahehY2neoM2sLToDsyatwdvLyfGjEqMziE5X8DfWoQruImj5JleIAPQpA/uAGJEa5dKQ
m88AQUmftWijDByPk3qRnA+cNcGvDqiC/Ac6SZCmCY2uJQQ6WpilJpiTk2J2AKxz89ixsLG05+FZ
HaFQvT+tYXCwDjJmzkFB8r6fNsNsZpnoyW3L5NQCeI2l7md3Vw1szpOMkipiTjgkSv/gx77mC/XI
pHebAl5Zd3qflufA7XwATDXi59IlA9m8f6YBiF93MUyZ8Zta0sSiJBtsP9KQXBRdDBRHitKVc07X
RDUhzRXioPc961+abH6b/q5MxYM1jZW/eJGxSiYriLq+mZMlSW/EoFZG3rJrEXyOxpKu+WZ4fj6s
ACQ3eMyUTsC7q1DgkRk6AQPvRy070JZGMfwY/HFJID37QqmNaDi3+1C0K+GVFHxxa7I1LULPb++O
HPvTbUy3UAstIITHz729E5yLlcx4XKv5xkZF7d7xNPTrbBfBz+cjP1VLO0Qx8B4bGSucJvVSXu4T
HQD2bYj5e4fRzLxl2IRcq1lsD0Ezl5udLmRk1HHhJBqPt77DRvelUjbu/BYJrTfaKkmd6V+vFV5J
1gySJJWm3e3y5iiXaaxrO5e4cB/ogEISw0bNGSlA71RbR5mQ4LpNK25eShNMYO6yPwU9l6yYyO3f
DrcQ2KgLNJ/tlSpmn9FJuF1pgFlYDPPc2rMGDNYzywx32hrUA4vi0sZg8HqxVzBTaPjE94EeIkwh
1oMvk0KRk2L74NN/S7q4TzqGfjp1G+beH8isEdF9P2wwQwGo1W0DuWAPYhQ3tqrbdKGUE+z/Z00v
+0WcTBHtkAieBtcv8iv9ird8SP2+yXK26Zxzy6nVt6gyCW4n/IBFy8HvkhPiRVGI3s3Esyhaiwg4
cfyjpTRWc5eC+AZ/q3PGkx9XM6d2jNQA6qFowbQXmoLFDjNpJh37RRDYu9oeFmzj9eO8/6gkfnap
6ImpqupOdFLuW8H673mgeBlIeDJ+b3JrQ0Ge8XA3SZTU+nLRuRifV9OxXP4WnZnqqU5+kQsoQga3
26Fa7f6G5W3dFvQeAjOAzkrBUht+o86wtA5pBo1TfGJfmqXdqxdlicA5gJKSvsT1ApAm+Lr0cQNc
bOJ6pghGXfwKMBg/U+OGj6nscQ98XJq11TU+wH3OEUaF+4TWY1r8qIz5liyqRAqDyfe1R5heOsBJ
ZEoiGjOvtMi74CJFhaMRVefeYgpR+YwK0Njcxn0UdHrGO9vCVFrflM5NtJ/n/r6yxRRiCIvz0Bzd
4R7RlLqeIR7WL1XpLgCwVc9+T1gN3asa/CGElYJH/UMFGYnktiQ2pPYhoamtgN/uxkSH2B1YOqC5
U6XfkxF53fPK0Oeh6pvv7i0xIl9HOkzCYruD9OTQ/9wJM+MRdieewfi0Ywa52pska+l/mWJQqqQY
t3jaEG9MkSVNccQWjzzO4oj5a3rzmoWP8INaEtiB3GGoq59D6cBjsMtqzUSQwhdZjWPJ1/KRQ2sK
U2rFtYTZ9NbNMZdF1UBTL+KnpkuBqy+vLVU3sU65MEe60Tie4QAg32lxYp+S55ysvcVg2ruFCV29
rNNbwNd5NDoI0ZIpSm+vxirsAb+jffx5lcBwdkDZqq04oxFAGkMTmEhPDqVcRSWuMLDxs7eIS4eY
KN7+EX7IKEBb167Z1BkOZSXgFgzQPc4Es6A6fHNOqOJ/Y2RIWrBN1b4xoi4fAlit2MnefWSDlfiR
nCtKIL2/1rMYhn78qGCSEbIBiJlKkEBsBVjkIbcZGBban0CdjAPEzQJScXgCvfJFKwu+dwIuEATW
ovFvsUxGB/Z9v2UsJno2YqmwoHK+NPK8LmcXZyhjUnrjpd38BgtdSHVlnKIgTXdll6AmKvEqTvto
Z0R1OQbs7GL7U+ThR8vl0M5qxk4lUUalpyD+Sz7MDIXVEZn2trzsLTjlMWNfGSgv1P+XHLwD7erj
9M8ev8Pk/7UpxQm5no2BdBL39QIgxXig68xo4xSIOTRG2Ok75N0cPMpyD98M0WMvjk0sqV6Xr5yJ
T6ciePQswiEvPzQ2QfbfJD5LEvB+pHQF9Lcp7CvAxzoZaNvLoFpxUuXW0WDpWjxIzwzGZA5qmDXy
0GjQZsupJ1FNDUX5YMGxQlsi5jpD4skmokaQasYvEEJbbgaOz26r3CUYRNA4q3nyIhcz2JJtQhMP
VIYkTJ5r0X9GjiElqje7VkWvk5lJpZu1znvLkcGKQxBc7KjUK1g+JH6xKEGgcHI7gfunLqvzTnq9
mtf6M4vjoqvwRBTPDR5fDuAEJ3C+x3sa1XBtr3mSQP83aEBVARKISAF1H9AIMXb2hzOFQuCIJwVE
elZz9Id9tfu3a2eq+qhmdzJhXzo1lN9XP10X9Ixkw+FRb+oXbGQM5Rd5EKkbWzbAxcw7EFbHonVw
MNK6UR3FWE9/NqZweOaJyRa3IVOWE8TAVt1cg9s2IcPW4ITGiIe+emTp28YW1xYK7hTU3qnR4kqR
PMRNdfXq4qfN0pehGmw6mTs4eLC5Vsd8wyyTw4U3L7SRhdr30wOzdahW3bCFU2RCytaj14po21KE
rOAGBkR7Gt1+h4awouvttz2afQUIh7lQn8dCrC2ZaDmOotOMHGplj6JNOm6PrOc5UCbsjm3qGV8N
7RJY+h7xMK7Fud9NvECC1T/0G04kGTF+7yQ60AiYdNhnp6cDcJugIblkO/LcPBozMr3pxW9oFM0H
6Yac0M6u4t1u8r8HQhq8bVRMhs9R2Ei58qElBBC9lhvBHueZPK40jboblHVnDJRVQKfRs1L79KL+
Ta7bvoqnVrxDJt90xOA1p+9oROYeMSfxWwA9cZb/CIC6GMcb3hfUz22yXpzNkFBXNdwjWnWVHZVG
9tIhN/X566kLF1Qa9HKpNr9ny+uVOBqqI9TtcfSehC27WecAIxojmfUSu2/zwC+Ku46ga7bNfNiZ
pFk78ij4eUIvTiWrs37k2k9ktqrKyB3D7upYS/IdJO/yWyeU1XiOGTrZFKqqJffzyM4OG/7AvSnF
2O07CLV6kk9hpNxw1uHYOn5y0ioqm1VBOEUdT5St1AnbOPF5OEaCjIMZjk9+zgbi9jTjz3BAtmQV
AqwhUiAayi4C6IUS54r2rPlLyaV0l1qNkHNXPJBXQ0ZjBEt6a6X57j1j1oqUW7B29zsYYsgq1ky4
NVqQjU4QECYiJNn2amCs1sV7oq8zCt8kjTVKIhQFE4LisL+Vi1dnCbMKQX8yMFnG+25IN2avMcob
HCy/XDuTuyy4dIF8Bqub+lr7A5nZUZzuKu7cwPulEipuPm9R4k4WHKoyk3/OzVWOPRQgkc6kGGv2
R7w2DmNFfTax0i0fRCTXSNMv3oimKSc5P4iml+YSFh4UZz8YtNwKbT4iUGPiRO4AjUx3yQs5PWIF
svKQOupjUgg7ng91ysv3mT4eDL/884ZLubd8QGjoB6lZHH2z9Sj6K6ZcqZXC5K661vS1h07TDDUJ
F+xCiUY6teJqSosx25YOf7/GjS2ybVYKQ8CAyKxhUL6s7Xi3AwPuHeQ9U4nJafmtQiXR2N7dTZGE
uUqjsdOiQSYT2Aezuw/w5bMlXlTji5QTShPNfaJWlbGEaMwptuIdQDJWMqukPI9GVDGhUlbkOpEA
OZaYb1XmzGofwGOEbSEREN6GqNRavMnzEeYyms+I+z/i0xYJEomKhtQYjo+La8n2Ez75ZHbX+872
PphRCsih4CV8sD9hw1rd72k4e09Phsb2GyN7J8DRRaEsQo71l54d1gsyxnF4jPXp0ncSSWspOOcz
rebZNOXbdMX8Amfb3bEQmywdbB0THm4Fn+bUMllLoWuvENcDr2xHyoiqyvFMisapvf8Gjwj8415F
aXOGTfx1z9HEFciWa8OM92RYRkaczGv+j9FIfB3HRD+SccBHUIG8raNiuXFCgOrMD4OSfrCPGU7l
AQ/Vo7qaN/M+9JdcI4mJGCGonbZTSyydeKuN9B5nnVD9lYWrUK5REnXfCPDPyv/zi9RC4yCQ4BKX
Ft0MJ1ZrOCao4r1R+d2NUnZpeLo5fpZuxS2wFbfrfe0PpFP0ikKEJT3yO+MheBG7ECBqaQW3DjQR
3EipXRj6i5OHs4DvXw1FW8P2bjWKaDrRdBZjYNCsLK6uOxxpkbhE+7wAADylAEI/EIc56p7aZDFi
VPQt5L3NPEk7ySADoH21zM3hF5SObDYtLjPALFxaaku4OHad2FUUacYR8PXvrxRryI5yxkdZvSxr
sWykIuJlI9+0DFYiS8NZunNWmsd05zxVc/CztFP062vkxHSEzAC0BvjA/Cuj5Hc4+3rb8k8PzbSU
yX6nrpE0Wo4XFUeiJqnL/jBRjlRsVF5SjR0ANZqGkschxArLKT2a8aRgr3vv4UFJOLMMqJ+Kl4ls
LOY/EV/b7Y6La7npHOWYeoa93u8JjgXDJNYfFfmrkFmMLCzf92nf5tywMfLk4mQz9/iX0KZEPEW1
EheM1oy3sC143ui1WkBTo2wNHY2geZHuQ5qxQYDE13QYzunBV/rDhaNjdKit5xVYJ99Cwq14EwNs
zTlLcOzrox/qPhkCdUos0Chp1ew92A7NOUwMGcaGp6xcsX7HLp82bHch8VV6jGGNPAHC+oTV38bs
9lnK3uyJWZdJCbpIlXvBSeJ027bzYOBod8jGLYP2V77r6kkvh2hgv6m23eXLcyaid7T6g5tN/zUo
yusDtCtBaCmT6dLWAxMh257GWE7868CS6am2STI8beP1FmbfEDVMbOa3LTRaYuDWE6K5hL/oGkcg
Gpn+1EAEn6ORu6DFF3gqLf6ihTi8ihPTQ0YihRh4NVhJs8i2VDUvxV9ABl6e7TuDDOi6HyijKuMN
xKjFixruoZg0w0PyDhgbo5aSc8VlqC/9KG275TgD/CXCGNJpCkDs8XqOAHkoNJDKn7Kmoo1/IC2F
kWfuvJpFJOf+mNpb8yIk8LHJ7KCPg3OEl7ny0uf6VmAkwksgs/vYgeMGlqO95SAmig/THw02mPzP
LhMxZM2GQ3lLO898pgyW4Ivdt/xL0HqTFpQ7GTElp7HV/oWHIKsdqVHPpzieEBWqzBWJ0Y4zp/bb
+a5svNZIe4s/u06e6QBgfAVrbPPjkZycUaK8+H3h8BkD1ZXqk1xoG/Jp5Z3AehGMnr8WJwn6xqwI
F4t06clUF4GeirBL8fDGaF99YUI7OaTFSK1/GhwO9EHzD8bhnfZW9BHXJxVejg/0X8a9RUFvkSWT
vCYWaHzgxaSZUVcBKGXJ7Xs/7jDbWm5uTi8EqbAQn7DJ/Jtqz/dxy0jm9HgnFi6dm6Bnlrir5A2h
Tz9wsc314HTX9NFnjLQsIq8BqJdcAvlg0jYk9gxsM/TfFPPDJinr2nH5Y677ZZfuvE/5zb9+f8bh
nfq8upyDJJSS8kjnRqyNduNh7qzjjCD8PMp7Rf7uozhdCTQ/8B8jvtANwYcBqwQ9xg2n4mI464W9
W3zVjcmx7v1AUL+ZLLpBWD7J4wcFHLpGqPfI6SYVAc/V+oRsV+aQvsDHkm3XpqKoFsRvVt+mMFTi
9nzRxCX8NO2RNyYydnXhJBsMi7VPRGEOmWCCjHtiCh32c0k7466CDsFga4dOVH1rYSwkovCwFam9
gs/JBvpSDPZ+BJouV9EuJGbqruaxskf5lzOnhtYdJSoJcAvBGVRWoQknu/ctYTQbzHF8zuPHYi8z
u+yaRPXx4JtQFwUvRn2WzNZ7vmMuzNN6DqC+UFHtvhgnO/ASTRgztLr3oXOv7o9XSbeATc+0GLHe
IBZjNq7h40v90Kjf8T+9Yvl5NbgkdYFPOsIr0D64aNvnoakLfjGEysKQbi7ZhA3lmDlzWcAOcdzR
GajipV/FKkwHK9GADlzrUI3B7+0JZTKkn6Yj0+nLa99rGM5Q6dpwJgxd140VeUqKPTd+vkCLAs/A
1aLMqrwoAGXGZuRQakfd71d5pOb3bKM+OcClenkbWNtoFQdhug12J90jgZB9I1E9sLLdTx7RuVB8
PInKyFPX+9GvlRIUaPoDzXl4GUpXsKwAooCI2QyLxpg2E5kUw9vY92LSsjZO0+kUv5YJxOImPmbw
uFFpeO3Kkhy/poFSE3EjgLfJFwooVjgG5lInNdEg9Fu2H6s+lctN9C5/uyg5PDjSQcVdG9FBYPA3
56JlS+QzOgG8YReE/feR0mPCyEqED3NsWf+Nu8tnQDGWa2sA1Jvj9vo9IIsiYpCwjzoDEYl6+wt9
bcPvt5wwW3MF2Oe1mGAlSjW024v1W0+mPvMxB/G1gSM+BzJev/J43i3MuH0blVIQVvp0r3VjrP0R
G1cbAN85R3YqYlXmwP3f2irzrruPtGVN+P5rMJxsgdd33yCBUmK63kvEFYR6AO/4Jiw/LwHKPDiC
UeNlLA9uhw1BfHyId6ZuZ9jXVbiyP1U2ZZRSUCwgSeJmZkV4A9dldvCSWpPyUPrgsdqCfiAFi3r2
XanEVZ9NNveApXlEK5ZJBye7rW7FwnNpvqBRPfGEbmqrn47/4QTiXSYQTOVMnpLKPz9l3R7iR79G
5pMVSXblPbYFpGH8UREgF5qPpMLjOgmBYOv2BMjH6Jp0pMMJnCNbg7VGQ7Nhn9oz3IIGVfwg60ss
8fQ+Y1lmbrb/sBxzy6KUFE7clgylG02kL/8Fj5HL+nb3hxAVMrvjnvFi1ft+ZnbNhCy9Z04wdtrV
ICbnEIli6noNpgOulG46F18e0o+CEzAKxX8+6vCVwIj4IDOKEWfaK+turrcm+f8ZV1LOjnvhw/FQ
65qYy6GY399n2HfLCXdLonRHpF+a034Pxw+Ozlifmk6ZE2GVQ1RGz8IyOhFi4mNA/Mku1xIvUP//
+mJn+sIIh7IR8SVOKaFmWuyVNt2rNt8q9hREA6ijWFG6aRKOT3tzcoUuqKts7+jX7+sGTtxn/ltI
gX4gvpZijT8+xYxYNzTftz452m5r/TaFKTiYzGPK1Mo0VwsdSoSJvDuzkG2S8HJJmsToom/pOBpP
1bc4qWiYQ6N1RB97LygLCGnSYQhUtiNgehrC8D1jn2DDy3IVBmF4+u4QXIc72X9uEWIwj60TTXwa
Y8xhAoYUHoNyprlU0YunYdsaTh/QVsQebxxmh7H7G7VUspNuBTwKDmfdXqvjAj+i9b5jZcA5W+JT
d1D6vYoPTKKbxSOr7l1nAQQrBP+zFuhBILSWHJSR6hfO+bYKC8AM+Lsa3jXTABoG4TYhx9Ey/YQA
RQm87pOwCDk6xdnSdIf4XfjRkqfA3NAn/9va01XVk26tUn7uGaJgVgYrsLpGa6Pnpgo4SyxoJeDV
oNEQUIhIfj5AhWODZos9O8qQM3DCddqx7vwtIEQ/9z/Nuv6BbdrlTRg5hW+PoYgzL6kycCdUeqEU
3IuJ/UwpoKMttIjZknKXWb9V+xj0te9ySTTmcQkGR+P43xYYQ6Emc8jCg/RWzRnyJspUFR35biIe
fRgcOtvylS6jqkOBptQcYEBTcoCPCWRJh0eblgAlwBwK9X6OqbTFMjFJCSsabJFuYdfJ+AX7KJ64
NZ5BJTHDpsQE6L3K72+zb5H6MQ699btlO6aP+tAmuUeSpfYL5JShuzJOKPCrT4D/VfB7FY+3my9B
7oNK9Zy1GfdD1T0Q8T1s6HUT8Fq9wFvk3imB9Lln7XzlySNOdXl3mG7yn3I0MV4NC1eBoiQP4FEl
VKEgd9HbMZ89zLG9qQSIfkAjj9TIaSkzYJ0NoHwGZctZ+8QokPQuP/yqnNP9pD5jc7dMpeDfWh+f
F31fEc8jKz3/dBXs9WOFZM8rN25Uy1iIRwD6GoGi568jfvYSQ2NJAaePhaXtS0HVCSCOTLMTfajk
3eiFESKoM29c0d/KOnJQLWu8VTzlOyiULRYjWbkyPY5EweuONzl/D0Dwo+m1NDVr6wjVaE14G6Or
2aAXh0jKSL+TO5hriFxtklPIM56Km2RSCMp0QYmkGlWfLmSAhR220cuVXdjl1lMOCt+nZmVvmj3P
kOEAZCnxBi+qpS3N2mHoN4YuC/XPg8+20s80YOE4nQk22InrI5PGS707Z6eLo92v7s2OAUI67Jdq
DpiSaBBrmfff6cQhv1JQa2qDBj+c5v4PJuWSQysQbkd44ZPBv/+vYfEqBV9bq1xQ/mQla31PhbSO
Hw6m/40uf+lt3Xm2I9zjaVn1gnhPpsCOibOCQKk35YuinC27oXwhCa2gE6ZZJo9mCLGz+By3dYX1
mD5QeBkgB6HG9cRoPE0ugQHaeumyw1can1/Y6dNiGYxSdqCtTXjl493Vd54QRrRvrCLq07qplZfo
Bg4ivqzPpwtmx8Aup0kHe1ELYqkHYhzg/lP1EBaXfCVGoAPsczU4t1r7iVYy0iJdBTgvTxg6UdiK
fzki5fDLttzzF71+pYfD9erVXXamicPWevdlBlvN/01cDTLtC+pvnl8SEANON5Ag0/JpmdukACVw
b7fdWxnMLmlJx0Yrd2GK2IICuBh4SaHh/92sYMt6Eh+MB7/hzbkgotoz1+nWLolnoadydVy3WQDP
0cuKMM8KdSSD7xPtawuKyqNceU8Vtk71FtzzJatgE5cksUnQ4yXnLBKa7Hl/oQFlNa88dipqpgGs
K6YAK6a1wjEm12GjP/WfmTb1UPPcf4XEopBbwyQpMIe30n830McPsKMLfZYI+NktP7E1QmFX/oew
2wIkB13UKIvthRlAtH9ajduAhYMGL5AsVk/MQxB+54R2jflnFCMwihlZX7t3l5VzGtma4JoWdkhI
4hkFEnlJAuzswSMS1wp/HdWWd1lACzEPbmX0onMTXMg+recPePHyVnKVGAeAIJRWC+mdY6qbWzwZ
7fS7fEJE6pE20E7/XtI2R//NjqgDVz/ZR+1Y3/snc6GGnaOf7k3HHjVPrNfp9JvShQ/bPsQb1YxL
4GnQDCgPzTmu8c1fqpNUhBdyhn9wLxgnNqmrwGtktpLwXJUObBNdLZQJJH2fud+9Jnz4KoWZXL9+
Tm9LG2qy0/EamBfoANNhE/P50fURqTiyyBXEojVi/DxjAcaIHMZPgFp7AmKd8UGf9eA0z38GC8Qj
oD3y6IGORt9B33F/5JaeekDmYCY/lipFR+fYbpExntfxGAgdxT+Vhho9vJg4YMhjKS3IyQ2NApw6
ynLomChFsZ08nu1Dq1uIZGGxDc9EDZUT+EcVfiOrtA5Jk2JptuVtzs27DAdis0YEmK6lcQ9R1AhW
3Bfg0zQcl85fR9DEQpfJ3JY/EyY/6+x4NIJ+xcVKu6A1pEsbo7CAlunY9nBi39nuaY2YVBugpRQZ
3mfDecF6SKEa41CRGeWvXsNoWJD3MKdc31aXr0G6Guo+FMySKIEdlGAs5rWr0Mh9DqbHNeFsLyCn
qJKAnewZcDCVfOFDBvs4wlVwpb6JY8judN/9ZgGRGzVK+WIw8c4qxfsEt5Fx6pARwNJ3J9wHUdcw
+6VgBuOMXIx/kq3d1EsFxhT3LSDVDOomuolZwmGllA7xUH+6O5cjXROreXVNO88kljGu8gct7FHk
JropW5ShSoa5xQ33PTpl92lgjqZrIxZNWc8ojUtdi4Go69eWt1j7tblb78mB5vRSH/XA3Jug9/Ve
0gPiW7CLGtv4Zt3YDauBud8xbyGKsAER3k2DfI0fA0BtN6WeMOlep1qrJMPZOcE8g6GEAaHGGhPh
iPOk0JcLQWb5x3o2xcMrCyKf2e/HbxmElQuCuXmIjgfcmZnqlb3IEsz2p+qD5+oagMc0wUUklHPq
GMo+/gkLg3sBmrd8heg4pCfjHLXz7L+HtbyzqJFo0Z/C6aFlZR3+EVn+30pYT8v5OLhxHAKieb6z
SMjT5FIdMGpKSs9qtbnr6Gjkdve9+AE8qwyKI/eHKEDQ7MKb39+kELRuWKXDpXeTezxi4oa5jFrv
ycaoTZKoCLxZQNAIpr/tRC/c8UJjZVQ0IU/fzINNQQ+BMEJS+f5qr4Va7kS5eRPDl6MZna9ABAy2
JQTjKNYkSK3r2PJuQuOGAgLVXyGApDU+LU8/asjSdn4Kyeq5DuA3s5ZWFE5aVhjvvndcAOJ0jP+r
GyIKoPvC9GCXtE54buIy6P+C+KvGoetvxeACymSrRmk7sr1nSBbln+r/OE/Yytcf0APDLqWXWB0A
G5JUollXNV33uEfzgrzLxr7DfRqER/2XPHvA4VA06+j1ZQ48zuZu1mH2HvaMEjRQ/omfLif99c43
r8Ht7EVFSukI4LVpDfpr1WBsOw72rlnbVO73mwoSqaL3Ziw5nLrZn9ggVCK2eMq41rb+Y0fr5xWr
YKjeWrW/a288JXeGdlt8sr6BbajcfWzkP7OEjxu6kMZQd84e3oKjPwzYN7biBung0kk/vcoQTMJF
UJNzD6L5hFQCSuqzKMUlUNNUTBHvxuof7MFjBWAqmra1BasuidrRjB0F24DR7hKaoYkRjPnUBrqK
dERxqpXRyADK22Jnd9gOir5MNJw8WO5UQwbHZTsqw7B3EEg7xL0jqMjQ/LA48AWXDt457P7QCIu5
bAyGlPn6Mj18T/gZvDum2LKBNp2a2HcXIIrIafz2f8BvzofKpYXe2pPiRNPw+3fL49siOmMxoxea
SOtSJwH6pAc0c+IxK+KqiI5pU9eVG5UvXXa00qEQV1F3W29cWvIEjSMpY3BKcMyw8uuoGiMXxaNO
cdXPyFQtoPB9sfEIXcxlGW9rpKenfaTfYSorozM+DrKcb6rjmT14WtfKb/KwbyxQtJCPQpx9jH5r
jrHV9OQLMc8JJsXyBs694B50kBFEoW4aaRJy+ZKgwmr2bWVoMitRtUUYWbQpbPNNkry/Z6BbaCQ4
fIi3jxXkrb0G0JiCcdpLsddT3SabxCqI+nPDZDNJYdRFiZ0uomPwZC+UM1O3uZmx8E1wxGpfKguL
sjCm7q6b2R/BY/wlRPHkadf5rI+a+GRfSdn7gBc5RPr2Qr71dz14mj7aJA2w+0FAYxB5n1+//wk4
q23Me+cT3u+YbcRIbEwzOYakRf1jFahlC/tSjDxYA6JDgfnqsu1sWWUcymAqNQ8ej30AGRjAbTM1
Hn+gxW5NMWekp0uO7ABcDWx9ltCny1bqqsChDuevBB7GjF3/2gz/hzncXU373iebfLlFI6rB5Tvd
vEfFW1BQO7PkZltoEusms9t0t8Jw1OVQb0stgtqZHj6f10nRda3AvUroHGx8jZb/L0wmyYrIhPcV
MRESo69gv5ky51eHvPDD/rNoS112E5ycC7YU0RBWWhnyty/abn7Lqk6Ns9g2i9wf/DsDDyWAq1ZO
oUJEh7CKHXJruojzZELzjsfEE28r5PCoiyRCCvqGf5U81jo6Yvv/O3xMJMbTxX1Mu5mL9HZ6ojeF
I6hwADjPCXq6wHD5RhQvWhlgPVBtH08plrX0bGRcwcAoYDZt/sAvqXpM0gdFC6X0xkiKUaSy8nnQ
/1aj4da9I8SDA/zLw23NXB2Qglg0eI3wY7KhsZL8zUsllYzxpUiSQZri4RXvOmNVK5BgTBx3Zgu6
av8jjp92NfJ2sebUcGG+MTuCKjXkh3lx3UfCm2QZ+j/AhL4s4qC5mpLWP61bjRwpHksJq11VMfsj
UMBlOGlewDU8bloH4eZXdl9j085cqueo2skoWD/1WrZeUMCJgx/B2ioaEqvCEBgq02Mi+G6rwuVe
Hr6A2E+DDT+fsyuvHIMcZbNnI4DsuhRxjprCVo6HrX4vxHDQWBe0+XxZB9wU6HFoxr201XNuAfsH
zIskaebWqf1R28LVHXuY5BW+65kwEoEr6AuSZrc1GHIwlyeZIY5I6tX5M9xchNmosya+TwvagUKX
+iA9qf68lhjQ0sOr+RW3VFFguVXHba9vwN3cdniN0BOoxQifQBkeHNHRNZ9hqcr1Xo408NSq3l71
kNMpDBc6GVwRjzJflKg1KGAzMqbpastK+EnOgVMWrGxvq7Y0TcXl4pfeik7VgjQgEI3XGKRS3Lzg
RQlD8iu40Gm+TGJHo4xeCETAYooaNS9YSfvom0dG/su3+NBvUsU3DlXLULuzzP3TqZi41ykgGmzH
WoDIxDzK/U3NL00mWbG+ULk9K4O4gDVTo50kRqNk3xHvKZzcXy4zo80sRVZTJCBCSGXI8jRqKGAO
aaV6HI+LgRH7QkcGtWZAJbIWTpE/nUVOXLvnGXBE40iHSpALgXfs6HTdYFEXOsw7Ht9J3st8GY2X
KKSDyeJCcWXNqx2sah/AaAzii2sksmPMvvUNjUEk7h4Fjg5l7CtE2sLu0eNo4s2zysANnNDoI9zX
eGMcvDnooqkQEvyZjVEOTLnlxTdH3y8YuoE8upWTP6MbVvd4t8CbU9QB+qPK5rr4/R/iOgOG/0uS
0rVESxmJnRi/zDEOW3P0tRoFzzOwJixY/XGD8wRNlx4p4c3iF8c24cYalPN233A3FwbbtlZHHKcz
Rc5rAjXazChVkvevlC3aV1VmymdxDFeykYw4qEVKgYJEnaeDZqAN9GHhfWmohu1nzHB0mI46vHto
LS8WA5TAKKLqsj8oUyjErBqLaCh2V6L3Dq347So+aVudoTMqJY9ilXRrYFJHH8FcwWPtJxIDg7rN
yA2RW9OHVxG7N6heP2Vt0ToeNw42/yenO3HYEFeQfYuj4Fl/d5+OMvZzr52jwHm0Pe4H6AWAYBbK
e58Wpccp4iBZ2dO6ER6qHM3/8a8uyjKXjjv9KROBXkeppznlnISJruSI2oi3cIHBvjvuXSixM/Lf
O9arkhyylotXeBnVz0tUbQhafZ2QcltaVZocqe7AqJKjm/s933i5UUC9xgqXgFXL7LWUXWMBITHK
ETojNCuopqFQqHVpWUh19JPVsJdEjb5NmDnl8t2WBWfY9lJBf36cKCtitxpYt2oaAp73MEm1qs5F
rYRCRXI7rLXVNaiNMawFCT4cLCanavDpZ2Z86hwLczrfipwOu/xxBkvh6qv5aoaahnW+KY8npqq2
+Sa+JqCFx5xcrCQO4p2MKSsH0cZDCNa1zWCZXprglH3q1pnmcArTPiOp59IinJBynJ2a7JTTnNOP
j4eTbV/1O+KMC6KoWgVJZ6pGBjEo/iL/hVvenVxWBTaXvLGcxeDgpDaSFjq86uEmL0OX4wXKgQVE
LlYfh5c4sH2S4dyhma+1HSHyxIMd8kgLhsY5MjLxJL4XBE9BUK9mulnLopE225A2YUp8iieAIAIz
i/GmPeSjMHpxJ7Pumv4bDp1+isOWVu2GTVRUoCloTIo9Tpcqx2t+Oemxu4QgdEIZlYs2m5cH7exF
8sifC7SDPuuSHrCaEZUCQuSKHNvhlpoTECvt07P2rRQBV4/eoK81sRPq0uFltU3ikrI3YSoSCR4R
3UZxJkidImhiAJQvteFmO/vrJmPu52K+NF/o6BJmJYa8caEWpBY02+rvS5pGdVophRSSyQPV7Bwe
MWxfLMmBWqvFmDHEFlf4COfmV8wUq4w3VckE9HKjJhx4U3v4xfE50SudqEgRmHp8X0yoDS9PIrVz
tq8d7ZjcrmoIQhFhU7LAQaK4DEk8fLaWVcSRhxk2o/QdCf1XqCooVq1Jz5UXbQhD4mBCzYFPNRyN
QfZfdcqXTyI46JJjV6X2DRHpKx1s3rixwoSW6j/neU7nxQHu2R+eiE3zHv4Odw+EWuPWCsW7P3Xs
XfsTghFQFXINhRfJY2L6Iu/5ZhnibMMTwUomHj6iQS9MpRmBxlL7SpEW1j77/KpfZoKH4xQefb5F
jQGeLcXdLCvscpBlNchJStl6FxAO0gT/hJCW2Sm6+MNZEpjX4Dwu6ZJaWJsS+8dEtzrxvSg4FF5o
t08XotZS9jzoS2RIa3XN+NAqEvbnKmsucq4It8VZxzm9AIRcv+V4hjbgOwpdssmvzyRekANPwIkV
RVCDBKuM2UINrFlzFaZznm1WhOPYb+JZ2FhDUd0+iABYTaSYb7JS+1nDKAf7f72rctYwnTPUob0L
zwD3go15P/JisonMX73NdB4kBG9UqALTylEPIVLAY8eIeEsFh3EvkfMwkm553um3D8Mxaz5AgxAD
yPnSL8r4RD1kn4f7yFe61RD0yLNcQldnzwf7+pOVc4rZ2ev3Mm17Fb5FTquoUTFxeRZve2MUWPIU
QZexdOKQgFljK7EvfCHiEwe4jgBIATkZ4mO6VjbUBLumufWGfdqKg7wXZNVxXsD6zC11AceyOgqu
Xof4mjGDxUoBV5GjzqKfgIACx37GvJptpkX5prTNCjV/LVEuftMNLd5SoCzRI4ND+ld5+3WAamBZ
qmt9F4tq16+3U/E7HjG+QMI/DQ7eVMccn6IcsdEtcskjceSzlneK60xG+koceFEZIjUCJl1/0Uui
cO5keOnBvf24NXfzErv02eyvcPTTLAKGgvDQsmuPmYY7qqNlomMxqzTcWKwA1crP525eRx5oFDSk
dkbXad2sYmKV1wc/MK1/FsN+I14eOUJdxaS9drITpBhmSij9Hbv52/r5+Sqng/vmc2TgWdnH3yHG
lV7mXELx1s+cq8HWydJbWlVUjBirpRmvfFgeYDz6Lk3cmJ6bwCk7vUwEOx186diUdWsPIJevotNO
FClCyBZrMj2AUODVtHk5f05riEkK5GCEC2FYRg0pcTh+JfRH8mqM1A4U/ZvaLYIeUA5dMrEaym25
PuGc5B2DD5TJu2a8vmk/EB57G7hucXl+SrJtDnEPISwDhaQuFGGnIHL/wNOej1KOFQsNw3NzRVQQ
ZM0+bsCkbKzuLBaovgErejywtDMrlLyrwUPmDyjjS28KQ61LslplGmlijZlhpRoeJZbA/RBw8P5T
e0rb7XTgQErc1kSV/6wmZkiHz0U1e6apDrYoDbhdpw+CrwfUUNlFVeHsv2egCYnldK0J6ZRu1aLF
+q80amhWDxraHWEtGhWdLA210ml2k69aSnIIxdqeh3/ykyUCBXgSusjtRvAl1WovHKoAXfX9y27r
fJ2GuY968nXw6dSkU67LCqchhHw4fkrXXP4+e8rC9ydXaiUprT2f+OnoR7vqOWp5K2lmKTluvDWI
xryimlnXe0PbTGCcQJiukr38jqoa8nnlVRweFRtclR8W6wi7HbHYQeD0F9cCrtgL7sfpwfuVpBS3
VOGchm5GsYhWHn8SstxTBHu1PEpQFNTrOqVoputD90kasli/pX9JoHiaeubJlHc9XpO4Iguz/Df0
EO7fxDFN8UbDpi31Qfmyke+107OgtFt5/8Ffj27d7lWGsHq4nrJ4Tv3R1av6fygZvG9MpvClKxtJ
uBFrTkmzkYpA+1W37dm5ndmaenkHXk9Ie0Gdd6V+6ut46PYk0wShbAKVh3rw/jhIFebtSlM0flrj
H90EFC8dhzpqsgBjxTtVCJn+iQJv0YBWbsc6MQAksGYyEIxhlFiJ2JLBfqBdfY3mV042vdVZvrbS
+zjsIa+DO67zMbzZdvEP8r9BVpB9NJ1Sm84drItce3Cq/V0cmaKIMwUXizBXvO1hrqLN1EHkrASw
l8iVBNK8bQTdfUWpFw31M7hHbIiddkFKqMGrjQuxjSmxMcyKDFgg8OukV5GdF2ELm/wPmBMsoAT8
PLk5TUD83uV1Idv9aLMT5pTpdt6IaW7BCzuWnuhilkQ7QY5BPqKA8RRfdvTJOILvPmYIWRpFGyjz
EIUNM/TCUgIpqsa7iBwtRzsNlrnoQ4Qk/eKe7XYWXCzSEHIz2epvXS7cH52ZTm8dEZ9vAKlKwQLb
AATbAigx/qxG8PL4+M/tavpqutO/WS5bh1A7IXPlQ/OcK/nRmKGI/3q5x9hMeOAevJNl5Jo9eoFS
2PSPxZiQkyn80l/Ahu+Va9ZLEp5F4gbgCsD67NrOfl/xoVWsugXEqTMPhKUyyNzkG6jcBkWPggZC
cJwzvRJWxxURfWn+cLQHQckFlQYcpFhMuIazd6Jg4IsgwDPy9OdYV6tt+LY+sUi2geix0lJuww4e
upu8RUv+FVWqyF06dqK1JHKbXX1f2EAnqLoxET6V3YRuEdqZesb9pL+ivTAOUCP49UtwBetirMho
5wpCUinxc0a4ORXdNJmdJH+G0sVovSiGgMMZjCg9uDIlQLLyjijMdoA978yR/0wjQafUVf++YgLJ
yhIEzqGdvgJSZ39QXZI3hcq+p+HzAKqipjb7ZcLHb+L9IqLNq5EvGyDqa55RExkvzU0d3whvlJPm
Yw71JleZoj+gLVXCqsH7/I82yqhKg7Wu4zUQs2oN2BHTO4SxmXRmFm1mMTU/T+lrwBRMko0QrweR
oGkeZbAI/72uH+Ly4UOtcQ7ni/fLWuwbfmwQgtqvDXaKpe/N80H1OGKq+2BzxKsfPxZaLYM4cfBd
qkZKrUeSNn9FbMPBwgOXcXX/4JbrNPfszuCfD3IAAokIpViHNetP4gRFOgTGH6U1+9k6XegdcD2L
ayliUUYSg5bKlZujQakEvvR/7HbHZNdv9bc3Dv5Y1ZsCiDoikYsjhopSoiYBG+2Ffwtlbcvo+VdN
cbKG4kzOR4R0FxPeNt3kSpjPIyStIpZLd+JnhTDV0ylE2bSUyf5CtU7H1ajAbCR/Y79hT2WBRBeT
1NFsNBkngAZhfXrzJW+zgTQsZr331pMEfxD1JvsCZ+/M9o4cgVIzyRM4lQQoKA+A8wvdKNr6jZ+s
TR3uA+NC5g23AvvQoxDoU5zSFqpYXXf8ZS6mXUW8F6gXYUATZCL2oElARUfoIuUXay3ZpbhQgv5C
SdlRIAA3ioUMMEav5d+Ip8oV1wQZvCLX1LoX7aak3eRdOnNTj9mHVQLfRXiy9fXMgUQDAZQ5nlmT
+5ECm+uo6hh7CTIQ79HRM7JtOiPF0vhp0XhWqd4EW4dYpbeD/12gItE5b3+6AoxdT4wUvaDj0NCX
+RsNVI8+3aJulSasRYP1jOrKznlI01gu17RYZWNvxIcbBFVqhypNDjy7tUvJ7uHGvOQqu+XTMIh3
8gpiK467ylKi67FLy7ZGghpGmYd9dkM2vI3n9JqLZLFybQohyEz9mSqDJJEelY+HYy7AiIRpI8eB
FUxXBwj+L0Q9DKFxmE4tBmx1cwYaa05Plj8IDuwtBTViBAFb1kZTnMxPzbB8UKSvdGqCmHgivmaF
NlxW+e8ATulSZJOAIB1X1MR9SR2JLJL1eXqxamBnrOU748ctD34CYcS2EkjcC1DP4e2KcTS6O+Uy
NQkhfjJ33gSIfypPhvoMhbIF+r3wQs6Fc6+WXk1YoJ6y0G0BtvybsGZ+bwzx1J5MdhHXbfflhTGb
mpAls2NgKPShwa8625piR3trQQ7632sqEnUdwLZ9bBqVj+ReRgwoCo/4sCx2mWkgqdIHN6Eq1QxI
i4b4+fyT1LMBherTLNq3/3oBNhwxdvpBR7XJ3yDgy3ELUhGM6QyHEyhNJXteeOulXC7DoSEgIoHc
ZJlDq8vk17aeV9aQhdtAGEU2VAnYgJ+dT+sYoDjgL5f/rrmDQ3owZa/X+LpEq2Vx4Xi1hTExQPxm
6TTaBNUbVmtSgkUxmuGuK+rmlYlMK2/KwFb+60D9VMJlFPZMuCjhhP+cWrGv2tIMSfq/gLTIYK1F
DXS+bJ1REdpbnVVgIv7pfPq4M0xsvemgO08sE7AbMMev/r/aAsyJbBgta5ivSODo06Nl6ajhkhO9
4S4KMTme4Hv7wty7LGjVguhv2r9EYsEbLNHKffnP5XrkjAH/a49WZLub0+tVmyQC1sDFVXYoOq6+
iC41+4kAUcLmENIvJaM6NHL2pPN7+y/0ToQhxkVIDORX9QewXgqClTlHueDU4ayGkeG5hxyEjCvY
zpBrVy5p/KJJciA/EpkRWZOjXK8ofd09r8SdTJ41i0E+U0LzcOLT9sHJiZ/2SLcHbAmSyMN79XIr
ns6M9rEouS2J1Ep3dwHtXMJTKHrtNhPB3TTestGvXSzOhb5QbRuGqZtfDtUKyX0vWbdaIs4h8rPc
cveZ7BUrG7hZFE6U8HoKdV9jNJ7WBhxEEEuCe4AnHS/mJKNZX97sRQtRttnFCxpPgDJ9dO3krkq9
fYKOmZmyhqIgST8vaHI3ZZsfymG82ts7I/mirzsfKP4b3wBPAirIZKwcJPpngtQ5lEWUcwl+Igvf
xNCDWEAotkjpe63uYoT8yuAsJt+His3HO9j2+7CYr1zK4GFe5V7e99aTFLOCKOmW9yaKsto3p6bA
bxygMjtzSKbQE4gJSQAoJHupuDZk0eGw7zJrqmRoW2o7DlfwXmEYz2Rx9iHFiwryeIaTzdUa4Txu
Ry8SDXdt7lE7/CR5jiC5Ku3PtrZQ9nVOLlbvqXB7AYLoj/N5T7eEmUQH/mlgEU5MT2oLIjzCJiMj
IhdqS/25/Cu3XnM18VzTAP24ojTBQFw9xMoMd36t6TOckTevCX3ZKiAkzLfLjOSfS1JKVc3oloOT
CwC5OZVBXpI4qHMWdNaqwAdDzykR2pBmsW31PY4MIl+HP0284q/+pBIvrDwsU/Ta1gj73DqyZb4Z
4QBumdrWFVJpmOEwMIU8iVeiSWNlD0FA27SeAR3czOV8j5Jl+kcamj6n79c5WT/q9MyYEWuGLPgo
LQBNJgBo7yAt+feuForMO7DiXyxoMGRJxm2BbAPtTrUZ8eSIJuextr1mlmYtc6Ian6Nh0zoRb8GU
A49Amy+T/4oqy7kNlWbK5Cm9RVuYh4W07r7pmR8KYGgB6XOYoQzyrbE4cW2t9Sxz/27iCsxhTSiH
S0LInS1/We/6y/ObcVuSL/ooBeUInP5nyaGMivfLiIRPQkrvv8aCUl1Rz6LWMpdmdyJU90e+gaRb
3wBxS3Fsl3sl/Vcma/uLxbSjmk5JoEJp+jjR6uOCJpcwcu7gUr++OgRZzCr9mmTVirezCP9ruaIW
6bqwTpfPKAN1Z11OGs5IBszi3XY8QeVefRCwnZ1hpCnCVK6KtHvjk2XImvFzOhDRMjeBi8ifLxfW
MQ66LIcgz2l4EAYTVxpPfn3qPLfsglGv8csXCslLdqx5unc/39L5iHGMhLOgisgwJ8I7UK2fiNcl
900EBJMXEy1wk7KLtvqIlhwZ0/po0am69YMdgq/ptFbhrPCTpYqCpmmP1H+fd5eHfvftYDkti8mN
s9acVAghF3d8BbjvwKEQnEs1/6IttZSnACnvLl7TWHjo2H4wYFNp6i39u/qZWJpTuAk0PuzrRUGr
5LbKoMRkeb8trpmAqGNg4SdGHvXxMuVxdB4gBy+fqbtOIV83IRJytFa/KLaY3/Bbn0wo9onqddqx
eBx0kdFrt42QcenCKdKbyCFPIXhiABzqGlxzICydbHo4NPTT4pyRe3Xm6qWgTBThH5vQvqIKe8jy
3PmZiEN6SAFoYUdbRrfj4i6zJQURYGaxgMqh0FDCcRJG2FeT71x8MDh63yfiDVHtbvLS35EmEUxI
l2SnA2SnBcNSNu77alIjrfuNTTJEc/tagVVrNFJOQ8HzU+khvdisqTDnDk3pd0pKY4JSzKOjpovG
7KUP5+idBsD4Ax0xRDycsn77NN/gDnwvwS+Wy798mBCbQKK3Ubqg4y+MvyspilFEKbyhcT0vHscS
cZ4ICGfKKWWp38fKoGOgS08BGV5DgIgDBlKQ4EgcFvSlEEVTP8FFmatNF3mN7iLqsJVsMPyNyrX2
t2xdkb4K75J3PVcLP2xhOevjWLN6a41JLY9kx8OimyCpWQ32oxiytaqoUbTz48Hroo8UbKsLoXtC
Yd8t2v0RTjmwOVdRuwuvAAN3w7x7X2gaamJL/d2zLY17kbwrXtDf/gs3gZuRLBOO3RIa8YbdEgfo
QCTqPzlKj5pzBnUKmtFdLvfgyeFYyE1Jr6K1nKKQkL/zghggCJ6yaqI7q3m2vj8a4UKrUhA9bcPe
Da9g75AMR1WQ72zBROl9ljBrjlhY+4zC6kpbgyrrfxc0cdC8+vdJbWIu2lGNhAGsLSDPQopjueUE
ozYYodIc48Q3fS0cz2Lfz/0aH1KYmpsN8t6bnOe7OzY2XJwTA8JAqCuf2VF3zTkHjiuzCUjyVgxI
ZdpSnSkl02a5pLTgkojxJSOeUysYcsV6/7sWvzXVMw4UvyU30DUhnLlA6anLGuFKuOaosYGIYfhI
tK2DxqgQ2PCaFMEoJqFZC6Ij7j+9XsWjf0q3gHT/YTRGMm8E6flp5Azx3Yg6PFb0b/75ja5RT8On
LCfrEOgz7EMyte7hh1PJ54+BKkfjGgpTWtKgfxpYZUCmnWNAex/rx3V3USwD7oxDMIDFPGK+sgWb
nvTF9/2GbEZauwy01N93DGtbzJx/UtmJu2AUhcMHjrr3mihhazxymNYBd/DsbBHrpY6i6vqEPoD0
LDQGGCTHW+EAkTU304DxY94/WEe/usTR0mlLGylgoHdFXvoQHycU7d1j6VsWe5bj3fwGsg7+6YmA
RXu/Uml3r2ULS5nIJYYucWsFpn3yVgomzLB7hy1SXpxg9VTjicBk1wK2IeJkZ79KRLqWTo91UZwr
mBLQLMIIDDY7L1fOqXMKdzE3XfXYGNbVHJHc2Sjc/fwPOZjLeSUwgcAGWs9rVVe6ZSCuCkXgV19E
51I9eDGSjGHfubuCJW+kT+YheS+DnaRKDARkkuHXhvUqg8DprUhtP23NqgV1WFVcvdjZlU7w0Adg
ZRl25vJsAD4l5TvQDqGyBTNkUVo9kTBb+4AMcIlyIYG/e90hCjjG/xXDB/b4cnWgcKFNiB2dTIUO
vig4+/3qreItpb4gsLLktPG6HPdB+4EjgUMSDcZcNXq8I/tcrNLBNqYTb/N0XVh+ImCWDCaixQPr
YnxOhc4g1nd0Yb34jmG3wcCLFVOBOHbjw5w5r1L7QSEkv77kGp7hVip/lVsFtbU+z9WhXPbDw1DE
xZDi7G9Jy8nfWJxENCtUe7cW+gWWGvVydWUBQTPmIfTzu3e6KRtwI6Iydnp+FVkAnnQXgcQn45sQ
CXeFpbr+FBIGLDK6fpx9aNMTBXYLddvUzrGpePyNoBq8Vcp8sg4GibUjvJYsvavfm+q/0iWAgxEx
n3q5E+6OQgDafjQjrr1OgthGo2dDovyT4rOGgvRMWbCXpx0q//le8ckfHjpgt9m5w7fwJHQ7eopF
q1Ml4Y9rnQA0O7scrZgZW3qwCHRjIzrZl0i9qcVMXetk+50YVil5OAmulRAn86qAyU8y3tszI6G6
cykqEPGJu01uVCBoFO4LH6bMZnxZtqWxTH2QLF5ognrwtGm5l/+vCyFGdc9dnLycqIVD66cfFx57
0PHt5u2OYmgvQby9MeZtfzlpe0PodUKusMXhtsv1By8/r2Yt/nBKZb4rVQetFdvG+Z/hi8ugvk/u
3rUajaYodxKM/M0meh7vqQrkD6Vc+xHrMts13qs/1S5wi1AYBIwDqX5oH6ZW99UI9CPPTKBcrIVq
ievdeKJZzaTmBQGi+U4O7NphtsTT37KZw4bFCo15KlEMpjLaIwtpyVnDz/p0nVRTFBDH4nMzx+4j
d/D9uROUVoOZBCWghfKUKupfzaLAAtz5G9jycAuc/uw/S6JwxBRTPjJZFUXFR4s6/m+o8QwqR3FE
+LOuRVLU6jbZwMlOOGB9i4Qu9YU0oYnYMODTK9uZEjM8yrzeCsq6AqvOzjfzHuQjSXFxDD7Fp0Jx
55LWxPQ8Sbh24HA5cPGEC73AHXxcBOP0+G/S0E/Z5ABB2V56Z/30RLzR2LluvnB83c5N6K3Ze4Al
IMVC4MjqUyZDEhGCqpudTGLfcFJwUUIl0Z+pcPx0nqU9nqfkD5r78En7a0Ku6/lti4zBkYSE6zvk
/MDlhX1HZ2y0Vu7dTCJewyszsgSfK7Zo20co7+uC6rYtPWHnBeApnwItXDE9ceb/rhjqMBJa30Jb
ZdlP2H2wVz4+ltBfCQPnvpF0KsPVZdx1+3Gp69l1wb+eMeekhZD9TNlBEgy/+FvoUdn4YsFMlKEt
VsLBe6Gf4fdZcj+djz4nL+l6j2pPK3vRtO6j5IPCnsPpkMdwV31EvWruhOfotyUUkk2aVy2EoMS9
IbIU2Tt2xWlfa6SVvtvvN+8qpwNOs1pSltppZ1NL2GqcWM+ZCn6qCLZ8s0gPuF2S2AQHmdWOA1po
oGfv5ewzoCj+nyQChlhK0NkixEijEfhLytWFB3WfYc8HMObDviDjmoHE5q1Oh8Quya1dVY8MpHvh
ncrXLzToizZogwhNhgi8dv3lgCr/rZc3hH6snWyNrOubhC3GJvQobTNNdA4v88AeShvG99Z/PCaS
Fi56WokcGaMJDFXiqNrYtD2xno0Iz2hINjQoQpBpWRcR5UycrEH2l2YGZ/gX7RUK6PP+QhCTfq5Z
ivT5D3Fi89beU04GXq089pauLhc/kEEqSCjzuP8g+SdpXGjNEbuAmaN2BjzSU7A0OccdzfzRZg3l
F8UaLVBSHFNlGtBOK2XSE0ffEsC7G8gIufrhOOdboVpThzp6crJ17lnAE9PhWHJTHZGHtqkKgRRm
y3CzQp+QTZxSnwbLxnLRXyPWHQfx1iQLoOwijC/3Cxs3lus3YJC0Lo8AievfAuPi1OCk7flKQ+TW
ve5xTQpzULVWAsvlJ2KRBs1s4mo7Tu0+32u+z4E9/K1KiFOMlJ92j1NkHFHSOfQtQOuM1zGWWEGx
moGwICZKUJEedFxAnTHiVaTcuvWbEgv0IYmvKGyFP7A9+NWhBl+j4zLN9nD1i2ojJaCll038+kGL
TYIBz9lKy8u70HIgLt9SsXuFt99iLt5Gehp1HHP3bDBd5/ptit7NipN8B5uQs0aQKYKLBLp7519o
NLxCEJCW9aoPFRvX5tg1hAoB+5U5CH8da4OmG8uQOoKGVCKkkCLwylbmeMH17pUXTL9R9Upn8Y9m
pwhVeDCI753vw1DdapFoTo+14CnbetZrHYdFDd7OX/6GmUbp+f9tySgLgFyFdHE0LjAjCaK7yqKW
MQCsvacoWLNy2nuAYLkBVker8cxaZ+e7dk9SnVjC/YXcGzC1W4RluHpd5rEUoBiKBf/Ceo9+Wvzz
A3smwJkGtphEC863Iubp9tAFDFpYFxski1TUeUrWhCSMPM7ZltARTS0CyXcc///D3vhCJwoyJ2YN
F60C+hCuGXOQjDs6RfbgcEs+7yzyduoRKYaDsYhcfxS+RkfilR4/f+3nfy7HXtsJGKitumyuLHth
RhPrj7yHgiyZAaGk7vM9baZrCdLCAa2vi7DvTsAzI/Rb03iB6I1a1czUTYjJi1CqquDTWS7d91mm
of6b8SxOYNJhgHa54qgRNosJLVF3VPHTu55HsPOiGbGkERo7pPXKIq4XkTZkapvJ5fZwJKL9NZMF
1vHwvfhZMDmtafrl7+QUDQbJY0ZLyVXX0gCOCsaW1kVBV8Wk+khKvZ82x64p07R1/F49/LGnC3nA
5bxO6wibStBVrY6qB4RAV5p/Ic8aSmioem/vsIy+Ncrgww2hHQ7jx7RdcUM6/l0fbxR57swBi7oA
6gtTjorPFxs/GO+zY+w1WJWHV+6sZX8Tgu+574fLQGzKDtcFRCU42diNAjvuudtZgi9WrVfi9sVM
oOXtHX7Mcki1wHFjDKr3GN1n5Dc4MCXLr+I8c2StxDIHDi1JiGhIE3oTFBFFAhLSlJy8Uyz4wQrq
p4gpkOokuvr0muIufMI7u/9PqD58HuCxYUwPgA1Kgx/EDlQmv6a6S+FbaVtBrLP8tAEsuYjDMoyq
fPA6QlhdMAnmzNGaMraXnQ22CLgvglzgvMuPtCXnfH44qSUc8G4YUCuz5oKxF2HgK8wIw3CXATSJ
XQ5b8N9qxeEjVMV9O2US/IwOlXm41HvRZ0fbJMJgzwQVfJ6c81UByVXDdQmt+iDq2Pbfy/WU3CMB
tYr+JbwMnGF9ANmGqI6w5u0fwAgxZ+Wr84zo+EORCtJq2kV9ZLqPJD8vlXAd2QEJgEasFTHSMoiv
Za9R98eMGAVv5MB36m5ycvhlTPKsQokoyeYacMz4W6H1Tf8ZRqjyi1aWNI1ec2lHV4wAOKKKQK/I
9+tebx3lLlROsmtWpkBO/X6TGWEJJZ5DKsjvHuFAqxjKEPRt9MAjllabWXHWfUKvuF863qA2TpNG
sMRhudr3ODi2A3YaWgvQreJEAjo/W1SmhmckJj/XV34b4rtZdHkwy5F8vbhbh5PMcskpy0YTIlok
E8UoPC7fPQtTuFsBYUmLiUutYuxUGxKjAVmQI3FtezuyF8neAVgTfwC2MLOv1lXVOyiB4LxascRe
P742pGcV7qJv/X8pZ5zfUERwGfPFjaLnXdeUGtfBritgHksK+aqf5c+j88m5W2lfV/HG3jDQOI1m
xsYp6ZR6BxdkoKobZCCd6GF27ZR12UrzdFFuQjOUb30+680KdYMCN24Ti9qZ2OjC9BDGmR9rjv39
sZULZnM2Oi3golVjFcgqX60/Fc1Rze2VgjgPXIWAikp6N2CdMTb5a3k35lE9Z9xWOV/jCR/pkMfe
t/w72jDhAB4N1lcT6SH9uqaKD8O/vhGdBhejkTNSVJfQ02FIvjRBw/iuRUKTSyFC3TXNMWXPs2fO
+WDKCewJkO8nbYre28mcpyg67lVsuYsTgWMy1G/PxvZ8GvD4NcVBNfQS2rb5yWqxVU6qzw8OuDfB
k0u8qPvI8OufQe7Aef70I5DWtgz/MdGSCrj9XlpWsrjON6NiyJZ3o5/HFNec8VqEypPFkE2KiB//
sm3wZZKmFXSHCFAbTO1sMDa+uz+fopRPLVbBspa7L4QAuj9vb++FbwK5MKqdFxtH6AYIAT2wRBCn
v3FR76L/mkZijApx9jb8YSnXJsYWCpTRz5vFZV++GDB/AWL7JoXIFHDYb1gO0tCRKFtHbNWB1Inn
NoyuaxWXqXvO+ASmvtD2Y8qy+dEMf0RxACKpb3D0IC1g3Z3Y+ocCEtWIZGwJkDX2Psh/LXzqkO4A
e4tvrpiNnB+y872UhE+f5CCuPqoOUenLDVgeZBGYLKqY3bBLWRSxD5hN9V1NvUfwzMiJwa2x0xZr
X2VQ+aa7FX0bvCnugI28O3kXsjQBTVOJtNJRMBWHDzVVwSlzYiKT37slmOU30uwuZZUIa5mJ+ZzS
khIugS6WyCQkeL9KnaymfcQun32y+kBqWovyYpqQcduvH8BIMCOkr9zywKO+FdgXhfbEqjodhjUL
oWIeDHdfGET6D56JjvydaHdF254o0Cp3PkCizYQUgDQT1UrY78iwknkZ6Sq9KBZ3D9iV31HMi5v1
d9PwpmYniu6QWgqs3uwy6QjpXl7eSsAfLJvG3na47eDLEb0DDmyEAyA55+U+2Jf77wQ8Roi6nSCb
ejyafPOa3irRMy+uBk+9MuB4jsSl37rDvaA1neUlhSQhBTC3wzSMOseRrEQ6ZyZo8g9zIEx2IK2s
uM1jw1Xv8QSc+4UUgbBayOP1GgYANsLlSAGDXQCwetxaJMEf/WWgKft3OnZLv5Sop05wfrUbHv9r
AUCctebfG2LoaujOCQnfA5vP+RqA07/m7z6PmBzP9dBGVJQZ+j6vkGy3uw5nfDvltmkEbFQPwjdG
zmCorTjW7DlicZEzdEazJMAA0SasTYulrSB12q+Z4RvMVkBoenKk7z2IARdql9YcbotCd6xqj4bD
7SpnYeoV1MtgJAeUrbSL5ErEx2ZJmsfhcIjXSmud7Fh4eoMjdDFWUv1E9zJKUiMg+v63LKROa0Wq
VTOkN8bAABY9+RmbiBXs8FbMVwOq+1LEh2XObrtnDM7ip/nNizQuQUniiNPNXD631ldl40fBkOWQ
gF/dFrGIaVsAiiGon1UpgccJhV9x52JWvu2iDHThaVwcIPNJZBLXjWLhR2rjz9J+id6uHEYuj67g
v8BbSptrC9mpOzesGdlXY58ZtVJbsa5EbpG1dzbxgjqgwhFWn9YJNSTKgG0+UPrlHYXBR/FtUvzF
TAERdeye0H52Be7O1LV+aDPfhnC5yyrUCBMVXkw/nqbGVF+vP/H9Lri6fyTArLwXWQ0b2YQveSsD
XYfPnjQyCMtWOy3upnn/IDaK8yYLBJaS3CPe1hwSM/kiSIsMjP57XCT3UTg5wq6jxBRumQiSfm12
G47F6N5ZPkm9lYWl8uZ4II/LXXFlnlCEmTMQsWKiJ2b1XCk4m8lo2EDnqSnFOWdOlju9HdCbZ8+6
S/EgNZJlDnrHsMXp4g0QUdGCXaIOd+/j79OqCaw/terUPziICY1JXZTJWWHmLaCjesy6Rbj3nOtJ
3YZP8MGHI9VktpKm6bXdlY1haJK8TPGXtwmL7dkvdFGq3qcQ7dLEzCoOs92si2ZX8CXzLDgoHv2R
YtCZcqqiyAtyOvCk5cgegpy4sAN/NkAPZRt9U5cwTtnkS03zNx7LDY0TNM8ZA9NK1IBC9qS21G/z
rEQdSznh0RGEieK4hBVIqIlbNdn6S2465QiwR1qA7p3XpIBQKLGj1LcATU+kzB67UseXSTChQYiW
eiUsW+ccVCwyroU/JsdDKI9AnLSNP3qVE1cApndaO8EGNqpzAcPk4d4L+L/rRghJiW0wUOwbswoK
9GRGqOJz6kO1bAuFzFpIHCxuOJOHlHTwtLIjaF7QiU6cFuSdbVG6soeKMEChqUxnrfQKtgKHlqlO
FehMTeRqMTDkKdplxbdq/fFIakn8/FezBFWY/hY8a3CHxNgwGG1CIbtm/xCiuSAVfo6t1ZJ8hbK4
dLD2cMP/M338uj+JZv1e2Qx8Tx7ziGozm3YdX0SIDBY3lkii9EMQ0nivxc3UkpL3wYNZZesc2UdD
muZS34AiQcJ+KbZjHAUoaf/neGomMPf9x957KxukbWGsRUc72h8xuXIqtcr9WYlz6e0OnD8wbtr8
JQcwLn2KPuOGj7gBQ6e/e6xXu24VZPkoFEF+rQ+A5Pd41N540CRLVn92WUW5UvoqX+4Y1SQ7cFfr
/JqBEjUb6SFX0kh1ToigLcASPRvdGXJjxAyGp056VVpFZdl81Jd+XFwkLtElIduVWljPXGSl+lXY
OKXxGSBTPWYqZ6pyH91920+bqbZTNmIOvtp3oiK1/R2LoPXcpmlX7lyaHeLjUCRuZ71y6307f5UG
IK1GesjL1xOJbSQZgDuTqfT2eopz+zBAh5UHIS6J+7FWcgc3IIlQZZkuAJn03yJjGG5u2SFWjA8H
9QfsbwB7F398Or8sCmZJ8ijHFAK52n4AWPrOD/zUU+t8BU1xrWyQiu5Jtq9LPcxD8IOgpCP7q7Kv
XRoLvhDYxv45hPWhyw1vCQzVtBSQJ9iWl8PTh4zMtv9p7LXDuP6DS7o6nffQz0eZPDjOIBtLUK+U
DHau+V62+qMn4cNAkE+mzvZe9q3ftcFRg8TOwz/I6iwP7m4PqZD5l4FFK7VY/SCPctu0htL2zcVL
AJnLWWGfVAoqKRDkA9H/HTGWsTpmm7nA1fqtLM3L4Q4H6i7AQmHIRHEoXCgougBA2ak0CgmbwBGD
FOBt9hQh6/e8wzerpihS9Jn/E4T2SBET/Smi7ni+wglGwM22OyDJsoGJBQVCK76lZGPu0wQdAgfM
8ET04Bkp0QkPvgTy6ehLvDg4bvEIswf54kNwr4Pwk8HpGalSJxDYcGi/7BV33d4cEkSwX6kCBHPd
ejVNz6eg31ONrPR7cNkGHNhop6YV6mRqQU4yyKSsqWVxF5HVN+tjfSt8L+zVCeDqBYH2Zqurr6wm
LnzBDNvK0+g5L3IUVOtFi3k8kMcrtj4fhE0xRu9r1hEH8wR4DS3kYe9vgkchPigXZ7qNojHR5eSJ
Tk1wgOXwTWDFmWGRiZb7QVUV+4mcWBVftXcpNZ5JCKcGD8gV2FrFt0Gx/iRyA/02hebiXfg2CZyp
8isSL0rKmy5ZobHUTMKtd8IV9bEZHAxHkZqeDjIlyeXX6JidCLRmXyHgUopNxLQNVS6HQP2mkTn1
Z7owugc09Na/cWj/x88bIBzpsA0b7UCcKTQLmwFacBPKhTIR48w5NZYpMDxVy8U/vuEkXm431O7D
UOCgPgOY+OvxjQTSR2rY7OB7wItqwcpG3ne4Bk14sB2gaBAo5FL+yaDRL6Brh7R+nR/v+4xHR5Qc
/2vTyiolIPG0R5XZSKFtv+DHMlfvGiBfohc0uEBnuwUi/xReQ+PUkTAMMqHAs8CBmH3rFNx7p9Bm
rwrjotxd9rvIb/7BWTEjo5E6/199ngUG6V3bf7ExcMsitHVDJqrJvhH9tVD6YZGqKDBwcZLvtZwB
bNIoTzVOVBSlcx2wHcTHuwzF8HKstyCzznTNmOx5inZKkVFbEb4VvlTrTie+ruM4cdKMGLbDb6rK
c8fpWmon++la9sxnEAUJDvzwHJlOe/kxvQzybIEQp2X+MxtsmWxFiFZz1KyfnAAr9SPhOAtyyDe1
RwgsvT6M18EcVolQVV5LyWraizXn5OqI69CFoKdjjzpew4ZUyDKGZBRaY8bs2BkOQ3QyRqNDjCWN
M8UoSplCFKl//A0uYoxQFvCFgH/rITfwQb05fDv05QM0t3J4yJUmZmv1qz6u8wmMpvz4cEMpwHCB
iJzezyLF+lzKt+LnaHIWiYQ/FzegeHaGG4uT10l+GGmjH1LNdKKj23DUmVoDCd/fgnbh7/pEPUYl
0ZMUzmCUcY9+HnYPHV/yUefX6zVpWN8pMoye7e2ewD6GdkB2Ye1G6PlXTTyhHIBEbnpwLgZq9yQm
ghnH1fwjxQqewXpQwEWAQ7GES6hzkHa3fdzSF33Ui5fPvXJj89RNlohl0VfTvfETYyXHUSHGGsof
drKbMBPR9HMGDH+28+IhAlthyWF6ky6f2eLtVp9VyNEQuMJyO2e6h2DNeYC6U8YC1RrhdcFugQDs
5n1YYV0wHWp6hSM1BpPUqDkwI9iX6gq/7JUVrVZ5N+upeG82TiYipACEwE5WqZy0PQQTkKJjt6RV
ksozFr9X7PslEb44GkXk+rxBfFvVTlFDTBaw201SinJlDsmmp30sKBn3hluGvw1lmI1nJen6q98G
9mPHNlqruArzJp/YvcSp118kELhuicniSX26vC4eFe6K36zF1cgu2hcxcnE8QPnHCt0S7xO9Jvuc
1RssKYi54DwaX/VQwiAPa28Mt87L5LvxVd6MiE95Fr3qBq5sK1MDbKp5UBecA7l2Pa+im3q0cuSK
IEYktkvSDck7NOv0SLTjnMvpdPztRgkqKF0zSra5OC6Nuz6zLGIPxb+mlh5WQ3DvO4tz/sWa72fu
CAiVGukFrOMgQLJcbMZJABZ26y/V+wPapAaeZufKDCq3dD/9Pgo+jNyL5JaNs8Nc/roKs6/yCKFh
4eQ3vlF0dVeBcsQxOfXuL0jzM+pC0tEDjE+HgnqXG92qEp58LcgJSjadI/3Kd3L34Pff1p/rIayw
jysHzMAJJqFKIekyer2lbhq4Nz0PrByyghXqKvs3IEC34lpWmdt1toj7R7C0fizY8FTCq9FU0Tmz
MylA18em6emXDZ0FHzm6HHUXHnIdNTadnrQ/23h6T/7ayB8cS1VB65mWRcKahV9LOGV402HCIq8O
58rQuKWsUIGiK/vEvOA0KD6xwjm5K9CFiebmEqv4FOo5f01wL1NMted893w6eyjlcAiqnnPER5UZ
uYw04BYLE81R5lzTCj0z4g90+dDkLRueiB1guzfdxB9LljwiZN/SDP4vaNH87E/VPFupkSI99yba
KQqc+l8Q54/DWHv8XmWVz8NMVvKnce7PlVArEgimpFKennlnFOmiAJim28ACxtQtSJEE48X2J3L5
FE844zNKlax6LQ86NvzjlyI808k5ND2FjsKpDbPndsn6wtYkoGoh9wsTWf76mAZGXGs9VTtAy7mt
cA18EhzGlugNdnLHOd1bUDwvq8MN7ISsNx2c2uLAv2joypeFbHmvuHc3I3Nd4vtpJGoZ3AexD0/K
irlKACeh8OkrDzY0SFA0AjQnqqukywEKKfB1XCVCGWiviLM+8QPLJfxUqpesHNrjNBy9pRdpKK7+
lqGPLTdhS05yrj0V8gduJh/WqfbiYxy1FutpIKqacz9vTsp4xQK5cwsGzd5K31VrrtzpfSaE3rlP
qUfJ0KA17AK7hBH+kRC5C7UOopK++Ex5axGKH9qg37bnV/E8hueHjMd1F3j3sIGn/aDZ4dfOgz0v
GlCN58pvv84wg97U0IDXjVQB7M1AIotCcUd/3vqlrCSAie8desBk9nKCT8pHallzuC2Eem+Hvpgx
xZLpLwlb47CfKSMYJEltlt6WVbt9a+V/ZOV8xBtIufui1/DxnkVNCeSUFh7oh4b/0mTznFNdmCS+
exGgDzth2p91CpxkORgczdSv5WgyjzS7imBwqteWMofHn5nli7vV/4etOrRXfEih5mnDnfR2o6iS
bH+7865VxQ+1vgbALM46LDi7psVE4KHzawxuZzCYBnp4CrwqmzhOFzryAVV8uUXVth6EOrAyAG1W
LPIoTiRosGQcGqYe4gfeIPsj3PRI1giGe13x8CV/+HXV2Fx1NjdBtMHK/PoTNlZVsdDCDhAkmvVJ
gRjxsEFAsqZXICRELq+QSCVtYLLLuhM+1jP7mGwt37mhzA5jEYa0dIIuKZzC8Pa01dUCk15Y8jSp
+hsW19PnK1Gz//Kmj/RKyqJxfTHOGbY4J8L26cv8luCP4racyuOW/G3NLvEzKMDYmPXX3LHhvDVS
fIDRb0jGnzK32S24yLy0R0B+81lQtAHA+9Ih2lMOBgd3B2ZCZrHo3xd2iPdWmdjRWwA52zRFQqf9
FRYJHMhPKyz+vWMZhLZK6AvkOBU5i3AayuZ5w6xXdmcBOG969jplAf5jtLh5PHMcQa1ElDUsDrzw
Q/M0WPfFxK1wkOcaSmEZJ2qJ75QyMmAAuvEwJp6AXeYpAacKhOluCX3nxZHAyZy+oyC6338GIjl+
QQ2nx0R7NAkPfXKCyiUTtM4WFZbVk7Kr/WWocQRne5r4d+SY2HGj51RfgTxsSWought7iNPsuFy4
ZHmxwEWkdOLrwNDH8qJCbiVUkKvCJWYoTDcMQuPy7ps0D+eq39P2RNh1Q13N/HoxQarPi8QD2i2N
4C214hEked4v30AHp9oNHKz0hw80g5c/nTHqgmGnKcIW4SmodnkfFlofcWKS1lQfBoaAaFtAELtO
Ll5TA2hFTAwqMScpOOkk2whrKCESFD3O3TW5aN46oU5soT7locPdgSnWO9UG+z9TNtC8LFvHsmv5
dZYIgB+7mCV3gnxrasXs4HpwCFuuHSObDEmwa7Oj3phFh4fe83r6gSFztZ3T07HiOu6rVMyJtqOO
KRbM6WGoKyFIhC+bD2gyCgFdCFOW6P2Js0q6Ona9dfl3X9o+pe7vkt6mdEm9PHx8c2UvbFbEC1Pa
98xu4ycmoqleNMea4o4buhcHV0jeU6TAzvcKbjAcjbfaE7M+iIxVYHEsfPyOLV1sQvGRpEQxLQZV
N0aDgGbFhgACEO64vfM6YsU6ghApXcrMe3grw7zbzoOV4EA/QP5cF9+rq7CLn7sM9hqJG2cJhaeJ
ynB5+CoAIanxG821X85idb1RQcXaTsFkqCggWDAFKbqEMj7IpdanBUYwtCt0ny0zUBWc8lCGkbOX
JcmbYHaQLXphajCw+tKnpPHqvx9VGfUTTuNUpDOGuYKvwnixFUHjoLsdmegaRxTfChB/y4V4J24o
er59pvwQ8WRz1dMUOPNaEM2hk8r+wWfrPR+hkjZC4vuXyrCLDWLioymkDvEATvS4Oak8kRnbzHu8
rNrqc3iBMsG2FHU6yy7qwVFrerBuZzWPEn5ZnhbQ+akpXbGcvNF3MwsjGAp3Pq/ezy5Ctt+L+bYw
mmjsxG2+g9qIwsBg/lQ19gVv5nt2Mex/g6sMVwW7EHZCGos30VtcjyWDL16yT8trEYV8M9Prp09e
9JfXdvhnx1ANLijLjadJSoGmFmcIfGBnmtABJKu0HS3Yx/v7tmNUAsVkw4AthZuVj1mpi47povNf
J5PSuuZCtI3imL37wFkrH8PlvbBsfU1Nnmg901drDGBfczUc73LlKjOLtgouAVRQPrYxQv+FJIMr
iCl+ATY6nUIwRsN+veDITKEzCTyjLc3/fKNCl//ywrRUZQuGf6firO0H4wdeE4oDALqbsPRLtcd7
17CM7qpZPIeYiEF9ieoLGi78osvft47gmkHnTU1rxGNEyChf/Sjp+dG4uUVd0EvJ0GkhlrAKQuwT
gQk3dJFqx4NvTGmEnACMr9BFD9HENQbUBH5eDAqcvIRUIQmDqE7LXgy3mApDzeOLIkEaMaFqeYi7
AkalwwrrcRl0jhv4Js90YgHw0YNMNVD+pGdpfDxBoy9POzP4FQqAvlBLfh8xUUXZBJUMZCAHb3Nj
4u9tnKgevmrGM2fLFol3W/8aavcDD7iMee9pgFuj/KvbCgcwX9FopkMIqG7/W+ovMebskytchj5m
O/0lqcG7Alzajxh56klLlRPP6KIhfbBXon6zOS9JPemxuyGjQ0qcxdzn70WnPiYlO+iEk7SeiXPT
5vmjTdnn5EdifScp+GFawI3bMBmlWtelhTwnVlUdZxdL7Xw2Jk9J0REA4cEK04VXW1C2KBQMmhC7
g0zFgkNGHB/pEyFn12/5XtOch/qACypZqMc6C3ArS7ZitIWYSqhklS5Rj0LyedTBkvKMsVaAboBV
AkQE1UP6cgVMRhD7afvjiIlr3aWNNlvCD+S6E/4WggON2p7N+PuVVytQ8guWjTU9ja/SGf0ar5ED
T5Ii+Ma8v8FpbK52m5leYpy48UQo0uNNptKXxj9nprvKa1Hj0HlnH/VUvvfq9RtSt3q9hqSstiOk
lwWbY76s4m5DTJQlWMpyAv5G4lafUtMqQmrsSn+nnBjI8eUBtyUY6qLDKOR5hIjHY9GalymGc6xA
wRLPr1KYK6qebPNQD7JtgRKP/UhYi/emNo2ZmAzL1CgT6lfFYmQVCfw45TJyUltcFo3weV1MQx43
NPgw5p0PEo2TugDApR0MkLTfETV9ICS3g+GfspMkm24UDdFx8TC4pdutz3KxLITTuxpnBCK3vZ9L
X+8BpFdWo7Mrcxo9JV3Grc/jfkJ44JHSU5aOy6PhyHlwN+qeZCx5D0WQLvlid29qfYOyFt0qypux
p3lTO5eYv5Cj1OgWgBknRfeddzZsw5wdOQQ4YTjzc54Ya7exiDIj5jl1Nc6urNxhZOlxeZl0+U9U
aCPHLitbor4XpIBXsWDgcv93Wdv5TAkf0MpffQXcil5BDm1kIwco5w+nbnnFS9Zi8PR19fpzo+uN
ZxYOj2SggeYQ1drCZQGrWuKTUu2q5GujCXKt0KVLuwhwyV1uBSFDHDF13lg/u9Q+nOsmMjLFKeMP
AdJHCDaEVTIfO+zFSRb97kyBx8yqKaAF2C/5Mk0ZYvhU/t8q3BX6AboY7LNETfm1ES0aX8PP9xph
9nY8janqiZcCUi+wKaVVWuXMMLapVlF35pd3f5SodXrvODxU+2+vNCnWtfUG4PJEt2jTKfBtcY2b
jepheh4IGkKJXih33LkfX0cuTYXm0IlK567G7UxsIKkOZOwIfo9SM5Yj0Cd5sWOUtnN8xf8DmkDz
ROizQGKohiHjHNDas4gov1GRY+kw/fbJuS9LEUANLY8r6iq7rUgtxGbTmPlgy75OTdsJx6KJSEQy
UXSqTi4XcZ8bYkFPd1twtZS/F0Q+61TDSIQZ/3Qd3UqU2C3PnGBP4q3f9KE/pPJf63ZaW6m18F7K
zaIfpXuAR09NGbBDsE1Ba/63wtjPw/ClH/s+HW9hMbffi9OwezJwVL21hGF2+sg3jCfmEnaQ4HBN
h97vyNqNOzN1cakhZwtIUOgVNIcQAv2TwL0wjKr2Kie4jFwZ2mCwaSEVkd+CrEcgDdET4ft7MpfI
PG+c90oWlgK7o377Q6pdDh4V8jEfRGRNCuwuT3iuTR9KeLuM1Xwa20rsjIpmQovYug0bTzo2TkA+
uskMqKVZYCeMht/9BeTFUuxcYAhzegR9vSMzDl772gf6zS1j+kEkVGUmh2FbcEUJinrok9eUhykr
dPKjWFI0l0LrL3N3DiFnsPad4I3mmXInWegzfimxt4gCUkKqQc4HC1rQXZwNiAvQQtLpIlQaDhcy
DlzJ5qwHtDgUJXeu/lFCVd5BUrXaJQVYoN+E1qOzGRasLsosPB5jDmIO8DCdbKdFSbHX1igcon9Q
+JQoHviZo1YwguExHXBVv4eb7f0TrgkTIBva70o1azwDnO4SxIlZAYpry+xKcvKPGo6n4iDIhx4a
tZj/mpSAh9CFnGMs2/0Z4FWIRKbqMxfMExJJf+2GzrPghXHHfDwa2QAv7BNzfNEPPgwDGmV2o77+
D1GNGaR0Tz3vCthB5vYpNeSJJEIm+MpeQTdkQmP9mj1dPY9E+l60YV1U5eVTIo2BmRp22ASsOhJ6
xJZFimqCV4XIuaR9t2KkAu1dg2Ut5iTbNKVk3+EQ09swuGtchg2zkVWJy45A1RvaEWEAIMQMmBVZ
Uu2Tvu6CM7IU03ZfhNiX+NVbiVcAvI6qJCqt3TmWzZ8TyMacKdZh/eJ02dXmZ33PQF29dW+MfaAu
taMve3N/qYbgK46HEXWOea06OUmATJQt1/UwUxGaCHrmd7bKrFQ+otfZiuATPfsi8pHVKtI3Z3R6
2gBpY2rO9IB9UuRm7inzEibmx/450h29vTp56WO+dvJnhMsTFNDgtSWrwxYvcVd1BbVKhmsXdg/0
gzfMi+hEeG0/vXsKexkL25yl7OMOMDugkNrW8PXR7+Nfe9SBPS/mW9e72Apsh2HqG5Kc/hckrrCc
+ZClmkqXDh5J/0k3n3fLV4ChHBCWhTZREBU8IjlZId7gHYl5L6EiSAXJvEeDGfWk7imMcqU5/52r
634UqG2cKTyBN55rEf5kqnVYVAd2SYvi59usDEtw85XAYDkcdR45gUMZt4mPnboWOOscooUfWX+1
OBSQnZXfCuajR/fz/NwZDXRhoaGq3DWByp/bPfeh9jzE6p/kS4pWo/991EtiFEUr+n4gKWIFxQQa
WZ+/Iyy6Mv5Z4HImXY+uG71Nq3wn9LS0mCGi84PsdbQ2NsiJRZwEYj4mpITzS2XR+/2uC1+LsGr9
BhX9lT/MLJ84E7HtKV6dABIxdeHHPIyJM5R3/KllSIwpSvdnLirDZRmrA1EA3PiFkfFG805Bfj1Y
KL4rLB9FS6UN5pvuBONEWXEN45EmTx6SPNjDUmiTj9czW9c2q0Q+5UX25E43wHVIhD903b1pdw+6
8q2tzfdfJo2ok1j3mLbkKgDrUGhDmqGgrsW+Ut6Y72wAQaM5Y+5Gqy3lAhqE+d1evNDkk/mwYWeN
t3AQ5MYjmzM8XqOrZBQwG2MtjlDtfJekJ1wvejtDHx+MLcTS6pC59vHX0PRpwhvVA+nbIQBpJAXS
8yEXupZe1v7JzpgT8qr6nBf4UfspvcLISkoe6xNXCmFbDer6clS274MjsDjHqUlUE8ZsA+QaR2zA
HKJ+HcGqMnwYZj7zzJNGbog6PSWsn2LiHuuwJsgJ8ebVoLHgHo5MDsaBLfxTbLZ4M1UH0uqi7BjU
Wq+Q5gjrVR3ejAFNyhKq1Es2jhq/fWk1DriZzpn1kGFUZceR0T2KiOqFKVOehM1OPYrIsACkEbei
I+HRyzXRh6UxG2AGGSWNxaGV+ZwIz8rs0B/S2JJCOtbou6NkvTnaznBRneM4skmqWk+n5yipTVwP
/kDZLOXeAd3J3vGaeyY5GxoE+Hv3rVF0nSqh4cvGyyp2UudmF0O10A0wU44dhnKFRFMgymBkFxdG
0pYQel6W4d79TOSMmhq/PCBdeZarpcMwR87HX6D15JHRKzFdqNv08K0l+PPAcJOFGaofmGQE/5Me
+RNS0Ltj/WrGeXOZw/EjlH0jIJRmcmJhU4s1m0uBkSieNM+7Ed5fbo7MhANQaBBpVsIqQMsEcbkQ
5kJ6Zo7H2r6tbMoWiohWIFI649rQYOeMzi5S5QZZUviL5bxm5Jy3fBJzkFKO70piEzwyjkewVOGI
GTjN33k3lZKEtQ4AUTKzXHV2khFmSV/QA3DPb11OTcZYsjLFWe7zbtHwAA8PrO3ty8p1OppiUaI3
iqxPZfSh21kD6+CyXW2JVzwqSvIBEQ6MRM5awKm5GBzOZbrPtbPQz+F/Xm9iwOwTECaCDzMr5uVp
CWUwNx46EHxhYWSMlh1LD7lSRO7lKsAsVySSqgkFRsJuo4vBiDZhS6+Z/SDFr/rSZ1JOlDKP5bvB
i10MtJGMSi504HoBpOa67LTXIkVbP0RPWo39gjZbi7HUEW2clfQkflxRp2wj6dW4cv2484IIrTvU
2RXL0u9Jyu/cTggGBvLgjvSquLvlqA8lDzbfwcGfgf1v01m6kQOXA4j6+Xzz3JsSJ8fo+8G6P9QJ
CYwV8nYlJQclDRWbUDXfz/9UD0120WnL3O08vsYLQW3Th1sX958WqZJm1oOaGVIHv3fQCMjgNuag
hcYsWXmojPBqWRzDCJcnyVSGV5i27ucVhXx42pKXssvW5/IGKAyckXRXie0lgYcx47kku/e1o08o
3iaEcUCDw4YbYlXffgqXrmLkPZgpcpB9frvH6Qc9t+s6t5u+k55X/Ys9iIWPXhc1Vvg7x6w7It7O
RY1xmESAdtr7rS7fUL84PZekyTjyoUR9lTUARY4ZIoeU9VdUaWRpISJot0gFnRYnVLq16Mm411ak
/8FLPAoUNcESuvqyExUQaWDCxiUYAt5LxFKsmuSsdoPB0o46au6Y2q65P5/VIbO2NRisEapB3dxc
afvbJz+wW7eTo10qcf6p9CgWMwaTv7ZMmvZmXDP/gu0gcY9Nq/kYD0qQakIKIFvXs4YyxVVjop+V
O5wa5TnyrMCX0Nf1ngGKNKjQnSZSJOfWhpLAOnbiebDQ7wyxydKG7zpOKKNO0l3h/vtI124DdFyH
Vt6tK9Rb0wU28ODyNJ3MlcjmaNZGrkreljkn2x2kT/HdOG3va0Uw1ZLIXe35KdqU2YQZjtQ8UMLJ
47Vu/5jJbPpyC6hxdq+SQqp0GpQKxJad3YYNmjMOxpYSiCZkCZCf+NpHFyPfZgcRaiU3iT1WrQfL
/VhcsZu18AojrGhF35Db162LKMFdU0aBvVrhyqtwbXMOJcNnmI6+aCIRDXrQS6YbWLVaa/AJ0Nfu
UHnNRAhzQ9HtxLU+uRVVmhIoYpM9mx8jlyV76pemKri0ezLIkCwi0fnuTQ6SN4un2qzqvG5xsdNO
rikzqNozn0auYqTrEWkueVyWxEv2AIMO9/UNSBJjI+gyDDDMY0Jp9ygUFMIKDouLRXlentbfgw5c
gAIg/S/mHQYw55uOvkeJofx2wEnanGgMzhdTXcMfAPWismJHpPkz3kqcrhxe9cwRBjwM57PAz/lh
YorEUo+eCy41EwAy0aRd5USJkVsPfw40NxSpE3sT4bVlzDAjrIpcxRbzoqH5Qk0uqQpiI4/kLu4N
w99L9UVsxy8mS6mRsuvm//LDTA5pZrtfxE1aCMH461pFdI7Ok/ZDRyEa8MOuKF/AEY9nptM9TKUp
TXTuhQcwKgN+532JV0aobLgOsPWm7F845GI6+kxU2ulyK63FMoyaVxUTnmAtV2amQ1wXyD9fG6H/
KDwjhp1f2pDDJYAIUYRfDuj6XgD+1WMSyBOfmO7kI7d5879o+VAPs8hqNm3fFCoRa7S6q9PvWpgd
psxzvOXgQzYVxKCHjTKZnRx5wDBv1wSlMCN07m/xNuxYCeWLwRdc7fnYzCK3edU9G/lulhdH/d/C
IZv4sN1GhTFPSYfLOYAwXlx+RKXkJ6eLQ0QTSM8/1MhOM8BmDPFM+LHcobzNrgBcYpGgEli5TsU3
Aayd5deB3o38/AM/lM+jq7yX8TfoWaoDGIFR987W6NlzuZG3VfvuKKZKemW1fM5GeE45hfTOsL0G
V+BN15LXxrQjWAggwLHKVmQG7jwe0Yu9OORxLxlM57736QYIrMLDWatkToduNLuO3056TCjFIpQW
XeZfjeDlWiP923bIGsiD7M2Lf+3nskZ1mpSXoPqr40hVnw3QJfvLllLiIFFfJ1ew3iTBsaFrOLAG
QJk7RC7khtwBAIMyehAw+aLsmLIKa0J0h18umcu5r7uohFZo5fhSThoZ2RSoYrHN0fheKt94Y9Rl
MkwrIiCNOpwqNDC36VIlwu4pdrryOLI8jIuwdTbdfyLsWBmPRk3qfEy5lZMkGVt4I7V5DwSDCCTI
oCH1hatV7xJ6qeeoLOtu7jS5pou0OL4HerPBJTqvRZHQ1clMCsySQPX3HQIM6PWTWMHXK4d9aC3o
ViVhmwjaOHifbufNh+koVgzXxwJfOLUCsznWr28SEtw19S6WtNQtfxrgExs1xPxpFlDDSbe5VqXk
ktPNCn0oMZzS6A2BzSFXhQlE9ZEdyN/kwOcmgQ+y4ygz3ryiKOD1WmpszltqkGn5bAd+ONuMoq4h
YhCZ7ORJje5+3uXhXi/5Gd56ljEMBa7hXIPHr1nO6Cr6MmBa6SyTVL1tpVx7sItRzvynrMBznHGf
WGEZtC07hbVncbCmr34es+4xsOe0foPB80bWOZ3cJGLngsVb58ZCsIHECKXp8d6+4Ut/QFxZ+add
nJA/jL1O/E8e2HKOcK2/jdO0arhoTKVMxFY6SejxKOUKyPymuaa/tclmnle2i/5rEuAglvoi+CxK
tI2zXFzRN6bCKHgojNfpidbkW9xheryT+YjKtWpNFbDQu4I9XUPWu13tVJ6jpaMPrOIVEgzglNaV
nnLFtGHxJGhbz27t3RBIoC72w1F+ugIkQ7niksGr14DhG++kgjHDbkbzlniohisBSnCI6FxBWnL7
gwLKTnbYHhPgskmmEj6cwcrZTcPSe527J85x0xXl4+xWPZpLQE/1HQG9ZYGS3qESMudkRXYRlihz
wbR5+a1Db0g2XJQyrFX5eR/yOIa1c8sOs4xdEIsmvufQL6h3+hexIzH7tvXfaNVY5n2hp20akLji
xArsOPYXkBzrgI3AoF+2wFoHgdvEquHcKj45SL9bBiF51BfVioK6+/l/6nzgaptleLrlSvT+VQpt
PYQTw/xG2m5kS0/MgzgGZOgqHiYD51pYI0Ac9kRXKoU2PGkGsqHoJf+r0tVacbOkmzmTCaeAvpvl
Szvcx8opFAbKlMXgeWuQD8RSQsay4WgHTKHseHcLQbk7/NHJih/Zn5IjZPiyLXhVYWT2YDBIt/e3
oG12d2813coq95g0+XEWNTjU0XXeEi/cf04v+ikTNVYbYe4Q6XjlMCfPtK9YcmnpJDK32ZexvY6X
J1Ctx1WsEhNRU/zJAES2GPmCOv9tNVSCWhQxnShkciPbe3teEGSlITfzFrujjzOmmTjfiGCD/6jo
xqfbclkkB9yOoPdKo1IosF2HV8BoMEcPVLhMuwcgDDOByB6Q4vheb3sdS7H3UieMxsWvEbzdOcy2
dQuo91EoMEAy5DYBwtu1GpKkqveUFcYmAfMeXDeo1knkmOANCcnzY0FBDTSr5B3NTqh5LelExD9+
G5vnaa6ZA/OPMZLblAEKEzXR3aAUo2BEpBTyrF0Ng+Cd3/t9qKJQyhoG3vj44ecXNv2sjsVj7aKQ
wn3fRVJrlNTc4aDRfwndrUSFZr5B4ucoxrRVd42m+8v1q0J+0mOsiu/1Kxj2vS9pQqWWicAvgby/
woeTNflcTVIzMZi8sMnf/uyy0EpnAf4Um46hJrxzOz/uQRX1XOE9mm9jMgpkMc1M04WIDsdzrq9P
hLaR9BXznJIBeX1IdIrrbxBxeYvmu4hmUKJ+Ty2OZa1xtZ/VVSXeAyiUqyyVrEyz92S53Zk0OEp7
Uv95BFIgpDRVHM2r5QylwXWoDoHKrTcuBBSPGnSPQZKxxuojOW3s3nK9PwBjUmqLK17rrw0649ze
1sE8SOL8v1BWeSXN+2if/faRy/5K00XrMPmU9W7CXH7C9UjJvzyCKePWHmCmOkQaAea0B7Nrs6+f
NiBi8iRxj4vI0vueGBft4F3O09arqNraFW723/0I4X41MOjorjKe1k0qqjDkasJrjanhxOZ2qWEZ
Ynu3bA5iZqBRhntZ0R1Fa4bFSQN8mOV6tzwX7RJDKVoFius/BdmrDuePQ3ekQGFFmbJjNnPxmLr5
Q/QqG/dha0Bc5Z6xhrzhJcqtuG8n3qYENIT/YXfgxI6/s2THz2magFXTYh7pn/zN4yEJhyi1piP6
S+dyYUHgOw2qnkB30IT0QE/2jMLDwRKbXoGauzIr2W2e9235gpFXzAUVPRqprf09o/WZD1wLahRE
QSzL5SO84XsCZCXC9pEc4bBgHlDY3lis3+NAAQvSSJtT699Fbadu4iUl9SzMLmSVd1MOY+LQjxFP
/49a0lvF/YoD/IR6ZGPyjAJPHEwAWQj9Otwv/5nt2MjeHtk3fSxhI9agJeo0qCSp+ijfo0h9qGuM
NGIY3EGa6Ksz63t57VXC+9/QeOd4vP1/x6ItB5dKXGAzbDqJRLhep/2UwHpWKqYI86HXvMs9Tv90
FVb0r04GRQYcbrzcCQTKKBQw4FLA15XvG+qJI63Ur3N92a4qhAqNpv4vxdg2Mm5a5q3mRwSc7d+K
2OLyD/0r2X5kL6dYxk4x5gWIxxmdsZ+9VH1GFTg9PPbxstGE4hIxbyXSgTU4hA1DBkhmWWX7+zGx
UOxgVe8mCSy8MRElEnIfrX06/n3SRdNX82qXT9i41Rw4KYuxpgXn86n1rGjgXtS+qEbWmHvCx7VN
0GtxcyLyaWzY/j7GiBT5zJ3VzVMDh3y38F8QFZTPJOMg/ZfUMcMdnY4jlE6p7iubii4Re9V4k5qb
G6+sxozYP+m+E2sYcPieKxr0GSs3wx00XaUW07Zl/OIzabNwa6vVPk6T/TCCedQArUh+bNIyI8b+
bBEEFf3Qpp9wcJ3xEXLOEEYkt6DVNs18rbJFd0kFii+y4ECs5F4/NpjmMo/VcQYy+K/9KJw0hEsG
LKLIjZTHeRc4Tf7x9OEO5bL5WQBF4JQqAWxJinwdubKC8jDsf0A65bVEAo6Px0uej+6h0WeFDFN5
4ojt/T+52xFp5/vYY/8mIOTKQHloei8gtZYfjUV8fhBZzS946FmYRaujN8Pcax1gLPG5U/h0Iism
wfOh6swHuMBqW9leheT+KBFnJ24y2TAi+VD3/SqR7rUtgdO+9xM33HGZIUulwruttzL97sKwvKGM
GaY7WZY5UigdGslx+VmIEppkr37xFe8/oRUyXwVpGA1lUSXio1qzAXvWdJceTjUbEDdz+yWE6BBc
LOTLNQn3JmYWI1v2zU6mxctuHKz9DiCAsYNaxIGGXI/Gb1IUq6TRihWXQThhHoB/OgvMqemP6eFP
HonGHSyfhFI+FbEnhLVH8ODjBpcJKl6rprtk9MwOF5L4P5CPd5rZBE/2N8PEal6PbzkpWC6a5FTp
IRzsxpspCSbgEajCoqy3h8yo+DDPK/bnyVIomPwRPf8pM+flfgszE16u4r+TBp3fiSuO3YZ7Fl0D
C+JvJVZ65/EktNh39H8Mwml/Qhvs8scQ/bJXqMIgnKmDzKiquoiCU5zNIy/2VZ2Z4FmZIXqAS4ZW
4aPb3E75XUHnuF1MRozXvjN+8lziSX0QTW3ZiAWzQmVkQGr6/8CyhlWytjZaAGmqikyT+qCLqye+
3Bc++1z0WTkF+3ooMrEBIi7a44n3c03L5oRNAdi5N7/JiDiAbQz7HkFbYKC6xIYuRNwKnqxXCq1i
czTshjy+byzRsllXIhCe6LWT41V4vyri/pAFvtTY69WiIke3l+r9XMmty1JRnp4T2ESWtwXJu8vH
vHQTS5rsCnBMcELFmJudYiUgsCuJZ4IVLYX5MlmiYXAurtusBpTCWAZtnNrRAIgEx/DtVQSAAqZC
Oqxd0ifDlPTCN9nR8HmScMyVyxwIBMpPYAHiexq9kOnNzyX5CuGvz+mTPLuYhatrzuRyeKOWysT1
yF7XlT+YJL4olCQFPmps5F1IyqRI88Em4rIm2QLkEYmtE3Zjoaq1Hh8Rgl1mrMffhS82d8A4vVO8
iwWRFA8/5J1XUetRomB10gIwNvfaLfTVuQ/tq4qlwpGh7JF4i4+YC8o3FMGa3HacrSVcI0oZ7gxh
uld4GGklTqAQ6FSzUURWtz9auJjEUcd02OfVotz+uLjBLt7nJ+f7PZZIjtH1CK7VZ+n97oczQlup
VlcmnJ/06RfmMcRIpiF52B78XWcJC9Wp+nmg395+uoBZ0rFheLYM8K2c514p0J6K5fRCbaORH95c
3/+XI8MeOGR1CdLGnFpYglalt/EGALGS4X3E2oH/sOHEwDp2k9aGoXXeEjLWVEdvcray+7fSwe7L
deFJ1jYxYijpuRMTGrCDlKx1gdIU1anbibG4lUusD2KWLxBK7n3FfbRVgwcH7wJFOAYg/ItFk7M6
4aAEIBFYGqlxj2zMyptRZI82srZlJQ+zZpwCLXz/iV5YXun/mZkCLkgx4OIC4Os1fG+56GEz/IOe
nK9JHEEwTpYyQKIiEzVEz//MCOKtAcO+N0Rf7Rq5oZPlj6UOtk87UYviN9LhBQ5YiAMcpovEAqzG
WecH2zAUdOK54sJIVUOqk942SWxXdY13HyFzijR3Fx/DbfnYJxBN6yWhLTircOYIAV2rd0SrpHwN
+HGd+uBWEcFpkpzMadUo0+xH2IBQRki7IpYVB+BfVY4yA3QhKgzIOykTt4FZjkjZvYBFrhQxBOSj
Tz5wBREHwJlspfEJM8zNK08I+XyBaV3d0+Wn0aWUhCPphBI5V2moegGK8a/SzcEbUSVR3AEt4V22
PzdD5xpSlmzXlAfFHS1MkyBeoa6FN6aNxYnRjAMsTCNQYl1Ke//GlEA91UhVa8dLzUQqq8EjCQNd
Ui17Am6HKaLCjK91oya/xEt6ZMBM8O12Pq+YN9rDkejaSgcFqkNj19x2816gcFeEY14Njf+VRQqP
RNWrqCDCawQNDfxYKNlBg/99GWTcfE3Ue38pHhznARjeXwyjwQrzjFCi35+QF+h75xe9VpM9Uvzc
OkMwpOmy7dpipoaxedDt+m0HVLdk/qGRFokF9pTTxsD+8TD+bsEgZWN1m14Jd5GLypP2HSiDZGz8
nMrt24uOFwxE/rIc8GcewiZfkJAUmR2udD/08FIprsRGdWqaPMNgb8MTGwBitsEjKeOowATSKxdv
SbhSQCCcoAg2N63+av0mp/NGCY+Q6CnW8Jd4+PY2FOddNqm5eURN1LKR+NWiCECRr7YX4Q9/O5tN
Tqsj0uaGhgCEFSamqzJjwSzojB+UY+JD3KN3knygAnvREn+0dz0l1y3mIe3l1p+ayWp00LSY72rn
XamYN+IgpcvnrgYkQ0GNZ3/lVzIsa4lTQ0nRGA8/+7zEa11nzbiW8qDfBSNm8Ho6NovGtFj3VC8/
wtvIWIvEp6dMIviESZMo2ePXumzaeQiYad0re+/PMDy3vgwsP3cUTkMGOFvMrrEv47DzkKxhDud8
knzLy0PYUcxuPMvotbFgSQsA9FjEcq988DlA/v0FQHrrL64humHk2bhnmvo+ST9RbEXXRI2UuhFA
K53Z2lmOrzewj5L5gLEcMu6F6ihdLml5yqbPM+hpEqbwJRLJtE+90/X/B7QcbhXWa806ksnSub/X
5ZMy9OkFZVY64RTiUE07AaUYLSSEcl8QinAKtoEv/dljhWolTSr652154+7+0z6jkAfOb4o4Nr3m
lmUuu1iUqO0Wz//DWsY6sJtc3YGIC50tXMUAj7WfpExszNf/Z4mCF6hijUn39DMNIGGtyI2noZE0
+vp1STXdYe7a2kvJiHr0i2wo/N/knuVm85ManYQf0f7SdqrPSZoDZFZZa7LRH77CfcsZWLjkz8pF
3TXk97ndKb3P17uMwf0Ozlx3jYYO5206FJtNaU6gkAUYS+y5vb1z/d52W7XY45raXa52Qmy29E2f
4TYGd9kUDzZ5ZbE6KNJRShR6enRLX4AJI9Je3b7FarmZAMH3W/7TS3ONmbfKJoAiqoKAJkCv8B2V
w20daGn8CMcr9U3cK7i2FkkU1B9QcIO9gbwF33F4sodvRWnHxf1Pd6JdeV3voXCnlewf8/v9WC23
JUje1j3bMl5V0y1YLIfvofCtjkAbvOwF8Kdvhy7ESWHpQW7M+zdHUeyKzi2WN97KxwDxMpQUkYSB
Z/7AfxrgK4hOOWKKP7MynHwEZsOcctViwQCHr+hfnvzrl+ho4zcMEXzRYUQ8qzi09tgBxb2kxQFl
j9exzNjohUDdXRJbS1+XufQSgt3egEd1uK41bLHYGHfDE2jm+U17ID79SDFC9GyzbsUd0O9ICUAn
Pw43Do+Q7HzOEIfQUkwL2IroX/EB+4qH5ItaN3Y8ZWDyZcgdkMjIXuj4ymfE2knDeN6GjOgGgnuh
+ysX/TJJMqu2qRX8qTP7bXQxLgqYUbDQr3RrMKOKFdLOqSQvDf72WRxOJXt0OUxrZx0GKpisIrKR
MId0S0scFHaXyCyC9OSuDTFJtgBX1R0n2xIStA53QYOrnFgMQzW6Y7O5mtH+HCMvIU7Xldy3aBvy
X/4sS04Z0KABMU+3wkuk0BKidIDL8JkKHE0yFC5NpmxC2WqlT8SPDh3aYlH75NghLL9Je9MQ+mUw
KWsXxkAwyoyPSCYJJTsqkBa+zwN7v05dGtgC7AmDC+7uEmyL61kmuHFp4sAb5sKjhXXwZIrH1lEx
x+oGlyLme5wyNVy7dAl77mpYD4m+lqqz7Ir3N5fPrPMIABEVWNEQ/UPXgJldMbGjT4PgLDmop5Kv
SvbfJ99zWIOdhT/IAliyVxeHfCnWhtoismYujcTQAK+S8aVI+YyGvbIYPky913MP7skvMfAwkCD1
ozCU3nYIoWq6Q2LII3BkeMFfARgCtwVTVObN1Kbdy8Pt6F/qDbgqlwjHknG1d6hu5y14K/8zDKVa
oK3nTUcGZ39v6l8FnWS8DRTn2ZvsIo4smIeaPw/MzoIMAPi/r2qXKyiu0bs885ADQBkSRT1aBeli
u9i65zgGHAzdQ7C6rSeUTqY9ROmdSmgTBnwk6CTrssfQ6ZTyTJWthkSfVA2b76loDFmtGWMIolKQ
5YIMkGw+bT+cYyJG2zyowSr8MW4+RUi/cr2+//37Ol5KstvewilApx4O8wuxqmlgbBOSlCQWA7kE
H+N25Fo7RgsQCrKdZi0aTlPLUq1v1wagy9oKYaL4Pud4q76NCjGKfw5YbvC1OHqaIT7wM8QE3MO7
jvRa5tZZ9Gw6jsaPxXXgQ8Isrb0oy6UlmE8SmCuxOsDS6cE7l5B5xefgPLieVhWsS7yo7kXXorrh
pBDcyVqmKf2SdK0I4kyWIc9/iY6Wi0gHvdpmRgdX1ff1S7ozsk3aUtjwQYWPFpBNQrBGJpZi3ZRp
/7/UsV//cW20Ihs90MpseRvlRL1KXljSuRFaY9N1Cteo4fsHSm7ey6oEdX3kDREXzoqzt/+DIG8h
U+Xi2lti9rdIb2TL3PF5kQJOosrgnSWzEtMomhXDjOfriguGdlXZPX5wSYUXh0ymhbRb6mGt80Hs
WSOTvqeJ4+GYKlXyZ6r+3+1uOJYmnbfcs5JqDMnp8BBMBafTB7xEQ/kmaHlm8Ox1G5jlZrfk9KWx
7SPq4VC043lbqZX2oHGbPl+jkNL0oElW5E/5TGhgyciZ+6hn+ZG3BPehB2uP978/hu60Y7pggoq2
hf0g7t7LFxLzOCDTawjMk2gcq9gqV0I6EH0aUsTv73LMv+71NlFJ57byfFdavXl9PAGJab5/UKak
MxC8Ua+4d7dFwWt3DpsY07/a6x7bK7y13wHvWzqRaK0gU5wWN1F/rggI3n2A5UDwGeLfNZ1TXZCW
t+2xNSlKtVDZQJFQFQuM7zJtAXcWjkWoT4TS5q9QqVUsMcn2fJFdMoA+W/eM7FCxItUiLeoSEYhf
Ff55xQe7yJH/MynNqt0h5PRnIKm5DOTblfOyfxhrzmtGYl50hvCv9He+ZBKXwESkJ06bjp29EWr6
rg+464jbAuvej9JKUic77hQIZqM15EY8I6klyFj/lPWtxeTtwT/O7VToRoVv3Kx7+Jwftcq0tZFq
K4VVvDEuvMuPZT1LwPyHwNsF2eKABRN0z3hh9afD2JxwnygJOdF4DLN3e8WjKeSY/Thrq4eI+DCA
+HMRrblQ2RWniaJM4Gc34eaj/9BuLVjMksgxjQSewgE+55H0yzGDWJyotyzyVXVydiSloNiTTU6b
maaoaJvZusf717sF9YTx9OZBomc/K5vRZutTZ+6vhVDac0y9QB4wAFQ+kyMQxOdxnfd6MxKZtvfh
bSsJ9KXfHtM8s3OnF3Z8LvQ75mz3gM1cf+fjt66Slbt4vQu2USikTqR43W5BZppYVjtdo/JhjksS
5hbfOQKs89XEIpHkGdY8M1xPBnaQR898HoEBRYGaysmABHIvYQ0Ku4edZtPMZY7lsil31EwVxFs5
C+elpaC889BrRnXRWaI9TZIvbrVGenj8UG3pZPH5J/JRDz57Reop0XCBEILWDxU8deXD5yUwtFKw
yDsFHrA1AMmF3L02jAOnuoeuYN+w1zX60PaZOxgfv4yjMZSsTJY1VBvFfowBm4AGV04VIZ6aoQIx
29gTq2BX54PXW/vLsDLfdnn8WQ8pVb0dygdbSJS/NIqXQbnYdAQQRAt3nTL2YOAODYCLU/y0Q+v8
rwWxLOcyzbRQyJDCEc1TmMBaakskE3cLYCrVljFNh839sm89qdg4VD/DQnjwP+SGR+bNrkDQNoge
g1gQRi/jpP4RYI3lekCwy8hjZ27mkyDm3hnHyGux27z6dohU426yMJkTes6qbd0ZtB1yf+TC07pZ
FPHU8jNfdCSLZZi+PrCWIeKyk8Ovnpa6D6Aqi9gB5WJU6J96SThp6P2OvtURbsew+/2vPcVm8uLJ
XEFdqEJC0/zc5FECMBwDwHaQ2Zw6HPxUD5KIwLzBb3f3+Fj/g/Ob9Ja6H7jx+n6Co4EfAu2LGhec
dvKhxDd25Qc533iP98korsuknRrT40/S6ykTscEte4MZ3qOi3ClbYaJOuULXxWzU5cJkuovRBC8C
gC7FwH4VDbNesA7j/+26tHqu1pIcrG/V1+d2Sx1lFfzB+5iXJ/xBFqoZCwqWyZqZhCfxqr5VjyIX
AtyQMOfHWZXcKQvvum6M1GSOLNncZ+EOHAYGgrHjAreMBVIZsdKFfP9eBD+Vh6rZkVxm7AsnUeKp
j1DP9uXzLnvwytUTTcxIBSE9kkV30gti9gyK6AhftW9n2c0aLry5q6TcgODbZznWhuH0EJ3hON3F
UUmPWMhqvRzLuPGVb5Sn1Wmukj7EjMjNsSlMHBV/HgjxzMUDqcggAqG1vkZ9PDeQSyUKKdwJdSG3
tchxce4E7NkCzVcXoIICgCvoIIp1tbl06NOQaU+rFpVJYUZ0F/WKSTO/kr5NSXVfElktw1Wmdwbf
EEkj6WzhUIVYpNss44HDzjZ63px60T/GqHHYkV3qEdm9HMDD88Eq4vupcYFIc4p3KN3EpJhN8TRk
J/mrO5LU6YagVboR+Qe8jiDQRK0CmueqvfvRh02RCiC4+p1DMtFgAGSsbOmH854hxIDz9tl0pKly
TNDsIM3h4FnlvCMn23mT2s223/2JSJJltzM087ir+AgigEzneDDbmpul0L5gcvkFzTfgsP5wVooG
OzkmjGM/rBg7ejhSyfJZiPP5dFqJ3AEefGSzGpcFkduGewqxdzwtrG6U4Uz6IqcUi30aiamYS2T0
Gm6J7NP1NXbn5wLrFaBVz/nEIfMG+0q27xiNaSU0cwdHSeJ+c/fh5DbanUDA82R7WQGJOpMgmn3Z
mXfhXXLgRrzts1IJWTpf+J1bOkZ0TJKt6qA5L8o3qJSs71EjScSxRU22YyZaaDnNO++uksQfDvi/
i5A28DRFVFguvAS/tgbHYko5G5niHqGlcJF3Rv+hdx2CkYdsS2+hMQ0hROvZEKarJh4GSjmLwi8h
avuow/6anwdLLAfxbND55BUNl+nElG4LQ0GRip2e3qOI8SvlxnEkZOuHOf8dxQWqEWeYdoZgJb4O
ORmDvk7/iwlk704t7rpkdnSRAjNO4A1+H73vJuTlIoxr1d5ikRmDOjj6HMg92i8KJOP45Q187p6j
xD4+Kz7uKgKouSIMWahShY4tcLmtatCwxVdJcnB1iJdgpZUIMnklfMX8BPfdzBtXYkUMXdQwPski
SZJYPqgyItbT6KwSqoeHToifauxz0Su3CZPmGkoNhcQ823UsFId4gUfDF9sR4ykSDlfNQbJBP+Lu
OUuRSgXlyXGHu6amjBKUPV9Fx92SPSFCsaYMM0WBoHsWbrbhmKTKwLRCBpVXe+AVwTJ51Oibp4Jm
h/cGQQLizG6iC7Iyog392DJKuMpDAcAylS9plm+wmlBSd/NxD0pg65cJA4ffzA2+hQQM4ZOwD53R
ipClfmuJ0XHFheVC/MFljXRAlfQ02OMY3rZNzjacmOroaJbUCHa0f/or2Y7ZK3oo3rkMgym1R/3a
R2RI60JALTlCDJWcBOqqBFBbuB1jy1gh/W4iaIMzQWitxHIlinHhNxEHo0KnNwp+YERJogcfDjbm
Pc3w7E9VCIlqDkWixE1/wXpd/zilqyWMRIA82hN7clx9c1Y0ZaTEM+AEc/SC7zTIjhD3u3Q6NIIw
r9likzVEaCazptl1Vee+UlUkeaZACnvQOKVIRH1RZKEMVHlN5h9Enbyz4gtg8ZYP8exsLr21Snf6
k/ig3U4+oyP86C3QkPsBvOeH0gDV0w91pcmc4BZDLz1Wjbee/pEjjSxYCwqRaGIByOhN2SINxnbo
MPgaS34FAIML81k+lCkbAvKeI7kbTHRz+F6V5/ou3vhbiWNMBOZ7EdiMnTvrYeHtobK4uqcdgfth
OCy3D20Le7bKQxSsOJDKjiZCojnHbGXuE8mknJnxZbXpl5VuhSqayTSCalRk8rhkDioYMI8WMmkA
pfmGTql/By8IBN1TKb7ARn8EZmc/rDpToASPHtTLof55KgLL2zQquCwqS2wSeBfZ3v3EyWiybf6g
ojgX8fCs3SHJNFkYfwKe6PcCrgCM/C/snbl7W1ZjKxpqjBv1Z/ciTufNIgsN2TPr+XTLRvk55HbU
KT85wnufg2YvLj3uhGa4rik/4v5vNSoxqgM0IkD/9nPPEscXxg+qqHqtIPRBAbglgdV8OaUO18Wp
0ecSFEep5J/TiN+aVtNvIGTBIWA8sVBUAueEGbkkDX+V44hRhGRsM2w2i5cKL0mro0rRJdQxov6u
ONDCtj2KywFOAD9ooT893voQ/CR3m/IdMHmF+ju5abyrIuAFc4BNRx3SeA5SwiZIPHSD0pgXOVfg
oFiXpsATNlITS7P7DeQrit05uhgM0REAfhVb00NA2PrPZYQuhN7SLiRXuJBNfoELpoHp3GiK5LXV
rdkkFw7bssODd0pdlmgel+CJe2Z3btm7RgD1xwC9Iv/0pEOZjSH08YrGbzI04+kiEzLBZDUFfcuM
1FrjEXE19lNCCf/9LgZ8HcGvP3ZAgA2lVW8XgsNFWJJW6IHzEnDJK59Cu8r3BNCsuWvjX+dXnwSz
u1i+KU+SqifvtcKfakGcIBSKEStkjs46ojPkSAg9KMCOT9s17Eo7sKLggnuQKvdpDmAtTfOd1x4S
2M1Pucn6UrH+qtHzs6zTIqLdYPwpQW8WWniLz8H2NyJPyoVlo/fLeLcSRmX958pk6AHI7pWM5n87
TCDLtKpvwBoS+8a35OB/pTa2FPUFhZjVMPnLHRnnPNj+WgOrJJNVZK81RUaY7bZK59j2RAqxb7RC
ZdQX7IbyR/vxRmYDGoVLkt1h5zksre+VIacB4bIhWKIVOVY18wnQPmyvzmCQ54HDW6VYDMc/2IZv
UmtbL6Iyi0UeEV7hNVNKNnv0TTNbj9JQTs1ZZK5tcdx7EeWVNXE/5n82dhNYjFjnAhN8A5fSXNQi
WU2nieOIvApBX3B7ls3+LptEXKuzJYhwrgS8SzGVibn7CjhyeL/o7+xY6UI3L1UI8658cMJRro4b
hRvH6HmB0/dOjOGRpZJVNFVQcQgN5yi0nWWkRQrkYj2L0j4ZiEajyBgnJMj2ik8ArDTRqr7bMnGD
gjuj6Adl68anpEA2xRjCiogA38C3d8PpFpcJ+4NOdQ/o+vQOKqvaaBqWpdLf91rVu2FpA3/W2Ted
Iqj9QhTYoNOGxhit19HFtNhxwlQR3aFYm8LRfI9X6ws1yOKaRep5bgTxhuZWuxjTJ2SslDlC4qNV
zAUTXQluGd/f0cK/6lI7iflPg7rwZAQ4LC/B/uZmUn42ZeKfVXilcJ2RQBgMbiwyjb7t38ED/T04
Q7gypFgJ4EmAsvV/2nS6Eq/Bzd1P/b0S5QYpF9izmT5zGP0vGzKPiLza+hH/20ZIGDVAtUnCTLZb
ZKU4xwA7p0VnDQ3EUt2UogzPP2T/nHDONGjae3Pv85dY/2mCBl4BoAMpdcoaAE0jWU/a34MhgrVP
ej96ugouHhFCzJ0sFPFHz+Nlq+rLQlmJP/o4b5FFSw3ag3k0kwe7+YYu/xozvFnbpm26gE/ulsak
qY0TRERQe5iuQDughX9FYsC/AZuELD4LdDib6p7cAO08NwSPu0KhvopoPK/XlF0HVaf4jw5KUHwm
qIDc0FnCzWx6Js/DtVrE1ftuiS08ld2Y+v2aOiK7H8tzX5Di4GrWRWI0ltICfwOf4HhJd2xJ8xo5
ReWKnCgIJ6Our58bJ28bx4r9RpkEIn03/L8alKDwFJ2l3Mgu3CYEPLyTn6b20cqOkrbRHgoAqEZo
gT2wruV46jgKCk2coCALmXCxZbS+P3m/D634aZdamYYzO2DgCSrN6fWo8+GeAtBXY61gzhrfLXP3
//ePeY8oh7B5XyXiWEBOWRy6m27NUfh9kt+l08dtzOqqQcil56hhJKMZhEjUCiPTDdx/Uh0xdiEP
XkP1jH+xvFXseHY5/9SaacGB15A9Qi+eFJOMmEIttMv8U1vZoU3Z2h0SwuzDiFpXNotdSU80TL+1
tX7DYw6qvnQakZFw20IJxWQQiba8lUkx1XZflLnhU5AyPB+o2bKWu3huw4x961daPA/3P4g/nL2p
sfsMv57dxcjInd0c0I4pR5UNdMuDL0yooP7tmNTx5NmZOIk/j7vBQ3TmcWEpJAstFNgrj5RzDsRu
S4XJWk32buCHfvy0bxyMHMusrc3A/SHmb2oEoFgIXK92VLvevLnoRzKoszmyxTK7kyTb7s/i8g7O
QfylfOAbQmhkhv/61L1dvBeMdycle+VtgskuMvgHo9140BbLMOtxOLfLaQ8lB44spk0msiHiO2un
XLeKp743BiWoFq79ngf/vsrZDdcVe43j0q+0PKu/GI9A9MHqlWcMQl2jabaOYSMWhAVlb0BOtEs+
Pf34JGpBuCk1F7LX+BcwljQvusw2UwhYQtp0A3MYAoqoYVAZhJT0vHj/YgO7zMEASRYlrDrHjkiG
kb3+UcpYcHlHny4d0Jk0cie+0lXtZjUDJXSJl6y+zMhyiFnsPYEYFo/6N6xNO5GsaD4SMChajXrF
1+nCMuh/Mxqjni3bQ/8xz3RvfzEl7dj+j+deT4bhVRgUHu/IaMw73EYrHvor+sm9KuBK4sC7zQZv
h3uPV0agHXmK5Fy2Spce183s3iZGx+Gice3qfoqml/+Nd7gYCyNIk7M1Qn7aIUWBCVAtssIUl0kY
ZnSV5sertkzyj7Nb/vNrnrbYAIdhGL6Z3GotambjauIzTYEyvamp6SFUUb/IA3T4QxMJQ44xp5AS
GkhVDaVsRew7UaNu3shdLfJt9vvIMUCyaUoXhDm4Lv661xLeK+xJSh6sc6CerlvbtINmm7oXmK+K
OrMikH+D+0LZ4LNXQNkDXB3IOCrQw7EhzwYz5VMGrk3GyVYPIEVeVbkx9qP30ytC6R+fBkXMIltZ
MthZtAGd5Oe4PRwVuKxoQqZbeQDTO34mbSWincNzJUemUf6so6EKsuRVNLL1F8wbaYfwrlaoAxY+
2Ovi0TORg+PMidp2GkKYh+uLS64ApUiS7nlwUFi2BY4iqvCDVakTw+fag4F8JXC4HswkOUyclsix
e8t+p70M/jIElvRtLlB37mdGmLekV1ZPBB7KBmacpm78baWvsIrhWmZ5xiTZXpTTuaRWwPQ6dJqt
noGi9P1+E4HwvIk6sGVuIxtVXNJOeuydg0tVHJejzER7ajcW54SFnsrHdqXkxEmYXvUTSQYKw1i9
D2myFlQdCtcZpje/7EOdChGnQ7ePl+cRdtnUpHRHxTzoEQFVYJHRurGkUGN/t26dA3PtWUJ0hCIr
B1tr/54+Yw/Mgk/E4x9LdEXfzDzG5BIlEEelsLSzb3Y2R5/aD6FH68w3dMBh691wvZ9NltylJDUZ
ovEHrmkM79WO0c49W2svoep20D404wRvOK8ocjFiNLORiALkvimlQjCqWdJKlW3q8699d9tsxrgZ
IdGQqwfNFkhO2MDq4IkPcO8Y7mp5PGiXU7uRYJGD16WwE8oqvVekdbcsZOXLauVSytEvabeSlWKk
bvWtxEfP3t0cvcwXjEgqc9bacdDhTLfY17jN3PZh29kkc2q4sZkmVANVayuErxiTtnx4UfVuxmhQ
jeXhYgza0t3P3PAe0OJdvK4Bo//MqWrLWScpZN7QGUwVxlv4MZhWGwv9XMw+YrZLEP1PVx5ZwZt1
Q7dPhtYOXNhbYa0Jrmwsvvr7es4Sh5ldaPwpX8Krb23x2oIwprV0fXsZJprLmuMwu3NDHee8/h/V
YBsNDTTz/TamvVOJsYk4UjkEXfrH0dy9MRsWQDCqHkXPtUO4h23CzDroh+iRcnaKEEEXQuvZeYJK
wUcq7EkGGQWt3SSmNp1Hjv0HxSuAGInHvzJf4rYf8rgSAHPwggFrXPLGukMJ2XwvLEXEYRw7j6GK
xjOP9V7x8ObpbnpExsZ/ZKUjMqVC5IQ3KQ+WqqOhqK1c2oDdmsuw1XtBmjaZyN7Eg5D89XMXS7fF
8S9B285TQrdS8tyG7BN1l9kCVM3E09cahwsVtVilgPZ9KctYNNXQmuV4s0XTCfWNLFE7RQuN/Bmg
QxEl8l4jtwNRVIXNepXFvkrWJbAunODMAdR1hnYuhtYWfHOv9RW0odJqEEpdYVk3V7XBVG67jAsl
DPIbfaTh6+uAPaHcG6UeB22OYnvovpdNQ7RfZ5L3QU81wzn+zpIqNQxAzSQquu6Of1/v5CQEfhuq
Ggxr3g/wvWPJ930V5wDFOoNc/HrPelTWfhAa5QWg0WNQK1WUZ4t4s894fm9u16ukTn8LiYhcKyEE
Dn0e3e1x1BcrOdTcs30KT7qqmqidKqNnYWO8O6Yo6K+egOUTei5l2OEWtFE5HMVPSExSxlBBzXBO
rnDL/Bb5MiqOEKTbWCX9HMnQUB9cpS09XqVj5qVH1Xw3ZitX1Y8/Jjwc9UORzgXVTfX7oI2kQnd2
gtPjtASyCpjszbQhnNOnCc4g62F2pZ4XVN3TazVE/kpMDtVp+3FtPvbBcW+px+wThMspmdjHdycZ
v1KnpcbbAXWtkA/EH4vPXzDmOG0bNO2UFrWe5NwJvYp0lNJqUpqKtun4MbsubsZuzEmqIAJd2zUe
TPSLc2B0GesjuI/KU4ZTNHxQeWy0GZXPgvcA/O3V3qqXqBWkcQnNZW3G07JtyqSNE7rsZh8aoBaH
ZMG4x+kZovZBqUi7P7CTfIB4hE9A0x9k5LRJYrz4ZU0A/9+WpeBei7Ebe6Hrbk61kyrfcxdhBZc5
oQdeu3SfVsaSGgJTFM0JIQ+6Pw5tCAI2oeK/cE2Yzs4M6kiPgKO08mg8c5UIsGGPxtIl1BWjB7gs
ryCCOsUuSCrF8lOzmwpWLqUMi/6T2yySQY1IxEAz9vp2/ZiiR6vndpyq+ZijLr/ZjViHnqjOJKEn
FzLyKWoBI1ro/54iESoOXe7cz8Vm+PmSvvacFEIG6ifA/CsWNVBrgSMl3/1I7rHJjaOFBAURViDU
zIzktfXQ8jbq+EWppKDVJajfbYTyF1YgjP1UGObxOlivfGGw7s3O5V9Z4IFQ5P/m5IyaTPYTbTB5
m+5KMorvgJVUpxVYjIIY1ag08pXfAwQaA37xIJLEaNIORiPwIghC5c7eigOJuZpqpfF7Z1EobHf0
pmWhBCCB3wQUCF37xGhAi0/xECcAdcd95Z+/AHa3O75MDNGSYF2khTXloTetiPjW1GHby8UO26kk
ZgKoqni6PWDj9C7h+9qAq5fbcEZDZwTDzilHMBTP4X3CqSFNO20KOR8obCqa/rdjQtkoMNxMWW1k
PjffpT1dnmBJB+/s9/SLzXmcHkq/ALcxOUWbjWkuZegMj/To7aD3MoELW2TGUD4WocCMBgWf3dIR
rNG99hZTKFLTHFZRXlKyDJc2ahGqkNIN06aQPP2hM5dQdngqsVXuoCW4ERT/JwKmd1y3y4Mfoy8Z
IMMucG9FMWoQQJXJRADB4ju0Kg5+1JgBkPDvXOQLlk09r4KorKBuRipKJ4W13XYVEArR8iWdCv0S
k3ln/l5B5IPo5sBQgMihde2dhe6s6nowmO0FOvEBNehQS3iLr40DYXZw2FrUbY0CIAs+6Yn4/Mb3
YSjWxmMebpSAQEnmxyWFgllFI9cxiRoy0c0cPGl5TLNZ8GGQyHRk8Sv/eebFEdOdfYKJNVpD5qYa
3Tka44inl726I1M+GpF2omSOVqh4rG159P6WRwzVkadALlyNY6Ij/QxjPVVciT74hOt3RVvJT3R4
1gDVUTc8ST2zBUEeYOz/kOkMGzR76u3XjI0Lt7xwfWhk/ytM890mzAQC/1158u8fDHS9uGbEHbpX
/YfxkKftVMz6jxGgOi2s7LmZeICp06mepmAkyvuxhePDRabHtSn4kS46rnKbIiYei/yuW15sqwQK
u9R1y/2qRpawB/tROrOqwweHw+nVU87WhnufKVq15lTqM0HxxjeuJHj+TwESeXtXy/TbmgDMioZv
56/plYSvYkaTjAFECD22DqjZK/IeuVIzXMGdFb+Diqj4XzwQTWOlvMbzZlbhLTU0BKVba3bPjqmH
pvvYqN2p7lmBMJdIvzzpJmGvX7p5VOqhjjYcHaKVb6VvhEG2X88tlPK8e/wjTVWcEZCCWeUHktTr
o9HIxHYByLJ1MbwSmRhMRA4P7zlePdooo1SqaJSclaxDyjUnVhBbaTBuMZ7oRInJuNdLExC8IqTj
14fcQYkt42CIKGqXw193SEmyFxRt6UQ9v18VNDKIT4vixkipFix+djxSeZ3FxQFgA6hJ9WskMSLw
XsEZ3WBzbHekXC9ycKuYyI5yTJEYvkEgfMlbxkIy0Lt5PBFxf1Fu7ji63c97aln8qxhTlyhS9LLN
4KIv3sAIjiPTlasHZHXXCcDb/H7fAU4Co5258O10QcBZE0vFPGMBTRaamLothWxSlXiMKWaam/3p
apLzE5aDuUZR+8jLF4VzWHFe/uI44QaiZP29Mz0HwNb6Mf9ze3pVp/h/WsyqIpMRQfZRe6ykA98e
lY3BOyH44/+SMBgA099WSokYJUujuEgRVQ4DHb6xf4XetSlha8rtohYz0tp5J9HmPbCN1dZvsiSL
9qHFQEz4uFgSgyqHm/TwngHoVktbFZ89lAml+Dmtys/u8ithVSdMdgiVz2joIirmAVmSknCIHed0
O8AFxSyN19L1oerPQd0hMSxsRA7qXGBAGOeg6UdvR9uWoRwVyONQI6fFgf8wORhSbJoVDTwRqIrQ
YRcUb5HP+orN5j3N4Ng/LaAlTWGWV2zowBi0RiHaAdvQ1ZZ5wZEl0KabBjszV2dT6Qg/F8P4j6JQ
thdS8+lxyjGA6K/SOZKggkkjBAmy0QCy/935tHFChy7XEXqP/T95QbdwkTQByPQIpabJhx6CdRyt
T06J8wZwVMofL1WDxJPWf7GgA+BP/aoaS+lXoGuF9lyr1jIwLbvV0JnM36NyxwrYE4LWL4sMUPny
0kVic60HTbMAsGfgkER27qkT+S29ZrviIxtAwToo+5YW9kdohT9DYub0+4PbTBC+lM6g4gLr+Jvj
OTlAnWLcQRKkWkLA3o6VErRnvftpjfbxyii9K0tntkP4gdoTvrUCKxGR6AZXaJkY/oKPnI9lJopr
dWrXlhs4F+0iPFv33C00ohM6MF8CBdRR/ZNcJ8jNnhB1+nBNsqDRQ7bDONfbPWPohmBKVoXLGQov
lexlzm585au+zwrijaW5uW4SYG+8g3BTvh2/OXGGIig2mkt3uAXiY4RVnNi/boA9GikLvE//PCFJ
j0KMWWe5dX5OWIM9NvqUyyB9cB6BfmF5vQb2wsVUq/7qiER3NLIvwCB8sNXOppM5MDJQ0SGYSlvp
5ZtQD0STvqmMOLUolY/Zf5KCoq+5jA5tLybfUQjGtRvv3CnRtApz+pn2+vN1vBjpngjSKoe+Rbqv
CghJtk1Hi5Lt2koG4Pob8Jl74WsXRKcs5kNDmEH/yZWzuk9mf5Arbet7Ix2op1d14fhL3mWdUBkw
AFXC0DrD+v/VKC3YIktQgendLmol0uIsfqmc06CEwwkFFnCNCuY5iX54y2hPFdgynJUutJf7wUqu
1VMZueXHiEcHGeh4MJessYzil6uT9yrCNoXGqI+uCj0OUGxnFBmknd90x3/Rw9+jIek1iKqKOzhQ
64bQPLfAdYiMHMMIXN35WnYHWGjbU/uUbwOPeA+kWJuJxeQOxTamVd+L7gAvqZCgMl6jQhr1dtvV
ZaMGWjc0C35mWv1sgEqVnoayKTHY6ZltlKSCmpQcW+pJFk48lOzMVlQ3LGkopsdNQYaUPJECq7h7
RAvAEwHj3UxXSyMRvAdDbPpQDsqJi34OTky2GINfKsvJE54dOxs3nyA6q2S5RcGdCww6h015yMrb
3OUYLBcUM/1r3jAum5er7rOWMdsyiybvDXaBJTPPAqUgqyv1EovaccvLq0cTE/JrW3bZ6memeB0z
VqIoTTR1qHe64yLwIebl5WvefrTDw6wOTTgzXF98wyqnW5LjlzdaEH0QOKqW7P9NdU/DIJBMob/+
yCI0H9Brt3ju4hVwmr99UdBOLgFS6nTRdqx+nXYTZdUv4QW4/6kVVAy74GH7Rk8ko/F8/9Lz1gWV
Hgx7ZKdt82BCKDQ11KHxI/CqK412CKv41XNPkvCo+GneE84Gu0cWR132jg3Fgnd1GvBI8iCRlY0d
khDf2oKrYBsRPx1Ho4UWqdCQFZMriRTZu04uzIiE4RHWax9dGdDJx5X274cl7/1qX04+se3/eaqp
BQA0Ed46fj3L5tnOcqOjgnYtBuUXBObCk9Equnpl+uivtub8s/1x3biEdsTqD2HIsOWWLza8jUtC
r4emriDprgmBu8dLQwasooi5zfwE1474Ak1PwpV41CONWtamZDx4NC5Um3byPQ9HSEH1QNTP9vxs
+DA1YIeWIX66UHuH0UcFwjrM8PJLTkuwTDdP5NH0GNILJQiG9z7Kc5a8AAYpcotR69xrltqyh/1S
jRRIqERdzyAW4s7rSAagYVIT5sIDTG/oWGYg0Q0Wv3aysYkg7rNtR1hnAxmtkpYd0EUNAeN7PhJp
OGFBZVWmJOqz/GkkZs7x4niKB17Q96RkauimEM29CkoMST44HxPiYwzzOJVn7J4Y3Hyt4xJS5y+D
0sqYA5h7wDdIjub12Liql5PPGVMl4/4paIIEy8P/GCQg1+oVRe/lABV6RtAc3FGC+iSwi3O01iOb
z+FOQ39bPgQW18MugMIZ6SyZxEqTit3iFT7LaO5b+YfiKVRUGFwUFChx8x4uuO9zfQ2LYXYemcF2
w68JEYWmOrs0RL9pxSRwmLx4R4GyvUvhYgWchIQY0pcmNPqWVclXIDxqH9jchKCeZvpzHCJ5Fdem
s5NeOKrkC/EYrSQRdR2b9E61ZT5P9S3D6xKLJmmKwPFTyKxG01XeWNjn+8i6dfkPbERhrsx7OTRK
vE8tH+59aEf8KhENqQiDQKl0GTkk5E9kWoL4QEphmJaNCu1WiioKjZ/beBwtfpquPXSo1PrH8d6E
m//muQtDUCGpTdc7p4/67cecq/kZ4OF2zQb3/cWzYcLdZRxNP9R1R3oWhiUOwFnKrfwbYVFFnb0s
jj3xFZVZo3GltnrTutkWA57H7WX3n9wbGkKi42OBHEH8p4H32ovGDPtklO7CO5Vnr49KAyyfnxUW
MJi4Fcw800tUEezuYe5KKLXtLD6/6mix1O3E0B1/Sra7o0RM8zajwKXy2zLQV0WDfiLn7viFnuLF
ojnyectjpYw9DL6CJJeaYXSYJAp6dplLj561qgXYz79AR95KiR6w9iMk4xtIDMFAxx1B0MsEExwV
5ChlROSgA/yEv1pW4eG/dL8eGRdg2nqkuGJPUF/MMZH62vhdIE6ztjAWYCnzXY5+wLxt0Xa4KNSS
vrZq9loQO7KtyLRAM6r/AJ6nGMMiCE20OHxT0TYE1VMa4qDKjqnPx9nb3aTil8qSOFlxLOYqnFVG
noYToX/4eaKcGirTzZmjnkMzWdI/Rm6IxzdB/SCz9DzjlpAA5sOBaIS/iAnZlME/0I1aSI7A7kit
HAiw+f/S4js2o5/sD1wEV/UQ31Uw/NeL/b//9w6fNhwu0n+l/fJosGq9j5BQFxNFaSdV9SUMh4t1
YdLfH6vDkFFlz1c6dR1Eg5k3V2d9rocVmLHxQXOkOfYz2q4JKIiPKZqWR697Ni5E43tnyVq9SHhS
uULNibjB7Ot9hPUAVHp9vbrFq+rn5UcGiycyIyt2wOF+atLjWcV0IRIFiQcgOlLO9HHKXbAjTtKs
pl5DM0lg8PEI/Iufkzn1L1Y1CmO/adDNOyUwF/3R0AnQEUwU9nomB9JM290LoEKieHjjqv6+XTX+
rTGP8eT+oBeVzUZqGUxXm78o51+vp6lH7hgIb9UWlBR7EWpg8Ch7g8+ZrHisWYHwj1EVRUvVLRyd
Kol3P1/DTKNgIT4WZPRdn2vG+UYWTM3z/mSkPPcri7xBGU/Bs6LNdSxjaft9qwdh9g8qS96PauIY
rg0gdapCnuYej8dzRLX3EJsZGEjpLVItdiUTwEdj0FyLBs13Z4O+PT1/GP3x20s2sghV6vKJbgid
HOOXTWUqN2ODc4eiMd5+0tGcn0K9gmi+Qd6mnOYNne39/P9hjOIGFaG2vJV+pCmTLplE/y4n1LsA
Ep37qwWhf6dqDtmg98S9fxfR/XJNYw1e3tBZRaM/eiW3diVYtzAFh8f0fFLZSgxeRhAz94imxrRx
txFu91FhLkFdQjTh/QlAjdtFn/ccBCZdrmu1Nr1X7VG0oM2vzrBVh0fyfY5RXhGvJ8U2RbQwNEWY
NNWcKI72jl0dWg0tG9Oxa0VH4dN2UJfztMicEbjAraewOj23dKYnxYn8sVGlDNuXqEatWHRRGuY/
8O5674XKc+LifYd9OHjNbUu7X4bqFkVPAPRHfKUp0odc3jsE8fFFYfHdbqVxp5GVj+RHn1ryDN8h
q4PkLLK1mW/doh50XDUXDpyqFM4DFaU6j9wJA0h2SXHP00+xfbtQjV1l+K2kR8XiTjaEnR6iWEsN
XJria8IsvBm3/CViHi8nURWrsdORXY5jK332FwomV/OpK+u8aN3M0I6DVQyoFiOiZ4jFM13ZiPnh
cCkccVQ1QsU2QwjLK6frZFdb4/pscQs+SfX/gzkE+NLNmbe3BEdLvRPbQWJXJHie6EVqJFFByMlS
5LtYyw94/Ffup5ZOfbNaj9NV8EVw9HhkZwRjpz6PaFATq+KgGvNnXqOFUIX1/G3nQWBF4LUDR6bz
mGrOeGfV7RnKQcB9yDtBoV2D3xqepL6GHGBuC/+ATad9VI68ssebGx1NIsqOH28rQP9V8ATzdCf0
bfoXUhbPPBmfoZoj9mO309diTjVaZyqmNxhvgeARTYdTCfUMrVrWCah3TFyebWFBQqALXWcA4R2Y
1FVLNQNm1g+JfklqYSvxhM347tYghlWkxSpjMmzPNhEqV7b1YSEApXF4wFBp/wwgGjlQPU068YAn
I9LC/NBmmD65pYyfZUvNze+hzAw70248+SxTrHtUygv76+0m5IRM6YR0H0L3JM011PcTyCy+L535
qvnahWNTJiHMqRXa0pSxdnAhyS/u9sjQLj03fcGAMdbj9HTWGxul+BAPrcSyMYpWj4+SFRwR7pBp
LLLef8dDj4wdn+WtbzAHA5BI8WJ9mP5EtaGyW5huEnCClrTEWOV1aAH55aFy0O78QWL2LG7TtTTc
i93BTXAUP7YG0uFHIQceqBYs0VKu2PEyfVzBG7crdwnfd+WYhrktn4XL8Zgdj/FHZRa9YCOKzoml
OwKd2ChNPDTpelji8FuBFFkG3Wa9Y38Dq7k0K9u3skMmQHILjebnYxpwUXHK8bCYervE6txUROVr
xfFonrg9FDBc+GVkZhGhDoMCakjsP7R0NW1FeFQRkdChlpQ5gyqjf3RejPHh7hh1mQsG7aeJVHry
9HQfdLZ9c8ps0jeq2zT8b/WpAMyc3hWp3HX6hSQOfsNoyM6/DKJAxiLisQS/7Osdxb67cdvoEl48
09ZwqpzAiBrpZFKOTgmjjH18MkSV3zBrfqNDQt2E0EyH6/oQ7/H/A2hXrrs5AOEhs9F7HAEr/DK/
20AfR4QwK0mn0cjRJmznIYwVm3uJMtQWFRryeakKJoKo+JzKCJHpsFluuyqGrvwc4xVII8Zj4lWy
C9Wy3wQcJFL6uGm4slTxi6teLsdgRzRZqaNPR2R7OcHIh/DS5JFgwer1HBd/pm1uV+0siLL3PZJJ
Rc3eMRJnikIw2+hz3hn0LmlEUHmqueqXqNMLzVlLw+PQofZVdgmBdEmCRoo8r5O3AEPdLQUHMamr
VQzEKariUbMcTCKrVZSeTHolq1xjEx2h6KVne5MBqOdR5sii/8Ako3xICfjWqCdoQerT+rIDF4Fl
Q1Bx8ohm9VEMch8s6Sn97JR0jK8A9yFAvHYuuoHxdjcbvKEqiXENmpsvhlUUTn11I1ZxLZ3SJ4p+
s/ccyJ4hrMghvr8Z4P+zG1rDzQvScJPJ9EYsN2sTxgWxOREu9KUiQTi+HamgF5MQvm/MU6da/byN
C8g5VeqeO/9VG1YiNAS/OzphgRBIehoR2tvLG1LrInyGHiUkPZ4zxQMLAhhPfVft+Zqa6lKhj7Bs
ADKKJza+XIvH2pXCCovHNbx0qlA+Z4kcxku58iwNPeyFMKb+hJKcoohqt6sRFR3mTSDL6/Dh1TFI
J+XDun63MGCMQpp/nUPkAFQfVchpamTr4BYLn/OMWYJg+5sGm1DL0PALx1+/ag0Z5Dej928AS8I5
wOZcwxw8eb0wk0lY8KEKiv4FD2KqCp+FL/JuRVkxkJxWl4N+nSedQpGToIbSuKFDzL288p/bTZvE
6nN+g4X/UK8NdP+IdhNiO4DnD9Hv8EWp4vZJ9LwzzPtFPrhLtW5JaHLhhBoCm/HNXRl6+3n7zkdT
Z61vlnVKa42DpzGZGF1Zx15SOmGiUtitRPB5iG3Ef8kcC9pVVTvUaQWECus3qpuKetl3709Da2YR
r5GCEuCGI35243OuWCKEwOs7Gr3cUlJFC5h04Q3rYXEUIJsgD0YplQ8D2V91FWkBLXYLlY31Lv6Q
d7dJ9rcv+1/qCuC5QbNXLoX4liooX8As6GOoB9sapAZElnhSHcnk75Z+I4vNjTj5qRTOhrkUQsSo
HUdpcwJc6wM4Y2qruXKj83IHkd0qYV4lgUdbvKltYM/FjDaCnicm14EccfsWv1PF2hVSoZctU4Uw
hm5hqVqqNkr9kdGSJQwxoExgTrPA5wBQtoGCCVPFVRx4nqfjJY+EzLrXgzc5yOLTw1kKXi/QzffD
UBzl3UH1qOO2yT4E3ljc3jlRdssLzV7Y123J+IwCi3EaXcH6tthI4GsjEEYjDFyAL8jja5Tljcc2
+rjdFMwxyXG/RkR95HxHGY7gBBImGjzVf9ylERqD+52sGNUCH0E4jbf7N068nKm/iNtWYeqLTacg
QbsHaqW88Tu80Ergo7eArjZ8V2nouYQHNdyXHiXXTw1JEFkRRQYEiOeb+ysAUnVwdWCEMulHLEde
Ws21oslR4b2IfPHzHx/4SCVoW7tCftAZFEAysdV1oPCF8O3L/OXm+lzFOXCWdXrFbm5DQmTa1AmM
vmvRAz+Zj4AlgDZb+yZB18NgRFWQtw1AKSboWHUMdVAqJjP+eU6NFDmAlOldyIhpRqJ7zZn9V0l4
/f025SnctBWjZLw4RpzhWA9gf5S0cfXqWu3iKbXKA/H4ARIsLMdviLTKbjc9TD8uv4ep3AUqNN5D
yFZKWDmOrps5ik/G9WEYof2afPUBAHhNPHO0ea76iDhVWslQIpV9Rg379Paud32O4lGbjsq2xrk3
xy/gMQjLuPQV620lKGH+ZzHBi1XmcUJbah6WkD3jBZjWKMmGBkhfj71EyG47DNJBB/szhQxWh1av
ao+3nW/VwYyEr8UIXAOa3G06hzQuxEW9iZZ5c3tZsy7kXn74f6rYBHa7xoejmLCxAw43vCfmOttL
BwctqhwYr8iHnDVTJpZXksUt3UQ7AL2BqQ1IrdW+yPHuLp2i25TIICGEEHvcb+67HnTWy60Mk4Kn
UFaZgm6/i4svlWcUKWo/QpmwpYG6q0frGRP1SpvXtNzelfvEjLlG2tBKJg2/xosfb8f5IaKskLCK
28RuCxYKLDDZ0hD0O5E6qri4iOo4SlIccR7qr3uh1hXv7yLWmya1j7kO0JOALk+227iePW7AmGQS
klGQo6vDU39ByRvN8Kt77dXdrWZeegw8OOflVDh7PYlWCeGuqhJXgsJkyLWkoQDakq7DaILqwyo4
Bf5Q3Tq4tPydygFux6h4S2nqMbfmleVBKvussX3qRvta3ZRFrfP6aNmkqJNnBcEgr1VRJ/L8f9i5
nq52Dpv1GaIKPaiMn1rlGBYWEe5DYzU6Mj4R4GUgYVHy5+I25XVzI2US0yuNaDQ5qRcjNgtabQdj
8wN7Qe2UcIh6xd1i/1+bckRoDrE4a4qH8tLj+BOfyyGLJwQsGvV9V4dqMXCzzhSmnPha7hK6NSsS
I6NlmgNXsaKgpwT/eMOA+yPkbVkUYHI/mMkfQYqVuLKLHtxaAHLyx0wOX5KjSstTmKUkv/kRY2JS
HgxA3niQLvucCudN8I9GBPPXQufKKAMhIkSAN01MGfshCXxZPgEP1RXMUEfwAF3EszYzw0cXZHbJ
U7nSxk2QPeFBYb2qv5idqLjA804U1HmuXQLEQg9tmnmjGXdBLdcUNpSSNFxP3MrIBnEjvlnf9Hzq
LMXrXyn5vkvnsb8jZXigdHM4hORadN24bi+6seYHYWnAIFpbXMWkI3MBzCvYZbWbCIVGUjiFRGdG
nHugdlDtAlN1Nn4WrVbL3TNJPZ6fszA4hC/KROxbuGtqGCT1q5y0YD7Yr6kj/1c6QNP+SD7NyySB
JBwu8+lWuzHK89nYX2Pd/2ztdgrKGS7a49FV0HT6z0L+VjVLpz2yNGNxFlAuY6kW1Xe1rapqPWgX
grqa+8VEmUUE9YWn8CgsT6ecCw1sG6Q5DB0nxVS+UPklrdtGilP7f8cXSgdYOZU9MsDO0zblhZiU
R8WWfrcZSuJ1hCADRsijuR3/7Xjx9BWujS41P3LV6GPu1ogFA6zllKd6fKHbclN59u6SVfm0rMI0
tOK3NEufo5meGzj7fY0lfpQyuRGaoHu+t/Sz+yPO3551SsJ5y5q11M1P0cUAIg/nH6jheC+3pqHU
9EaRoN93fXytAtsBAGwjfX1s+E17hXbs5npbebby7tvIxBkFaVtAk3DTctlhbNHG7dAWxugrJWo1
HcETN8jJ2OQsX3gcXUjEaeuPqcBFi2eJ7Je6tAgRF3+BdRXk2kCKKq7nw0b7kuQO07vQ8KwyiJrs
B1/9rVooA8kVtqvIQTGkE3yH8NuewKmcaB0N9h1bYhJirLF1viy1UbJPBQUJx7ieqhy2DuI62HdB
LeT/9WkQPFgoCF9v+zqKLy21uVsdH+Cb3GYzmN0AtSbVD0MlG7XZOhK5WXltPeTfP1K3ZnyIcUbv
g5hYWVNB4ZupwfmqW4bn3zXehz3G+dFSiYVJuyW96KRBHLEKis3VBSOnFGufhTtm1bin6B5o4j19
9SJn7MZpmbVl3PQ7gM2MKByKKKfVlSS0xO+/Vp5pF9YPy8IS0OzT4SDFdFzjeor5fGRhkGwFzXR1
SviQLIW+M/jn1NdkqghmnyqzzsmO3okPr8vo3IcqfIQ6cPNZIRSE8WuygpSSW51Xds60PcjG+3XW
iXb3yPKciW0IBwDCSOPdXCn9r7Xm7b6uUOQHxpwciaKgRUqKSxH4C2eWVGdbUFh2aEjtglrQUwjp
kCrHymjLuRpTkckfHdKrnvKTFMgok3DFqx/NtGBSDFPd73l8LMjQwCa1LvbqjF4cX3BABG7wcWQh
TndvEy9pFJAecdjwpAvfWVnoqa/zEcVrYdCDmSkFe17NvdRyjswLuHceEldHUbjqZXo3MdQ4MOg6
oJgoQLIql05dyb88fhmPv4zmPuWTEbGqRQhj6v3a+LOJg+yxydKGYAOUSyHhcK7gA5xeketJdTe8
wSO0PZI8HY891y4Rdcj0bLhRx1U75VoubPt1Hx6tRF4KXJx1DoxYRWkUiufIs/9X3oRW9AtGifaw
oLxtvezLoFgJVBUoCisFQXYO0ttHMYt3xA4Tpp6zFi+c4kZ3tnchfOiCsIAmhECCNNOqDI5j5fGO
MB3eTl6MVPDZhK4yeLUqOyKL1goLcbQcziEfRbnYqr8RFR1Rr21NgdCp/MOsj5Qlib8Cz6RtgizT
LYA+f6uX8fzQiGc0Z96ICo3M/ctBfeqnRauzmTrZE64srifX4mrDWBl1w58suS4slc73Xpf6JkW8
HXFEh84EJ/tWtIKhG0jcesHUYd8pxcxAjFyPCHNDZAn7kobSyZfjlk/PQ1vkIlQuoS42jEg25zxv
6L78ewGySL11PFt/PseVZlkiwUIzFHg8ee0VLaKhw63NBUCEcokkAYFwMzCfohQqADfhxZytYori
Ix4/sw1rz58rmpbLW+tdQLDb+D3eh+JJUAtCmfaA/cd3WFjIT9JDFDxSlqTmy8hi8dcMC3e3JSiX
ijsvrQ3MvRZIyigeP2q78+jKHjgFOCMGFsRY/N07sPMtzfxmqKQriUhEW1OTfKqE6YHcluUb0S56
dEhFm0qDJ0H/ANTcEU4WJAre5W60cJrE83z/qhRq6pQG+CdrI0GFpvLszsmUM+ch+XFImWG4egtV
GL2VXgubv5aJRQXPOYbWzKej3YrXQqp8eJuQHKC8M4AjFKERl17YQ/hYH8Qj4T0Kxi42bbdFn0W5
4Adqo0o1dP7nX5l8oYGQIVlVfBXbieTFOskm4EqcNOlUNsdh+BqTtf1dEcWP8wMkBQTqiSWMPMVJ
6kt/zHHJNm8lrjr1h/gUGZ1FsjrZ9CdJhoI5TQ1r/noXQx8HSFagsFYsfLCuvGsqoQRQnAAmwqkx
39hjf9XS3bmfqAepJeatH9uIxhFqDXkVbun0fnNm9J6MpjVqSGmIfPOiupSDUE5OrstcPm8gfCUf
8WzSaLmgC6xs87uMwjyMqo8NP6jEzmhUhCYcaHRGVKN7CiaERZTIK2D24XlVwc45LXUrEfqEdsdV
XQnEA1oZLmZezAQaMaLo1GtQQ67LaENSLqOQLbhcxfVvb1/3avw0a4BxvYZ88Iwraw0jEhN7X4/9
lpwp5Hfsm3/Sj2Z8bn1NQJYx5uyJswSW/7nPCa7OmDGYCM50NIjq4+81iV4L5x9IGU0JWc1Gk+m9
61ZpXDHq9odZPwgUVkfc8Lu+UYjJQnZ6EqLxzjCXXQox3EKx7VEWhZF3ZtFFGfFN+hf6hPjAEIuv
R1lKync4ECWcwBJ7H0hsqXZpspi3uIzUevNYTCuW0R6C0QSpthlTxEI0SikTCERNrpCifMLlEv3D
gE1CEbPFkyu9HnNHRKH1t7lQqbSNBiV8kxpK/vSfR/7UauzqtmQBAosjDnGYW42IU8u1GnG5G+Us
pZKgJiDvth183WtXrGapxWcy7SDB4RdW5LbgP1KVGTy/FvOchiU6P/idNonmqaIyrgP9CfegRSjV
bjOCDK51lGgylDlEsumM50YjUFY4St89OcaFkXBW9FZ7dvJIK+9M7K8WLpzKyLZcYaJqvskuAoUO
6Nof5H1PNx5XymvYTOpgmji8jGzD0zoEiIZSzhkpHLUl02jxtiUrOuyEDL6MmN/GqaYSkSGcooke
GCtUbFsTJWFvbDneA2Izl137aNxqa0XGJ6DkxRVxnxykWyOc88Ucd0y13geEm86yICC/INqaAPBM
cT+rb4hZtYB5FRvW/zBi5UadGyMjO8nhJKLi3cn2MfeGB5VecOWuBEfxIWs80ZGqHrHVzpCkIfEM
vDXL3LX8g3dcv9TZ1KM+budu3+9SpDgdpNNmwKdUym15f5NkBnKrdUnQwxIQwqzVFjWeCHroPkg6
cyw+EwLGYAfc8hw4Pkbu7F4sbxzE9Aw/+UVs26c7cJa+8Az9ImSUf+HmAh1SghhtgbglnhcPGq1Z
dqeYsiT1q/IsQHG4FpYdlJCdT6M0/nTTEt8/pb7riCJwQCB2l1ZQU8i9Ioqd8Xa+VPEyxqgUz+mU
jRnRuuiO6d+cooHhlyRFQdSt2qdxhAXKGW1bGXLtcKh2n4fkbcdTGRYgo01KeqhCNGU18DHFbid8
eKlO82fJuU2KzzcGNQ6cG/3XiNO88KimaeJGETAp2DiWUcvrCiTg0gyG/A/Ny+LLQl2kx0fc/X+P
YOglrFlElWZj+KFc6d+vjZrTZ9AnB/JVJtEJp2E+WIwWwsGqQNLsixUSlI0GthiZKRYVy27zRPRt
gS925xgZPmjRhXA3imtAibrVO+QpBZKqHGGM/GTtiPybyXIp0WgDCbejAaL3R+PfBNLw/Fq/hmld
1ePv9Xj9X950OA1Mk/+Cvnzt7eLQHC+GesKtmXl9pK5D+Z0C67Tk5uQAco8lHXATb2GbQ7IR
`protect end_protected
