`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kK7s+W51Sf3iq9Q14zoVxoT5XitQfWjtZzXz9PblaZjxgexCPHxwPdN8HyM4p7I+ZY6YQRtiD3V3
pJ8bg/euGQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eGAXZWuEzASqV3f81RuRUZism2ELJ1gUKQIApixFPS5Pozo26X8r0d0wr9Su9IaVSlmrLQMl5DF8
xVSdYMgQQHOhHnA9pYC937Qm/YApUSXRPAFU1cSQOqdP5acZlwqwcqp582kufpEuNduusKvdWbPf
EfijnIlZB/Wn0LrSEAM=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TxQYZsMixNq7plTbwecaz8p3ipXwLcPnaERyPvxHpTt35epWsvXlyeVzPkCTulyLsC5ouYastNGP
q/v+htfVjCHhGYhzj5m0zcedzXAb3XPZNtjSvb3/DIGt12BUSjtoSFnN1gw+Nh+3q+JtVDhE43XI
z1M7R/ZAY3+GGRnU+8Y=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VpN10r5VKnPnzN4Wt6g8e5a6Yn+zCb782KRzvAUrrQ84xth9xf5B/QEll++0n+jYz30moLtdM2xX
xXHlu9csdMLIFy9VInIKye9HgdqPdgheWwr3m9sqNTNIhfLZ9ZzjpNyPN5vDZGZNEESeCOeouKq+
8cffxIvK28R8y92YxFJmN+3Zw4SHxiUCGUpi4qx6m8EQNCDqDhIMam4gyHfxnI1MRrNwHFeG54lM
l5NExfTN8LHyiCUzKkM6JwRsU6Az/4E5mlKofnsEaedEgFfrXuI95F/XB1jeQGgR8QBXKt4OMObm
9S6H5pgSsnETnIeASxJjWQ1q9zEXcUnY4mwwmw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nN4362U/mRmXW93fQoq2uujCxL5388DFI7YHxYSex+C3AkfzvyHAXovxv/+NdYUq8pWO4uWY9ui3
6vxRgMT9nl7RM4qZkuXinfv8mfX6ro2hvmHexVRQpTfGbd6gF8iAA1iPzv6oE07JcCNgqlPPBI2W
h3bjfG08dDELy5cxS7l10LY8Jj4eM77Elcx8fK4vrQGGEyRxghTap0MvM81OBLYV44vhZtW/QNa0
e04aG+qajlp6nyhF2hI7cB3DaA7LsDbiZJiVrtxB2pyKUU1qEtowtkQGhqI5m5Ot142VN6aBDHHN
MOn5gryzNAlSsI97lTNkvnPkBk/f/mTKK+XJ2g==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DW0FWZLg024UjPuExIjYPRs/W+gp5pfWg/6rCtkSbFjzaNMzwTkn1a5mgMTB+Lyo1Uoa+DRHt0lc
3oMcoy8rfI24MW3t/+h/YZmGvVILxNreLtUevUsF2EtUv4dmfwhlcoCk7+OGkQC/bgv21GXFf+y1
sdTTUWAji4yFbvpuDFhQak2k3SL2E+ve2ec5nKqHgIGDUz0xQNqogiZZLL5lDmfUlqhmo/stTCP1
EmOzqFvLVHJl/NTQYmdl7PQ9lYCDyIt0XkwhnJrPHPoyu6ugT01vxemr3cGBxFkqgcjfAjRIy/qn
YBjM8LfAOoMFWvSuLuVmsbMuH37ksxD6kewCtQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 779472)
`protect data_block
gsdi5KvPfYEPKuqIsaqhTn5pZA6awZMTtnsi1wyL0AoA24/cABtTiV6UE/LU98oFLe8M0Q+RY5FI
D6iStY4heGa9+vLGfvy6izJLLentgBFbp81l1Y/eCUKWmgoU+PEpp6cjKan1Crmuel6YbZoMTF8q
2nx9MY+xyI2urUAYa79Sic0soPJIC8zApVMTZCHnT6JtzIjtJfFlMDWm1yS/S5fYPjPU5rThcI6w
wYo/I0TVRxmHops15l7ilDu+85z7QEmfoSEypI04khNa9q5a8l8eV8MOCnoRwlBj6k8P16n0inAT
cOZCUIjGWxiyb4YMLtfMZORYTGPFmgpOCgwM3jE71N1Ysrk23sqdSk0KQaUDFN50/csXbTjsxUz/
+uwE5Mi4JR5nu8nb57SYviN7B063Z84a7l3IzBq6zR4oamu2L3QvKzpcuQJ9HFyHkVYRN00/op1s
7fNgqh48/RneiA7i+HC1tAUI3FfIrpx9DnKSDBrFYncU4qdoHMzLMxmeejKBZmjK2uHck9uurs5N
knuxhEmOWkfj/Y51KAXtuCAgJnv8k5F0iUzAl98A+AQfLN2JiOAnehFzdTjo1HdKFml9EyU1++8g
9ZuMlzQ9vHk/wlMLE1+v7tjc3gDubHxghO0LazPFq0aoDGZxKcPtBE0pewjk8WHreT9p0dDQqeOn
WBQDjj4UzqTbVuI4blWmaeAtwoLnjPyGy9BmJxI+Cc4sdAMK9LWJRaZkQseNX8+iXHh8rPoOKB5x
yQx6dt3/5NfxvU6s1D7/8FbSQLQl+9OvfF+2XfIjdfmFVAPoa5Vu2TG4GwSB0u/uzJipiPi9hB9h
V1trlEL2AXY9velHaYZUgIFLNO1eS3etfInhIj4dJ58Ii1QNzqvSpa/xm+7lSH4oYF+fKhKgSu0R
W44b/Xlu8Wzc6t6B75DPu8zxA2nFGQ+SoqCuIE8yunxfLvBErovTy82tMmDaRY8Nxv8bessoN54l
UbMGAO0dJ/yK110p0CFqYHiofUzUUSxOkKblukdpC4xkltW75GSfDWNSwFsgk99Y9s7tHusD5z9w
0GCfxkccFjUWcUeJ6phFSzoQ39MH6sxbsDhddLVGMj8/5C6np72b7NaecxC80WyWml7E3/LEtte4
TCyPNI0L5ITaEasu4SM/P85ssySguiyc6EBH1AEWSRrzuWbaCEVOwj1Ke0sFQM2BFl7NCrlvcJTo
227drUl9LJC/m/Vctls+PK4ef2/MKhxDegQLCs47tGt1N7MpfXt92XmSR5z7EiNHcW+4XVh91Alz
gGBI6l5bYyhAcKktbKIranCvR+INO89UINGgWutjeA9qYobmK6XH7qHpQ+wIXbekgX9jMYsNJkd8
tG7mafXfUwRINFLCHN+cR/at/oFrXZZxc4uwcg3bkqMz9LxRvmbTfs0RryeS2PEL6TJFCldJKMSR
2TF+WWArzb+cuo61wiyeuOAHjov+c3Tj/tl94vxp6zmP6totAXX+RwNegkzUGN6rue2UISMKN2Tr
HXdSAKnn0Zl/+R4FFDy7I7enoa372WTlXk/1qkS/vGbFGoLjt98uEdWVVks19fYv7Uh+JCv7y5dP
Z8N+if0lKpF6NuDzBq6hkd4jjqLwh0kGWOhNb7tRGGmZVS0VJxmSkL6aXJRQyGEZrLT9gOrYPNJu
hUP+3YapWVpJSXRieHFC3u76xrWmXoGPWswmR/ZZ2XUCNCFiiL+7dY9V+P73QKox38z/TlnZ13h8
v5523ka0PN1QgC3CbVxFp5cX772jDt8jdYjjKqcycqyoU3ADRuMhR7OeG0WZW2nomfXV1guErw3W
hyNsZEpP9dUUt/DSH869+6uY8Mmu6cB7dy2ETcAy3SYIaYIfGiueJDubmyDJEFOzBoY44nrgLUja
XDhK9IRHhMUyA5Vr9LtQguQd9WMzUxty1LL0kbTT6E58dHkhUVsExIsO5fljPQzboyyQJU+fnNmk
0TP9JgN00glumUAA3uqHaFzZ4ifRKsMxzuSJ1Q3JcN9b2p1d4EOz4Qr360IpfQ8SBSG2XwsryCMA
6NUF7+ZAT6otsZglBW6l1bott4aqZT6wNJ55cTspgJkpCEaPdOEfZd+mRJW3kezDXzKYNGXUKsYt
JzHUAyS3sIHK+ACkZmnTM4K5DbreVmgH30tZZsTttWeYi4mmRgD/yJCY0jjrqvNg1+GTF/ANR5tB
U7r5NSOmGMalTInoJMUGlTBx+gRP3X2W2vGAoRggKq6YtcJUZ7ygN0q4hdWaY+T+aJpbew/vjAfp
LnJ6DnYS9Rje5ch/MYnwmcdYJigPAx5lda8PLTihDo9AaGqflVaxW8So3pGE9VgxIDzUanMHWHv9
eA5QxWliPyME6JfOWKZOJl/CKBUG9DaSAWCqcq1dMrHKBHciIkWQWGeadRgOzgFULRtBcPMKAfVN
QjeCslqS4FIAJb07+X+k1W687mqDErvwKaOlt83aN1ZT6dVbmLPHS7FrdwGQwKEPKuETLijDCBBc
BFfBHATLq4jjIKI4MQ43CZ++l6mLSkrULfG1cLtQDoO7/3zAxf0pX6WnHV1v3kUMem0SQqqjkxjs
ql8HK88RwKKLbewrEjRn5DdK7ii7oKa5VJ6Ub+8D8sQWTCkYpeRfKNuCCjltNDS4272YqFVg6wCc
tF2nT52rpLo6bxMkylOpqDpF/m8Jy21IiogRtVRy7AJXg7ejQX6sdabs533/Qd0CdTVWHoElUQZT
MfKzyETaRPCcMvdh7izQI+QmL1ULl9wkhaXO40rRdO1Y1dXWSUxh0uE28rCEEf8YT8PtnL0oEISg
J+YALU3MvTXkCxhuZQvPA0rvEAS52d9ilPAcHvwTv9RMdPGER4HL/sgHGMyhscusDLhSuVUyLVUh
uw5cqQJkBB1vFpCwa6i4SCJ3RfXkBsPZQ5PqwYnoNK+EA4nwHw/kVHN6WnEpBXfPKMR5Gxbj3kMG
Ghc0uXdoeXyB/K0rvN61Rp+BCu7yCo5ut8CKsjWvY74ZB3ux4xNF2RS1ec8Q+GHw+sb2OHrNGamr
RXucOuZSYC4ELoo2Mlk3Wp73z2erlK9B1FkZ1V/Jp9bKL0ln1EEkbX1CeF8Yr1tXzpPFIC4sNwmZ
XoKvXDbiqYmh1iD2I2L3HlYgLbf2vRkHSRRglkyJAxl11JCw3Wju68ZFtLaM6S0ba20hIhmDM+1X
FBW6uU61AbDjtpCMHQkbibZUYYAHRw4UCWEi9xT5hU1PKr0L7gKt6k/WrNMCbZFCwubBDLol0DjL
xKok0hNwmnrK/V1snIIypfb8y4/S9I5bCTLGh/fP3NNTCyy+6vfJM1KgzE+kg3GIuQ6zfc2z3tZc
9ac8dBWul617DcRQyO7LjyBcdkPSgtgRO0Wjy6XaHIvEOZO7IR5rfsE7/8EV0NU0Qx7c1eXZ5MMc
iaIZvReY2VtTSdGpXchsrR0BAtYfbCiqo7gIomUNAHLYN5f6QTwl+A3+4xYKHpyQBET7hr9tRNOI
n8b6wiyGKOtKTvA0uTBk/lY5J7PDGGQ/++4Ue77A42y1Zs6sIjBuI1X/1OVtsBv2Q/vlZurir1Vq
DEt7CRnc0YB+5EGsagrDGUcRgLpCgMSqNbaNctA9IJjweUjcf66KhiOg8YKdHWUFMMapS7IOCWye
XghAJ+NKYGr2gBSZp/gKJ+XhqoSfOWV32sbJ5LDzQHcU3yK/eLbWg6FLKefxllm507+empSWZxpp
0t3D6pIJtYF59NsSfgnT11ZDN0eECLkoa3vmgWnuI3zU89YmJeUpYdvGntN/tpvV1sVw3pYFBYB9
9Ph1xqdQDevzmqCf4UX+bcli6VB1U3gV44l7ziQjEtq2WHMt9ay5G/isKh1XfwfTMwvyNJxejWHp
yuL4iPjQE5WF+jUatbLnVjljZJ0tkLrtU2mUTPndfaDa0jfgjbKACCTz91JnLyAIJw6QpV0TrYuH
YJNxvJIZIv0e4TC4qJwLeC6XiURFHKgOso09evmKDV/S7HE3qvjYj3/yjp89QdpHUlTd7hGaZ0kV
2OZThVc8mob6U71vWvkB124DdIZjRBGvn2nxe/Rq+gu7+mPm9QH56DRhPabSe41KqQtgenSUn86m
FVzKAJFNAPc4WUlm6JR2n31cAuFvbKfYYDk1fHLfnka2yKnbh6F8n9NypZxPNdhXpGYYnfwZ/vNi
FeQ8o0ANqZA/nXGXDMmIwtbPbI4fmJjleIPAiy8kRlbZxLVzEqZH1lbC4GLLxQ+bD1VVBb0ykie+
Bph8nZ2xyUYKoShI4sO2bWdirIlae5qJiEekDBrH5rOTN3EOZZAH8S/BabdUaz4rDRJ1ySBqawug
cyPb5IwhlNinQgKjaHUPp2ECKuib46NrWCqAbA64QYfR9KEs/fN3VxkxV8LeJqnbSCosouI6Fxzx
8gFdpjqfH5jBbfpSJzTITuHYFhSKlBcYuZF7w5kXxpq3bdDM0Sy8I6oGRXLzMXoh227mj1xLB9M8
1++qCaT0MeKwtVaGY9iFfPt9XwStCGztXL66+v9rt8qglBimXsva+zu4v1yUfXLsfP0tMeLpHsi3
TJ7HjJtGOh8CkR2i7nHsDDieqNvZ9d0I+4IwzeR1TTwhdRfiXaQFXgI8q+UDv1YjA3QGJ5osZSOZ
F+Gz8vh6LkZRXhF4HBg9IBXBwi9Ftpq/r9dzt+QPHdwUkPpI9pzEfs26a1BhQl9yAvyup7rPF8l7
NnBvlUX6TaqKepTQ1aVxZfrgAEus3Vo9GaNAne5ornHx+2VUefsa/JYRptkdvzWmRRaSNzzYhh1l
fbezVYZKEcrHNbc6P5EycgQbX3o/lf85J1VVRI+DZMhSMXyGeAwyu3bffb+yitJUgqrrylwHBn0l
n+psB3SSuj7/i+J2tH9kRnMKO6oZD3E753N0HSjirksCteDkrRZYQaiL/YW2ZdU1eWIDRzaDe7tO
7HKi0JsbyBa7ZBE8rMcPOqYHOykakYix3YnnNYqrek/IPN9r8MIucsCVZsuevwpHFa6jNmlrCIc7
bB+zMHslLuAPK4cI9bZR5C+02N/TohTLtB9vdjSV+fHNXOiEZzAP0nBcQY6LLsKqq7KcqkgjU9mn
+Wt4rzrjV8VejwZJDlv2GSYZIWexX8q5qYDS2ElBE2gA0IYC/8quNVODT0XsrMt23GHk1XzFUkrh
vAciGGn9J+O4xNSTgTI66aU/5fGAfB86UDc/gPHep054xaDFyY1ufMRmrx2EAu1MYHVgsqJh3bra
j9pAvROowXQKbT25QXTtdjvDW36fzpc0+hr98zMW9HsQBa1vTAb8DYaGlZzAvPVrhCWVpwUfs1Jc
16d5A8oMv4Oy4lXrcKcSEhrnpczDHzFzxUSXdDEhYyV2RSOLg5rOlKNliqifUuulLydrE5E4mFc8
7Cv22lkwi29qv0+OQp539Njt8lZ/3XnUKa0qK46HuXpLkjs/3ujZzeSO5os0QxTUEXDVycGQ9IYh
JyxioWpf4YSTQK+ncbvndmyl6c3/AAWjVnSRpiDuODh0emoTEIU0q9M3C2OH0u1Ar3rP2fYgRNLq
SZIHJmHgUSEk39HC/8SaqMe3l0XwGHKJJOGvnlREUzfFv9DC5S4Q24mRdT9NR516LyIug7bpH6jb
EaOjXTtddxQoLWlSG7pR6E5Z3AEZ+rBgopo0yn1c9v8idZOqqveNTXFifDsVszy3u5TPzlX2E78Q
2+yL2HHvttmT6eemDtsleofgJBlPNLOI11TnzeEgowxvKYXfeeAAGmmeChZweZx9ybdnFGxbYuXg
XArwVhX2ngqnaS4TyaR5k10LHDOBVkm2Ghx9p6j4ypEAMkR6z71rBP3C33EG+xvjuNyH7TkpneJR
QZ5LAQ3MGFu03zDBMBdMFv+wcBpuPbe8mjmFycglKjHec0oR5+PVlw0zaocw0i/95WEFQEQG2CfJ
lNeKrPCuDkiEfbS3j1LJ90BSAwln2AlvR3bnT1kNCUYpaaHQWd0B5unNlaoWZByKznC8btPKEfAw
Co7slozKTLmoHJWluzfneMIsDtuM2px6nTwSYRlwrH/H3yHLryKhERcrp14kwFfKsY4i+l+zBz1F
I8txGR54RMPvcM5SYJ2VnqF4ll/BtbopPamE9bXHSoD0rOpNPZ97VaIEJEWPBdb1GesXbenDSzUq
ReQxrvQ4dSDpc2YJbJs7UkzTDOixFUrv4u9ALpT/9bhhrl0XXJd1yohgcJPKNH/WmTQXN7dxLp8B
0Y3RZFxPgWsTjPuARDpFNx2FV/REJjFw0yV6YSbzLgvIrkMuXkNoHt/o6+dOPHIQ/RMI0BHGTJ8k
icssiXhpSOSlbaW8ztQCHmtO57HXERKywt23NWMTBIJqOtq0AlzVwvXhEwP/rmnX2p/kgZi/WKpS
TfP7GDumKI6XjEZ4zTxB8ShPqC7DbV19M8xNaKotgySxAw/C0e1zAtj7YQNE69ERLgkas6hnt2hn
h8oRmnVwRTynRtrd12GofFLAhAAUPm4OrhGrjmpxImvf+EOaJddAruKi1pPW3Fd0QhNq2C0TbjMn
/BWIWZMsPHijp5qmg5mZS/UQ0ChDIA1RAUWfXlBhlq7en6GQxonLnokvmQ7xjoCkf5TGPx3kmsYD
NdXG6kIW5gJuyvznsVIHD3Gtb2v8ioz6jHw97TcD9saJM1FRoqZVlJFZAsKRyr4G0iCKBuqClmh2
3kgCfTWE3LHkaN2xnHC2JRgM0NMpvviuqg8WKkH9mRymWkUurOpvmP2/GO3oeI+c5xcfUBrdtGj9
Ud8E8eKnBFsNdJTk8fMRMlmjF9dnsq0MxTwbrl7AC/Vs04Ns24sy+yRz3jj2QNjI2+/rJoRAziWe
A1AOzV58RVvaOf2u+NAVl+tZw/h4qEvMUqXQ2t47KltOlzqkBM1SeuP2AnuixJZ9Dr6IvN87r6tX
Y627nwmEzRAFFSd3cYgdKJm0RRgudEVZLJzAuAZB3DtKQtsQGdPTR6LHGGE9rIMPI/UGYUuO54FN
RiAyKk2QvsvyueI3xG2ib7Ra5e61Akliu5EaYIDy36jJNuOeWwz0DJms1Iae6pR3Wqojbie986tD
CJuN2nJM1QMMd3zNQ0YqOnM9w6cFdCCYkRWSBmqPPgzu4eN/+05FkAVqaz9GImmYw/WRNkRnvAaQ
osMrM5LmDsVYZAQKGn/ZN8hGzQ1RTTDtlM3cJ7Pz+Dtn1RaD0V47zSr2c6yiSgnQpupt+FqSQLRW
WOkgKgVkVm/WaAY8dXEHyOV/l6ybJux7estwvzDCb8uk263vAZmRiuwnYyiZ18KP+tT4tZf3DHpF
P0afDY++NAZeObARk1uDc2M45Wwqp6WBWCzmtr9gHolZl3bm9bswqjYrGAhgZUwfN6JjIWRq7rq4
B8zB7fu3XrS8SYu/OQjmiZbqgIFj68b58NqXFdc6t0vzYzIzKhep89eRSIOsze3kOPWFB7L5m1Yg
8+ZP8WAz8PpktlKus1lWbp7ruTuZe1F8a+4U/K8H7AVZ9HXtWzcLHMypX1wEAfsyDbBO7krk8x+W
Rv/NfD74522YK1YXTjFfzMl3JPKJD7CohyIdSrz08dqqSYxaZ2LjNAzbDcLEKOidTj6AAvqgq4yZ
hJDV53Csp3R8cMXeyE+2OBo+Z+TUTx4z9bHLBV5AxUSlcXAKoFSYCvRpT7TH62hQtaf9QNqs7z+4
Ta1xz2pecRtnenBPoL0fLIhjlRnV3lV6NfxkJOnEfy4Asdm3U51bpbUuS6G5zfaxXGMZJkNYU7xS
/Cl9qwzNU0HRLS+OKTTHxiJNNIdbwcFv9tStWeOHUYmNJEkXdcb1uMSN/UZpRKwDc6FFmSVSuxAm
hfTcD58lYZ6Q3SyqLiRn7kerkTEUkKOeCvFYxmlBaCS2v2X5IFdl/mUCoSyYJ5T+PqiUMcDXZ7Jo
JiMNIqraD02Avo4nmcKlF3dF03JZV3hggrZb8wsylP1vcupuGDaF+LKd7zXhuDX0RkBT9mJAzOaM
i3CEhFEKkeBFHyj9nkamb6KLYqmFIP8Y5ame6db6vXfXwbUBproBgwH7hbUtqcSjQlhbrwEFQ/Qj
4ZjI/jmJy3lxf3aCVk1W6hjV4cGGl+KB3e0cwez55W4KQ/pQHfhOfdKc/elJGIK4Y8XPfa2TUKpZ
4UnFA4QWJCUQkX8JdcZGsWNkiZp0gCn3mxLN2y7yRdaCrGiZDNz1hvmcgYjB4a6WIugSW3fikJ72
MdY8s1SrpcduzcQZ6S5WWUL3HGBdGXjFC3mXe69GKiSNFEYpsAizL7u2OJW4U4Rmi7MmjgXzLsgA
sJUZYR98+Os22KqSmJAyBv89azPLc5gOR/TaGDbVt/X2pU+6j23z7GZeFaXbQG3lAReaMT5WksGu
JUn4SmdJX7KMxX1wpwt7JruwcmYq4cBFE/pZ+TE8/LfEUU0ukx1lyrRfrcHK9DtVQL7RlfT+rhWD
1jHg/8GIO38yy2aQ2QsTtG5g+qNiFuqxYyzoozVBJfnGuBzd7TrfUY7iGNY1urBtN3LBXjxltT5g
hINfPKog8y/PvDYFa4Xk90BEiqLGMJO9VZhSVRpo2TeVxvIwoHkZpc8dg+fRrHiPNA+cEeZBFCFA
XLe8+znu7y48I0jA76XfLq44HpSS3gMUCNybOqgHECL/5PINtrjz/anfgnawfkWP8eLeFF6jhP5S
Ftve6sPdgOxaUeP5A6q0xxFm88IFztlP6Yj3LcMoUqYWMQVCJ8Kt451pinKlt4ONr29hXfIf7U9C
t2Xu9QDGPiyJ8NuWRut92r/7IF9Q4jTuKdIWmDda8NikbgOO1WpAcUhlb6NbVaydirv60JqiLC/d
W0Tu2SaH5vUuiql7aeUlcZJzzj4NG9l/cN7rvg8Htx5EW/pVpYwg86QD/Ba7JXcAnVKTgWzIIrS4
HWJ840QundsoLlFpauLVqVwb43oxYDVqnbrRqF3qLKLy8Ji0JwIJdkVjvIfVRbXKxWJsy0lO+72z
SkDMzWsQsFAEpWLkFmCbbdoZRQ7oddTsuI2rhDEnYR5q4Yol3tutHDa4iRQMWu7ccDajWyr1sIVz
iAFmIGIwYD5FCFiH8aJ1+kuHe2bMxSLA+b9M1O1ZPvggpnKfzyh3AgfUuDxE6a8ggGs5SVY76cX6
Uw8FceJbmB7IPFXXRbjIDp/mwzel8q6M4+CvILQ/Q4+BMWTI2ozc+67JrdhYkjB/kYaUSafgAo4D
NVx8BR8BGaEGA6IgoedzVTaN4+1WYIkKcvFzlm6VXu794Ub0aj+GzP0hktGGTfbF+++XAfxcGFzz
rNAorcW7N8Yyey93VTNmTnHOIkfiuecEG74uUQvZ/IiUZ9Fldy6hE7NP+ryWrg0PRG1dCk/h2uIJ
l8982/vY0pYYtBgjn3Y/8hHaEeslN62x6SSBLNK/GjrfcaXSfLd9bwnAgfpZNNtGpL90BVK90aNB
KqzLpNLYXQ++nfe7UMSUjeXQCq1R2KAkbrQvUzIZh+LGsRSiyNyn+jcF9tmy7bxHTDnflxEpv8tL
zpL2+hjPQZ2l/JG9SNYzXDhhjjTdf79S8hH1EKfVXfSC5k+i71qSY9P7/x1pimT6nHWwD5X6HALY
+W9nR2KRzsuTlM08cupWWyNp/tzVvurH1CrvZnCOwOfAeCxFIWz4rUcQsNHRqfughYjv78WvZoQA
RwtLmot2qCyXfri64oo8RWI1+GVsq/VQh9AgZv14ouy37tzfuzMc9eD9Xmljrc1rgdM9TSf4Xk3g
i9ktIgMTtaX5MUfCySAVw0J2JKwfaSblB+rXoMd6QrTeztcLca8p9ivTQDfYUz006t4vj/tE1SoQ
BKxkTPLJ+jr0Ct+n0W6peVnG4rBccVnjFuzpkUw2BjSSXYM8yFVy/h98lsZHGwXxVVikHks5fXg7
3kl37yqY2k8+yZHWarPAttRCpol4P1/kUs6EQS3Vo8EyKRrDQKs1vSNxv2fInmlb6r5k2K5iWpiN
MhwQ60HgAHL7spbaY8fB4hkbeUw1zMaYFmGAJpiY9eVrqYHsUKIwrFW3aJ/EqXrIYP8YIBBq/jHI
A6IDSiv/F5tgUTUvs1RRjtHtdTonenJV1O5SrLrE2G41PSOUPHlfau6ndy8Rr1faOCNVml97IEya
kyVFAT2hO0AT9b7NcktK+D1+s6Kmnn/IcK+CIW9DpStDbyWaUtI/KUoS0yuaG+3P/Nfwtf7RLjF5
Kt/5eJ5l99aWdPZJpmjR6DE30CXyNMP/iVjtJPzDYEf9amr/OSfHNIMwihIEJy2uPxDAnqysiuPs
uK2EH5UVnLd6tqOslJhX4O/mTL0a4ZV7N/TwG6ZxPrz8fg30p2tYwv7QKb83aQUCzcKXF4T4qo+A
aRo6UutcClrlSwkxM254EoX4Y0TOoE18Oi/Rby2aExh2Qr/1Jz3mg+Wzaa2YCTn5ro63CKeBEP1Z
JVhRv2ER2e/4pSQeT8wAjXZaDx0bcmMD9QqBlGerCiX9CES3CZakvcBUv5Ws38Xm1T89ypA456X5
qCt84g3NRdzpeG0I7tVrveZRVaw6zkhQXlgmirF3zuG4Xa2uItPGflG0w+Su3aPffLvcS6M73p4O
avTpTf5whp/z8i/xtg2BGa57nksRD68Hk+TpScjWjjQG96PatN0uweILiqt5XeNw7lOLUmORAOwj
qBynBPwCHgutIoAikFi29DmJFI2Bi2aHkECwdJLAi6/VMOTBDhd6oKj3yuTc92X+4jklBFXAzNFE
smGZCJLOgP7KZ622VNA3GMv4X/Px+bcxe99MBoZEpre/z9Zxpz8farohnKFZsl1HtjjpzhTm1wzO
8j+Itd1oSalmY+y7SoQbAJ78kPMnqKYAotJTjQE81uarzpevyvwMs9nvYnPhiYXwhgO5Ifrq0UHd
8Jvlqyb0nJjSw+YBjS9ExkQFY9YLyeS3crrzVki2Pn95htAvBDSFfHkRT0vWUrLxO7Ju6eYYEUJL
Pgpqm6y0qcoYZcZLIKBlWzkX7G0iFs6TdQGuVlYknXgTcLeAl/A+zabycJxW7HWGmKsOLHuxdg81
CnVF6NSNvFkNAcb9HwahKWOB4WRK2pHlHFPw2kNm653BBZaEUnkevv2jTTszPiwtNaR6ZfDn7ko+
vwun74RJ4gCFXs+klhrsZs6Nd7mY0x5QAXwdjnQ6QKDfuPv9aLmQCAKTg2gzTtohWN1OyJlhTdc5
TfXMa0drSZOBAMDNsvMr0EPvS9NiMYX3WJAVJ1XvIzG0+7NJJuzQp2OmMnwb6Azma+lscKVAx/u3
IKPWxZSaZ6HlWOMSbDiaSAM8qtEg6psafGYe25hZt55ZsiSUu87fD1ixYyHOPYQy642MUoLXH2QO
7R5uceHX7p60BCeW6ffYg7iKXSUrpLm+Rof2Hr/cULAhtb9Nz5RNi0dOlfxBQYSjHajpjkREdhrW
Q91Olj5nrMl4GJT41vdqU/a23GTRN8rFbZEJEIasNlb88vTjvk988jAeu7dRpLmoztw1C/j7hGGx
1KdmYhaizo97wD6b9T43ph1loz1uNoPHXf5A+nhuWsnE4FX0c1tV+l/bOz8xQjDqb3N8BE3bw1nH
dpSYhuGJ4VsPVSeFkeSLZTaFG3sfZKlgPgMQet24qIHtAyCgjcx67WFUfqzPIrH9tWjEKtZ5RGHr
d/xQrbabnLk00/kn4/D8omWspJ/Vrn3zUBx1g+LdnNTAzOp9X29oH8pXDWmagalodfrbwcL0mmd4
+4QkwOSAbrqfyEqdvPoB+3HClaSxZ2+AK4c9uQqS6Bi7ThGWLUoTQ+i5I5jdcP6TqgbJAxpVjyTL
b9flMpMTkps+d8W/cT7Ow0nhTy1hPw/3Dr12JOkMw61+Mp0SEvH4Kgv7mMK6IEjK2cs+3KN/vhwR
wEt0nYNCicw6mgWTxl5sljFd0pM7CKrLGWMFIXZvDsyj+Yvymi/czhUq9EC4EMwQ+oFL4Zs1lr5s
WvApMwjGL5qgWI2YGTyHmrGRk0nG3A6NOeAl1zzav3xoymxgAJKvwyACmJiz8k8s15DLk9paeUTh
xVEAE3TCibKGb8PLb9P0DvmkU+P6yTXTnU/4jA3n5JzUrXs5SLSgtAIkkAIf7auNy3aeCwSxRSy3
raft/H5qcEuKmJuQo0ncrJze2SaM/pvu+SY6jxvPLHQJZQMc0JDJ9FHp8L/zE1qw4Y2+7P4nYert
bN4SmPN1sIeVMVGBG8P6A+J3UrbTQbDjSNr0Fz/r7ZzmCueo7+UaUN+mGmUHcGxUp8GOaLB3VdT6
ZUx2K/jMct9vzVTXQ4vRcxv4JG22OsygxHlU+47dEszMksiuil18XO5yg5IhWK/NdsCkmV4zrcWT
azb0CtJfL6bh430NPb//Jo5V8Ahi1YGCJUJU1YHb7kOEgiU2wPrEh51sDI4Hz+eTjvOm1L0s7VUN
RhfBnjdZGNbFuy3ft4JjRXNeC7i77Pvp/wYKEgbRydYFa9REKF9mQnqix5qcS4Dxcy5nnsdM86fN
+i4CAvTPC96yuXqrW0wIxi3OCQdQKsyrL3WMfDruiDIRf5cvA9ErsV+Fnzn9WuLEXt/gF1H5Yo9f
v5oMr9e5yXt2jnHVH1k46MBs3Tq7rUii27rRM93m4JTyhlI8FSfwo+NuohhjRpEYHP+DXb0FJoQL
6cn3qZbco1KiqzxusMUqq+phHMRmvL9RAa/+zoNWxvyhlfyAxpfFz9t4u5qWGEjM+UH2N4hXQ7SV
ak5GTFxMOVSXHmVrXfjjDB/c5qNjzdtxOTlQqpw6pEzLn5tZ0xDKgqRX9lKnqom8T/Sn34MhK7Y+
ElAan8nkLgLLhK8DM7obsAXIFx91HBamWCIKhstSsSdq+UuhhN2ywFVrObDicKL4uCGHG90pzOax
KlJEm+KF18hHU+iY8IbXPx+nsS/StxjGCwpZrbrcYf6bi7uYYVj+csnC09Hlz2ukVf7sSDZtiZKJ
G6LoalC0ze4Xom1Rs5N9n4FAs1jqQOVkGKHuu8HEDSpAANXCKwCqCXTDBD5lk8z1mMWnHSISgQG4
SOoTJNAvfwcjNaTKPiu0BYC/nTTXCXYH3PCob0BGf6ElbTl51U1c+7yF22Fm6ocViKh22D+blVe6
2C22jx2KhKKZ3ZZ205pJXmvYgpxXrdSAhTT1MzCovvAMApE4w6/488yCULoysfuypFLt07Cn3kTv
zUWTIDKkh+FgldlRtKiUpxh3ActwVRwQ8mVYdpnow5/Svop1cOLDWugS6jvkd3+9kWypZ5AsI8n/
uR/URGLCD4zYRt3/oFYPw+lREwKTSOMDAcL4+ALA5GUBeKgWwklP9elJd2dvW3WPdEU2GyOo4lZv
cierwYWHTxpeW6DgsU405+OAxWv014RqQavOLDp73W5xwrG9XhRFNqYpMULEKETMMO1XN+qWbM+h
a97O2RPQe+qBujYX/pNuKamu3GI0RetylCsQkNGQvnRB9WJV35UNG23n2gxjiMviphTa84oUjA6a
n5nX5l9aXigwfj1s1QDUMqutjPvaNSYu0ngff9AojOai9aeEhsNzTTYyt9r/+/2TfKkvJXflnzmG
wIuaBNmMK+FsBsZzHPa8EjYr2pd4TRxNGlGVdgPQZ0k76LvZZ2/PDsca/V+6LZDlElpTp7MhPzrm
BKcwm7sPPWfaqd7hybrfGyUunlrQDNlGIC1n5/bbief4Jz/FtAdNXJhNvXiQry9u36aqD+Iqfl0e
8iUFh7IKayAd3Z/5C2Fz5ppXlXxY3gG70kXhzC6p+eCs66V5EF5zqxeWl3y7ZhBpugrcDqPQ5gzo
4giJfG6cBqHP9j+u7OS5+245iUO4XemkH/DWwHVQ011CrIAhPAl/jRQzXcy0qxZ3mCkGZB/g/HtJ
zlsSgkHWPKN3qFlyudYVjg7ZymrznI1fHJSl3CAiTykSbSU3UkC99m0uxa4YECscTY9SOSrioMVj
HJXI2My8Q57lF0RovsKKPmowxszeNvhp2Gsv+9UdfiM2m2ncj8n9wGPmHjZXJetrNe74oNRBa1Ah
/1OkwaBVUFTNZlcosZeEbZTi7vPMbteEdw5hb5dbX3BD1ceRFcACZkSoS1kPT/fTkR1zsvlJR3ju
9TtP04tbNGxxAJepFJBUS6EUqNrWWpTzjUYHAsEyvpoLO7kB5Qhas9Bq9KEoVJwzGhCz5oizFBgL
e8EbkfaMm4eDriV+anb96URi8HQEty8QJAeXfjy0nxNamCmpXY/8ctWqLPcAi8tLzm5JmTVGGJqX
ZHIOJz/BeqBIlUK4AAt9n+N+tP4tO5G+YXQ/DRgkOh/8M3vyAFFFLfOIsp+1lfa2ZNrUe+wJ8DlO
+u4Uvp7srMnqNKUTK0fg6j61dBsu7/Ydsfx5HdoJZdJykbrefBusbitEmV/7MoBk2qCWSXQgwtBu
PPAeWZSB6+jxKt37zCVqafqD4lHKZQl4RH2838Ptps/SKWa3TI8shtydkINPjNp/QvPxjxsK2Uqh
m4oy42rFQN1+/N8ZE9iTXYL6i32lihvi3daLP1NiS9p41zSa5GBUTds+h1Ead1fAbDZey+yQfhhn
JbBIuj5W8ZPocnTLip8TSJJVr5q3SRiiDHIvw05DT7iDl+NV70nTaUkLdWpdWuX7GS0RxPru0OXl
RLYAZoqG6Zv1YkIJ1aZNPa30NIrpndGO5Gl+bXP8RVQtt9LIj9mOFISSkxxshhiu/L2VJafABrus
H6wvi6GBYLSv36NKulrH2PD2beRimRdOExW07VUGY+Fciq9x3NiKuopyAfFUn+LVPPyvZabkBsQR
4uuhKJwPe+AjjphZIPdglMOKKqN80OGm9DCTEFkrYmCVefnHqIQzXAr0O8upPsK+faMBwAhScKJI
jj1dm7W5JBZ2NIvXIYOmS1sKX3QDl9Y8KfTUSdb9rc+fJERJHN4N7oerN5cQczJNgnR85OJTlo0p
YP8nIR4g4bmTVlWoMTDJSRQVMjGeA8dh6jY0K+He0aNX09I0LwQ370+laTw2p0F0NWb1waEw98QL
DcoKIUfjwNiYHJLVviH6oX+NyU0rZI+AciRFtSx9U8tGs2Gsfmj7KE3NTC7jCsvq5UKbvwBMOhSB
TpkZwDq4botFLxPnAUlaJDUnynIN43ZOcuMm7Fwhte1/ivoufnMf+khwZQSdvLUFDVSt0OxyYjFB
3I4SL7mB/d31sNLfvjjArbh4zRyp2CHu/ZBBAGSS2caEiUZ0ppgYuLTdLbre099E57zmpYT2ucB4
jUWn8/xcyuZcPV3jJ9ndrYcbD8BSA+T+xIkEHxxh+Pr3cnXqNyYzDz4HixWvYqXRPH9UvrIjJrlD
m8FwlBYwTE9L8sMMbJROS3JinPnTRwqmhIpkfWK5uIonc7GLFK23eXGEpiN9aQY0a1hkqxS64Xmj
/xJRqxpno+F7izExfo8ujIkexd7xEmKGC6lqHrliCsWPTQXARJWb3uTZ8pRrJOSkWtdjw0hzx+pT
Kb/4tbSOjY4VN9KGnmuw82ahFntbuQ/AKZii/JFbxWsucz3LUXHjGzXv7LDaNJsR+t0ON8MtFuyE
iu+9afpIZTq4X0b1SIVBOev1nQOAstCsKtxCgqGyXmr0AJoKgSqzYy2T4xAu/K1z6STldGAizS/h
bj4qc/rlD0YodaVOAQjZZpQ1BREWJYrzVijcKhsXI88KiJzK90E6zj5mW6BQxpeq0NMROGPPkMAJ
TBwj0ebtqft5+CBMkjxmJZ5zf+q+CwKLCnhXwMuL8w1HZhyEzC3eKxTg2za/dvfCxEJrkM0C7v3g
x0eMFfcDcBjTo4fgNl+87hbZPGb0uycsrvMOheHJrsd9PNAJRCoMEgGzLLMaWDiHfQ/vU1ulFGL6
rzUOC0qFQo+PnU1Hqmq5FhmU8o8ySaqnrcKOIsnbfe+YrEa2PhP8Y0Mk9I7b8SXsK3Hd6Veq+TD+
755PehehyBzXSFeD5N5SXdwWpSQIjnNLRnEYYVCBy9SMl617RtW3JOtuT52IzT9UNuB0ZNiYqLyd
hSX9dN2Hrtghe7cgRewgQ+HRl3emH14UubCZ5ONxw2GacLjL5i4Ok8qqB49aXoe3xy6wE9RC6+C+
WTtCW826eKVJR+4F2lGKIANbQnK6gCDKzDZXDCnU/KwnJHPxPwTJ5VqB+9771MJobnpoWdc8f5F0
Xrl0xO267RfkOGdoy+9oC1DJ3Ho2RPQWaqqn71/b2y6vRUaqY04QgLLGMgC3GRD/spOELbKCfCoL
MerubRo/C1vggZ+Dl85EOrPixpAZTdoLhRzV1W89KgyE7cUq0YtY9IAQsXT9GkbREcYx5MmbfmHP
jlVHhsaBm+NRU/vNTnBAjduyIzrXo36c6WVkKcxNfdvdZ6eauzXEQUKp2aCGJWaBBODOHfshqQ1V
GPkd6lkWkjF4JbSyYW8cfpE+0u+35SY6t8z9vzC+6CjV71tB4+0wbPPkhULUZeeZBi3b13E5MLuy
J7oAQfAd+9lm+4RCUfB2f3O7gb65an2Us9ayQLAKDGRYqmIgKWi+IKG/M+z3kHc/eALcFM93cyIz
0oiTGh639PcufCuli/n5nO75ylMTDe1oSboCrghircCMKz8FUbK1v1atsyGt96DlDOSwAJbFbixX
GvFN48hAP6AHnNUM8kn6FMsxEImRYEwmoaoRJMQjv0KA+lArOjIb0nri1JsSKminxkjJEtbI+bQT
9FRWNuDyIicpK1AHWAbIxVAqdnJc9vBq6Kvgtyq1SPfiK9oZdd4PJIbbDNkRM5C5LQz5ba3XrfUU
pXWpFiY5MCQIcluF9gu/eENVfq7aTJxdvAwpawvjXbXVutwNalSNVvLgwIBKq4K4CsKVaiK1iIH2
lepZeb3BZ8moppiTEzHUI8KFxtFQOd5JRg4zaAyYyOwqXIly2k9EKmleC0LObOmeGnJp/JkY3cQM
DsfioUQnDkCkbuYJdZ2v8Jq5wQ6N8KbFyk7xDy3bM945PWZEJwGOdkl/oAZYl4Tkf/u7nYTWYlVL
icramXxg5w/9gMsW3Vz7sPVJkorhxJ/kuAN93bfHaK2an0QnlyFNzQe/0/BNW3pf4UY8LJdjuxyh
k8n7Lz6vATZe5Sjy5ufXM3z938SBgz2ErAcGzHspxVwqD9IHv9QU9JkOE6Z9ARtygG6EKZlsE+QH
WB1b1oNcT8H+qVrOZOIyJqi7pz9EivlOyFirCKPsEx/U0ILZRNPJrUVblunAbsqJrnaB2+xcYyFQ
JImarBsQHeIfVS2wHVV5UxLJ7OWMKryA3JAggtJO8hMY/+9fu5CHwBdbMa0N+rqXw8JDr60OVumr
v6rVujQZbduwpwRIDhAZRkGZsYWIaTmlwGMONNI9AL8Bd1x572oo0vBkm8XelzL8GI7NLWaosKbQ
Ud6Iq4BiLCol1Dpo9SZ0/2YCpSFnbbrZncwDErbeVPQVaIKV3r5ZikRjC5LaITktcgY76Oq9edQd
DDFt/A8ACT8J9brq4ol7bQfHoSEk+HL7rJLhmY7JxbIBqCk6IKNQXC8gu1Ve71vlrJNFf3xz2JWW
e/Oif9LK380mcCHZo3wCjuKKOjWC24UuH0BMTQYgQyT5lErI9ZDvtAPnDqiu8nL1TE6+s13RIWG6
wWTG0NSHTiV92sxyRhN+hyIpNxFSSaY0EWb/UuUOrjAisQMaVnbb9KQ2l83oNbnrKr+TDTX3lHxJ
hRJ9hK0/0I0+u5VfxKJ4m4XKJwl+yqqQH47TywnxfAXRWRhDAyWviIgvxPBn+xaTFsnMLtu/RC9w
nxagBJ8CaM/CQnMV5mvCcTlmsSzARjFuHXxjT3LiOL+YHH6iamort+7RoowvbERp49VeMvJIpJXL
xgfVjT48YunxSu2mi76wlihTTyD6pVH51Ic5gO2ct9XUaqsVpUCvkHohnBlUuS5/uI+f80NNwU0g
reshrCotStFgrXF20stTHK8IIFox/tyuvBlmeH4KPb0qhrDHb28VCegOpRZWPo+hHyKsFK1Y9bK3
qvTtHaWvo/utIE64kFcIzSBz3SSeM27TmgMsPsBGgT1pSMHadT9txIR5z/sRbg46v9FYbihat0WW
ec0Jpvrq2Nkif6yUwGdg5lYW9Ox5lLWzLFYdvs19AEJu3iWj7HxNCOvZbuIHD7OYOT4ubstUNZmA
W8hkhFDUXnpll/iD6nZqht0zFHb6JEUlKkJ0AvexZulmILzHLEQPC2+C0roxsYuChIgTkZYF63J6
JVXYP+nPtmEtw/uioq0ehhzZs++j+cYX/gJ1LMuabhpSAFHBZkrC3RlANHkAXZa4myI3nDBjm/O/
WQNtUXoPU/Iu2QkLZl1Lc7aKiXPUXswpyc58cGgG+sKCvfhirPnpIWNwLaSJWI50ZmlQz151PxfL
mXl5pdmhVONf5MK94zd1sT5gCI8NGNKElvtWfTIF5H7IwxC3DtjT14NR4DLYzISBwZQsGrElIZkt
9e2k/uCpS4DgdS/HgVMRi//oeUNDZHD2wXNS2QdEPOh9U3OvsZX4mNpkON7dCQJf0kdtQKjh6Wcj
aW1Kn3Qwu4ztTGaJSzhtkBJr1lSYNmjYn0Up2I4CCcvv1JdoR3AsQCYUxdQZeFDEL4SDaZvmmBZT
8024V1xEtGVb8oTgC4MChkUybKjNra7jRb1GmUWeyhiYeWFJ8sCSmI1Fs+yW9qfKlZXsLqAxjsaC
pDkTbSk2AvBOWXc1wDzgRTyvaerJNFEy4w0EQdfNtFuao6QPht5p2UZCDln5pa64iRgvGO1Tlq8Q
Obx98pIEAO3GI7JNHiPp2UwKxQz342/twwCaHp0j35tVQSO2A0UnAcNa3DtUy+jWyYoiXjAsR/cl
aUwpp5M7h31VOApEgaQ+zNKLD8ZS/Q4TsgNW5AikWTalh8ataFL96myBb3/h0gn5snbNn7ZcfKBk
+vnQ6RsdUPY7Bf9aEr+WtvPZr9UXHk0Z46yCRW/NGTBoZKYxrYrtvP71zXqe7uPUjRwzzq+jVW+i
o1wiA/ojeXGiLw0TYHqKqnTi6FbyuTkcaE6SffRq0trndUfrGmhi/ryRgdQNO6OTo5L8YvU9DAAb
8hCFCsCUzQzwhTYMQIt64Aoei+vmXMxMwykJNYCtpiWdlenAHmjv+KtlTVMw8Fro3NcSE9SutJY4
Iw1TXl2m1I7av7GvAusd/rHsm6LQ1vIQ5Zceqr9g62/isw/2XHYrkcfn7xsSVy2Leq70Tmsjlvhj
MpBeW4ltyFv0ILzX4YA3jHeHDQWoeyGnGF++6toMH0YBXa2bHxIIhFbG478AD8f9Ex57EP3U4UDn
A8UHuTDVaz0O4XCOrsW6hjFzPe8ck8yZQvdv+e+eAkqcEGvo1e0wxDq4sxA72TY/XXpKewRGaGH/
YuurYaR7KqcvUe9NnX6BIic0GkSF+fTL8v3/fnl6RxRGkezB5GS7JjaVaEiRDoxqqYSDP4+ZvPrV
GP2bKUOmkwCXbmtK2IOilTlpnzbl+/JruNXPkg06xhzi1+AX32t6mTRbDkDz2rO8yT45VtbB59ZJ
S0bn6LCkxXwF1Lc2U1YF/sw6DjWiaNZ6FKJksQ+PUedJEK/+xnASZdKC6fiya3VWIkZ/++zUv2OL
bpoHPpeVN+hi2AWeXZUne3zF1LETWz/Ll2SsON9WHMcBK86+8+xricozfZCRtENzfddBA3uxgjS8
5vNJjsyafqtigJStsIF/DsIBjsHwiWjgq0uzcJOJIQ+H0EZNYvOLX/8yggucs2OJaqg7r/h6tfLc
2sjE/uWgfSiP20ZimLCi0CbPdEKqoC1XGoeiOxCptM3R6lLtpSzJyGxy/lMDvE6LCKTyEK1VhQye
AEbZS8hJRbRbw4QWpL0nwGXN2yozxroktUIHTxaT7IWaDaCtKUoUyY0D4hsSDMLkjcHB4Oars4BN
vpteYHHZUGCWin4AOTcC9JLa+n1npcSw3JLPTQdywL09OpUcxZ7mNG77UUtopiHK3DLnEMdyueoH
WeRwrFsgEZzSb40uquZaTwWc1hKGgCQLrT3SMzfMiqDcdKBf0Hc3ZdTfYb/ktFKhaTg7f59G1T8c
mIbfUfu+rGRW8ngQfsAl2cLiHPUzVsFAIfjyT9mUGnserUW6PM32RBWUb7pHjLIs4VVXoxXl1dn9
U3xaHfFOLpDoMFmMR0Wd0ujuVBILDyfoo4U+QSpcfPWhWYCxcU1YXBzsZc2wm3YNRyzPg1zaWJl0
LlGX69R/g/iOSFEi4Aq7AKetaY++NUWs66ZiugBA8mFhAAhFMllnWJ9mx+MnLlI/rBZHP+12T4Mp
FbqSlOYKQV7poXNNjJ39g/R7XOPzRaIRLlkWP+TUrLvrez4DLlESrEu/01v5jpjIPkicb5UdWe8z
M60U1inh5KdcXc5vrOs5GsgL/joMNak0bYgaEHinxzYUkpv/eLKBkNE0p4nAl5WWrdE84xZ4eWs2
8K1Nenp17NZQ/gZ7mxl8zOebRG1sxHH2GfNac4CMf1ixoLzeuoKEAZw71exU2p7psPQrs95E1kHg
vCiPbARPV81kP12MvkKA5+prt0eisXma8oNXJabMs/K8oYzXwgJjnu+pCdQ2pddHWsdfFPwD6B2Z
ik4FxjxS97vvTI6IVRabHcQT3JFRBXHvWyvPmThkrjNtVAC2l0XjFH6adbSKtbOxSInb4GvrTQyQ
DdtlasO+IMWSF3Z+/hnhXNJtJoWQYIjNykNWz0+LKDkNajiY2iurDiQy7g+AzhCSXrLoJNiPBWcy
Nl/LMfHpV9yyFwyy7N0gTAXW1K2G8aFXUp9EuSsEi5EZkrg4Eoj0TbazeZGAITNjHYJC46ARpBoe
BTo7a0Pb8iv5q+C7W7VskjLRbTnpqUE1EqDGB4iBX3dzF9JAKGEqkmzzJsgG18IFTrK+0PLSa5HL
3YgwS/EPnCEWTBmKo//g2k0WIVX3ZhxcIFN2TEmYET1kv9kw8JTgYGolk6Ca8tbOYoNu4ytB2UkH
peKD6xj4zpZGAXS/xp6TcQkbj+1QvF/LIjsrBmEWaNru4KwbMGYsaLEVkbRSSeBg7skHaLIGfwi5
nQjxPGj9FoLL7vf4NQs03kxs7qf30I1cEcXqX8xysWJIHlL+o6SNV0zK6q8NRtWS+fbYBEXKN9Nv
Zov1RL+yx+N5nMif06O4EdoGzdoai5oFn0l9y3TBRuEZG/yubT1yotwQYLhbvq/fG2rtKvtp7hwl
tWL9FVpsNOfNxfNr4DB68+2045radSCIiHIpd5dvGUH6k9RT8M3hPrtT+9PQYGmXE4Jkw8zyNITD
Zj2luQj82JOAKOBOHD8G6iZg+PSalJ8P9Kn+t/FF0coiONdkG71HtiPue5mAV85HN2BZVC/8tn9J
okeLE2FaOa8iUXqGn5I495Rbvq1wDoW7vWgvXtbrxIF1xCHCMdZHSzV31rjw2mXS3MnJAV/7jvUb
jVcAsMM73troNBGIKIV0QcOokUiE0sJfVI9ESUFlzZdp9ztLMLRt+v1Hn1opY9dFhdHAqZxoDD0z
f45SFPV1KdwIQ/fVUwQGRTRoCB5UPn1FeUIEjEdEK+yfDo0kp6JzReO6wOzghSlvN6ZbwCRd+RyH
VVkiVXu1jmzkGpksxOaUQ6m7PysOmJcMKh0orkymxdkLea5zA+6ATyWLwS8P0FNf74bUPO2yrufa
8wa8NAbWCzwYPf0qNNCRaBWjmSuUe/topr8e2xtbyMpfbO74Lx2ZhcbEP/FxrSjE0IYYTj1DjuzI
xdHnD7LSdRfkdXApBUZq419b8EiJShP4Agrm4EBHcUtLFriBOcGlXdlcWWohZo3vswU9VWnSHAKy
MAc+hDqQWiUlC09yIHs6x+v9fQLf8kgSJ1CY7tFCjpwhAwFwBkUmYwnM6gLT7orm+EfK/azKvEYx
SdoxYHol9WCCUppTFdVKhj0V2Z1vTY6JM0AuC1JfbCcxhF3+8DEeqqYo+aRAkUTfY4mCv4+G9+3+
k+pgtC2vLR7iyspU/yj61jVyf7nmyEmKtQvdlkPrLPGcPIQdMG3AP0R4asxJij4LXyTskyhZMMUE
CFaCizFNP6PSHgEHXyvTqFjD9fWk4MMT+qBzma/g35fnnnGjDarFCMvGLlrapFCuWMLQB5e14V6P
VMxDbCZiy3HBqJw8zCeN0lmDQ2CWBZAm+KXIYqV6Sfas86blUAj9JMWGiqMjNXhwVagNL+gd1Pj0
amJ61Y4M7y7rVWoF1hrtGsSvc3ox5bUsxABXlJd22F+ltJKDuZAoyBo79wshRX7e3fzggcSR0Ui1
hqFo8hGwDJ9M3Zun5+gKcmPrhysH+LkUIlDwYtXZ+kbZbToOllz6fyUEZWs8mjpfs4rQxxWMqeGe
MNuGeB8us1mbLf11rlp+/Mx5MitDNrMajNxSm6QumkwFn2F0A8beaK7T9NpQeEqmr8O3nZrsEptE
f27kqQNsW/uuiy04zOVWLW8XJK2ypqpbY8U8/bwSGU8VHtN70mFtX9FDtskpzletXnYbf8v3ovPx
oC+RUNDYuuacRM3nS6SC19kVmhl5x1eu6ZGbYUgIzV+0q0mf7Kx3IRNHgYg/DlPkKUugmA/Dgre1
xte16e+vMmhQKavhVvvBftfLeeK+TGJZh7pvZ+jit8PWnG+aLDkxMr/NsxZyeW1uZtj282Kl9bAD
t4znkZ1ThVmU8370H3A612E2TTElBnwAY6Q/03LEInlLHSNoCRupPBx9bKxyo7U8+hgQs0+Jx0RS
2IPSQYjPRw5zqa8FK396ZimY6daryIeAfMEwYbugqpmILDRdjSjEPzJdZ807QMHHWdwv7ocX1yI3
oLw0XTw49jqNmq1gMOTpnuFa7wYyo4PsQnZqqRMiw/cfgTZNwSdHjnIK7eiRfA/Gjr0UJzt+cJli
VhnjaMi28D65JGXXALZVDUO481NkSCHQHJj07fb1TYWM6RWanZsERKMKZt+rulDdEjzA16iW++2k
sdOLDInnWUo8CpqAU3+4DqK9z6pqF2RxkoE9/rJGyg0wX1P0qkTY+TOkh3z1V10O7+N7Rdu5ooh+
pjNbcNTgK1Td2po6IpHSFuicdwei5yvKpj3IZMXyUWSfC9atzhxrxWCzO08bQhTCOHFQtGf+999I
3K9QiPJHh92YwraE19d9ve9rZ2aDo6UtJFrY+Sg8xMLwv8oAI64XjZOIsRFX6OuZcocb7DMBVAM7
DkK9PiTBFyk7f4gV9HOmKAzSQuyjYkdhndsncyaMVuyWmYOgvgFt5PgPUceqRTtIlu3EJxz7bYYB
W+xH1HvrIDdq8uElLIqKfGJ2tuxwc/19i53g7IT310cNfVbTbS7YQModf7WcicsiXtzg2C2I703Q
Q/oX6rCbgCas9StPp8Zbf457S3PJSOjFFiyyovWH3fiUuojnfzvSBRR+3iQtFyuU1O7i+tdOEin1
nZGDKTxU2Qw6B4O+z8Y6gk/Z7R2By2Gx0bV8uxgPUAV1/8lkWKlyEsRQE3h1PERrDrHO9e+nNS0w
3xCzdRRhp3Z9F6q4Z09+05BpMwGOcQAMxwMm4PwKL4zQG/evNzqhaPt3rGpfgJYA6PcJ6L1KMv6i
uXeDG0V7fbrWPV9eMIpPokOlcA8UectYhfFbcd7GJgPxgB63/pNPbuw6eQ7lYdATs4WJPNtzEtt7
CLmZaLtoONSCkPxfcO5UYhVLo33VM8fiqIcvwUc1VcGX08SGQJMoXpsqkGhFWy8y3ptnLOXOwNEC
Zm1X8EFE0OJYUeSdzPcz3KemfA7JHYuLfFJMyBkKH7YeabG6NcUjX4iIMUA8Cwrvqk8smQuBzu3m
2EOrSLc9sAN8zyEl4ZWi3eECCRBOfTK2zZoDmdbuX7bMsDQlQtlDHRoHctrRQlxIeGgoANMAU0WK
hW7IsryQ/YH5cJEGi/BCucereaXWKw2UIErdM5NMKuMiCQ0ooc+HufmcRUFBrU4My/mq4we1K+r6
g1iAKAgXsAsF/Nkfk4/q+3rlS0Sqkb6Tm7Kv/qEHq/47LLR5HQuNP1L9lmoqi+6WB3Ahi9Z1yUnB
N8OvHNOb+48t4svCHHlzyqwb6Lu4HL6trPDQoAM4PIXHwRUCZwEUIGQAONQYam5cJKoiDCPpbTlF
qlwCAKicblukP8TOqw2PYeuAFv6sTXfNVu3TuD9OiqBn+t3OmupIZSdNX3li60UpzrzdPtDJomVx
F2gchYqTZ1MwuK//Qr9v1cJ/JEE9C3qc6abMntZE8agLu++it4Q+C4QHxQZ/Qn/1c5SRrThStcJh
2Enuv3j6PcmAFdT6yydYZg1OwYzpJrjeDDNCLqFByVie7sSNtRP9YnblZO9Km4T6UC9qanDtN6rr
30INFZY4b4gTGQqsVvwGIT6cLuQO8O/tpmM6BubWGuMStWK0gpfCzwdZuoIE7UCA7uKoqZf/MOIE
SB5M53w0pIiiTVmABYgWpA5CP1DXQ0v8NVqMZCuQAJ1kO63efHAeoZFD/lBH/CKrL2rhwhsjfzqg
AeBqSHKUFEa4qAC/vHRfO8Wb5DrBBB8DULSEomdqAEOLXqOBGYqGsaVEeUgP1SBpanRwLTvoWFkh
iqFf6/pno0etllPhcY05MuwhQaUha3p3quRv+Gdk8uzRqwawo1s2hS1Ychq0evmgvOHJTvwvGNIq
He6mAYP4wVJxYtU6uAWxpe84bTXf8jhWYFCkRNzsQzQEZBxXptkMite+7BQmJW3vY0UXMZnIgyfW
MR9xx2MPrfReYGFfG1HuqNIFNXpCuRIoXuWsBxu80KAtmG605j9y3u5vo7GGXEOlwkHJ/DCqf1vk
LFi7PcE+wkfyXI0t6s+Ung+GjewSywAu8sqP8lUsPp2Lr+tU0zfxF6/BQGHFMdLZBCPYCqzSoyBH
uXCRoCBsdCxx0M5tN1ZJG8h3DKdx1dWMywsDeiPm0GHm+KqXKJ79jsWsbcNFpIEoJOjqXn7k9xCK
WfpL1BGqd2Np8CzmP2gYmFgA3HKUwdEOrFby5DAkhobFEqqQkQ8dstpL8fd/H370e1FkRB9m8hfq
nFcUQr59upNtgiQcIkcvzU0CYupeuKCN9hqapiFWpR+/DalR2+bEU1q/skCEqmvflK9fuacE8TMa
c9iQMgCCd+POP24k/hFs7B/uRFjOi05DPVJsrgiw2cqjIVHXyNzwchqHBVq5EUIDmOBVQJsiWyUd
vUYiLN0yJ14A0wl9LLa4UNjCWeQu8lcgrgGdwR+aWFDaQBxqR1O3udLYa8S/RiDt3d4exNmMl5R2
tHv8HA1r0bzJvZKSOFst4eWYciaXw8umO+bYipB8+iHJ0ec/xhuQDGVPZzXx2R3XepB6/NzHBHMs
y9pwkyY2/zzKPIgbUO8IOCJh1UhW4HsXDZfgKQ2xUfIx4EpRNLOYUoWrKlJF4B993POGy4qyNjWV
sW41X9uIEdxYK/PwRTgcvxIZhcShICQYAqdCrVZj1AzLYRPilzf0tentso+IhEtyLt0ksD8/uFlP
OtXMzxUdLgIWMMfMCfGlYI6VvQqgNLmhvWrE6QZiXrlN0vnEckuCSNqzDQkc3vU6eFF/l4ucEHc8
+LCyatJtzRW9EZ9VBxdYXPV1gjbseLqaqcQBKW7RkIA0/T+YJpSUGNeoDC4fiC5Hmrccjg70W/EU
WnXgF2W5T+lXpVn/cdrVUGiEEbptgQMiYtJNiCeNJz9l5DuGfnU3GjMD09WE1lRwIvlq2jGo14jc
jPIol2Noxp7rHxA2OR77AtUWAYmp9PCxgiYKlUfz9NgnLa5u5npdRyqLM1IuvtNgMfYGFO+TYPUj
ns8HG0cVjw/tCW3KY5lsMEhDq/Jgn6LkzemIFnQh/Hq9vpkmvOWYi3cwpnFBEusW4ipMIvsRbIN6
ViLcbiRCrzhCuQLgaYsIPnIbjnkwWeKdxElKyC+8bdDcNLQIu5YYpHeyd+b3Jof6Nz+lY+YoevvD
C8G0SQ5+tQX1cIrfUHspRmTP6k/8Bx9uTX2jq0/Ptdvp89FFH0sGpznTCiOBbRdSoty4xeEb74m+
tmA3PT8+bhpfwVxZ3fdQsbQ+TnyKESg8cM5dj19S35Q1Ri36iyzkyFIgDvlhlCtcTxD96bn+ZGGF
N+yDhRBylP2J9xSsA1SZYBgw+CO+3YmwOVEKXA7rQEEZYfECOumYSqkstHb4rzIYvPscf6hbB5mL
TOg30qM31iwbN7atFShFDFd+f1eYwRVtyR7BTTODjwaxnpmdbZDaAXKVsu6Brjy12dyGgZ4kd958
8zCFHdfz8NeGeUpF0fb0Upup+dvlIxWqwbH/uc+VWMcVlkkDhOQ7CxZgJgJdvFygyXzl5GSQhRo1
0MUp1MYpSRkxrl7sFYPghUAOYmWJZ//JrxpTpMwrdex6sthCGMqeeoi4BHPK6Z6yglaVz/r1Q9tp
vqyngwPOHzQPud8Wz0r6Vi0KOyotJrjnL29Tdd0Vv9TH48I0fBQcUp/hDOenT6RYQU2SvAFd4iX+
gL+o8c8jzDItH6EDeQeftMDbILewyfFyO9JiOXtdpWVZ/FXNXfY5gRXvHuWJLTmzrTfsFErDqlCw
5SVmwPpnjkcWWpt6DmdVbJwcolssyCT/SoealK1PKlgMEgM8WbU8tDskItyR3zeaHFklWrY22Teq
1we8v2TLwffD6aZq54j/UD/RjU14ZUNjsNBBtPt4dhCzEjBAbEnA9D86kxcuFlz/T0az8UAS6yXR
fZ7CuW/k2PIi29Lk+L1veAaZUYY9hff0G27xZDIIPdGOtXK2dfjFkj936naZ7EQCdlgxVKPbUe9A
lvx8T+JNmOTKF/9JJyqFYv1DufuTcOgNAiTDnxwI5xiRwT/TcFiG6U1N6FKqF8kN4ZtWX3xvbVKm
kWv9pEhrRqGJLCqVNeR4Dw6mkZdzkGzOGUykhPCDbfctJ96jCtwEopjWc6cbSzghO82bRTB4GHQo
tg6JDDxBpU5uYkNARvVgGJhXWp4LwwRonvkk9s/Todkw3cpVHvBXfbrY1ccpLxDLoq78rh1fFj5t
MWf8YCNduytEsW0YAFsQ0yCZRB/lNoycan4SVq9HZ3M7NwIYSWO5o6Ko3yXYBb9yAKEXWHMaHRvA
8wnal0h3knF8robWLYxLBET98rUvd/pH8THSl4QaIkK29SUxqDrD/TWNUnIucc8vNqZpxTcc4oYu
4JvaIwuV8i8GgBpFAhQntR3GcdwMKXi97Bmm2bcFnnI9zyxe/OekD48NuAMIN1kFnkrCAE+kjtz/
ecvibtct8ArsPpe0nf1bntqAsz6lT7NLIkBYf1MhT8r579avquRSyMZCQGCkng3CmrylR0sIjGeW
CegUiGUBMkMQMHDincAQdJZK4GTAQAkYnd8M73G767Dz+pr2Q6NirmWScEogwygJ+eYZfwpGu0jV
Vo2+TIF1CTG+92+8NVdpZK+Mp5LGns8ed5GVjEAaZff5OMXVuTIflgFSLomWRyD7/E7aMcmPl7tH
bODe3nW4Nh8VTD1F9bkBdykqL4TVlKdN1LGrZwoUyzUT3rPGF02vhZrDu7hGxBWz83qmCwNLW72g
3Ffuaef/jhpnQ+Q+DBEkYtboCciBdS8FGP7IdEwKTcNDvkC7C2JdnheVnbU0d4HDb24XJettFXdq
WtHqOGDBAPYV7xS6avh73+H9dVBQL2ABDUBaddSE/uirHYgwRPx/zGy5t2OWpOdCjUVGJLGpf4Xp
6lJlYFF65Ldnh4IibJwxFAGbQqM3dpWqvRYHwJgokEnCM3lZXDwwl2Qz96vVpZT0YRh65zZ+XZHe
EfCK3+ZDnXlA/M3pqUHK3x7/6Z2phywF+MPPuboZGHHmk8A7A3hI5uozFvj9/FnzUZwempnUryLq
A2fWphhHCLEVFQsAekz4S8k27OothMnkk6JEGbF2mbYDam15GyTpCW/URCCOYyd8hf2R3uxy86JP
jGD86L3laVJqwC4r3I89N+SSfm9k1eLGNSUYL8Sq+Ss1RhLLs8WvpTW4KKJPIU8HisZ3wF6Whh+d
9SeFEr67w5KyCYRcTDyEW/nWAM34mqV4HggHnd8TZ5ySHpTZg5ATD5Opj687unuOw0ahi9mnndh+
vsUngLb9lvE7SOCeQ5qgxJ4FKp2JFxxLSlBMCx8KcKXw18fazEc6voQ6qEnrI4XInXG51vNBCXVi
01o/EJ+JmNc6uG0xnWkz4hIcZyi3J+ndY6//ZLfns5OD+wPld1oyfj3vbIVPIy4k2FxsSaSIJrJd
sIQhunoytq3PvUTBvZYE2Y9ELhY15t+If211ZR1M94VIpnFWQEg29G54CwDDd1s3008tV9r/6QPH
38jy4zU040Gce9SasL8ESHXr7VCMGKjgliDHzrlIIdSsg2haYjqrY83OJzc2st89QXEVKCMzKmfD
/95VTfjoWWupXMoRMs5Y5QGrZ3YpMysQ2LPsQfBL2FJjl7WZYZR7l7e952qa1CgCz59PnEkhuLIi
7+lAap4HS2TF4ZTyHplnN0Z01/G8grd70LhxiIv7kzbUv+TqyTqdc3oWr8BamVZ88J4LxkbHKVaG
IRCQQZuvMnQgz4z47pTqqcmNQO1nbXJg4ShH0dvebhuw84OyOkDzkQ+cWZMmwAB49zz1VkAoEQ3s
2IVgiTff3QSiQn/PtnzwBm9ixpN4q8dogYZrBQSjogFVrSvIOR1osTsFxye7DCp/onIgGGNXjMBU
1NjdVQLGsePeUTo5fSMK06ylbJwpqo9gh1nxN7KptrUAeO4zWFhkOapxQo2seWmeKCUJFVxIS0li
kMywytZaO7mAMjx+b7nZ0/1YQlPi+mW26RanZr+foNPgrdWYXzK3UkkjJT51QoX278fR92zxM0Gk
97nPgngFBhGrQkqRMCYpSJo0TFtYZOr66EPi2qBQF6a4HaTL/9lWk1u7N7uLK1Pl/TQGJ4Omz3Y2
6H+j/Q/C+pLGIBWlLl9Qr6leQF3HO5LMWh3M6E/woxEb2tPWnqCrZ6fWdU2R3Pp9IyfBN8cxniMJ
v6M2eyzkr8C5huDBkmFLmIDY46rWBtQrekpTGyBqU1mj/5HTU4sr2WeLwms1ybYPL7IkWoxojB/H
QCHSAc24+AhNlilxZT0A1CpeQxCtcU5YjKmcpbMmR4q0B8abQS/Fn2bBpMILyTFC5E/VRY0jsicM
/Mf5t/ulHfrEYze8WlEbBoyDyjgF1jp0ju2frw17V9pN9XuJTluxn0D8vYV+8DVhINPdRxPa9pXY
oPfX0seR3wh74YWqhkNjnBAlVZsfU49wZbjIE0hjmmIax9Jek0oDEFII+ebGUTDr4GXA1IleOvaH
CF7q759m+pPjhD9Uvpwt3LltQoaLSour1p5Ll/xyVORamoga8iTwFSqGDwDlS5NjjtT5zv1QkzuO
QD0zuy2GjUUmkZvzrB5c4DnNGUiR2x0mg+glTqJTYrm3u/7PSsY0DXuWvhjzV7YW5N9+rYZzIxou
5FLLqSkC/4tSoFi5/ltWZA5+A6PcMPxpGu7BrO+OXTjmrF23HbMqbLFOC82hUUVrZ7V6edqeX58c
wnUhmhu2fAYUBDUJGQaqAcNMY1gqmtUQPFgpCjtOUezWc60BK1lalV3x0hfub4EwY7vUpMdh4292
FnvoRPXyhLTvssBnmoRmhPwjlHIu+trsaIrIX8QxHofF+9pREkoXsEl1A9jEOMtD9HiWS065B/Di
s4wRBh6JJPeexvpKqL6EzIEA5fBJlDIVW9Fu8egjvYGv4yGdjB5LNlXyjsMjKZiTaPCgh9UsjkTq
91ksv5RdwWeCX1ls24Jckgo+/ZJXd4OojNMvDWGqH5YrWVLhQpuPUNWmSAspo6gWAPK0FNhKL9VY
fZCpxWfkCFViC/unqiCAxu/m4haTs8mECSYTyAQEXm+SGHnfgUojqgs0AcJunX7CHUD/zZRxTLBP
YOLhSANu4izGPIkXk+lvnmY+81u6QEW3TxxKZy2B/4x8DYJ+AZJDXXNDZzwpPaYmo3IWyWPhekER
wraRGOx7ees6gEYV6D5bCLqPmrJmG7YuvbH8jIbQNZEHaz5LeKkvRf///2WAnO6LN5KdHuXO3TKU
YqZ1Wuu24oHjG2QHR2CRIUQVJ9cVHzg/iSrRo11YtgEdxiHrNMrQ8IapgBxHUgV94cpFA+IX/WvX
Oh1YJ/wi6fHlFt3Z48u+TUjKATiAxFqijf/LlB/9WLr7RQ1Xs3egxjYmOIbEOIbv75w45mX/lEVN
7fUeXQgKZlNV1faLQBHDWEl8KehQrhZb+grbUmvfN4slxYiLhsCCNtm2/QD7m4/siRpb5txl/sbs
dbUASuj1AsSkhLYwbM388vkfaVdciNO1HOBL+w/O9BrQERqtcUkkmRXQjeAw8cgg6x1FZ3lJ478E
iyMkQsLS9BMFR1ym92vXVOozbR5cSxLLqr7v0Z/3qZUcNok17QPZSeb3x0xI0dPT0NZ6QXw3TyPU
Gp/Xdq88hOweb5DC8op1JjxxzlmYgnvGGL/0ZrxZyCPgM8r0yExZdDiRDdH42MKGSQYT90NotH+b
fLslAcAItRfMskyCRxMay8QYxdt/LkIoRykua5otFcQadPoBy1c4VVopfXMjT7lef+TSw74Xgvlx
/I7FFuJhCMQc8KputB0Hhy3lHJB6LpZryuMJesDquV2qcg2bwfxViRpuqjOFgfsW89vRuqThAjdl
dyLRoGWE41nfUDTy17IqCSf2BGHFBxPf1kxQJg7DAz/Ws+PHmkZG2XK80AW4dv3D1hAMSFTfWUTj
mp7CYFcZeFkxj/r9cH/CDm4yeumPb21IFoH49UC+yZmzS75WgOkifaY6cry3O7kRmaJ07VejtM1g
W/TavXLl3fKTUN9hx6BUNXnIR1K24X07DGNXGjjHvFe4adDqZ9YaHt6BpPzSQ2kJoRed/2i/lNz5
1HAgLQC4gProhfdJCm2U6VGcrpZs1EdoTvo4+IX+EQho+nFymNNUGTzzsFopcE/9uqPbII4aGWAd
SOpxc6/uxLym2WZOQhhAw0IZr5fOrLIWPQTYfh46n5r5RO0bCIuC5LQRvPN15TL9aPqtjGWY/7dZ
gQCrADi2FChCAQJTnKN+PSy6J+mksKLysW+XOjUmGZ0sHXoHWqjkoJqpp6r7nk5WRS9Vhr7+Pl4w
fqYuXJqxv1PeKCMD959SvzYwQYeiYjuWvFw6Iff77Bw/nARAkVzJ23de07ZlCmhH/yhSS0ubrv8M
/xiW1giZBe11KwV33KcNh559NLv+FNiExM/FbI6C0/uWglEJtWpGH2WUEjLL0csoUOPoGQJKw1kx
qEnYVSClLLPFg5gjR/9aVvzJ2oAe+DgXeuENHi/ndlGATrZdilCtysdrZAYwTvi3uEKk2HH/NLCY
XpJScLkTkRLbeuHi56iNPxM8AVudRWgyetcZ53ApXbz4NywzjsTndsnI9IiQt1FwxHP3/z+5ak+E
7rukL7Vq3FlzTUPfgimi0q78HgLCgOts1SHB0QDErXGX1kt5X/vJdTYlK68SE9ZlA6LiNeSc63zc
99AjQuRU5qrkcU1o7uV5gwt95aogldI2yRPZLg5t+xuFdpH+waS3kO0gAvFqIv/TW28crgtq5JCN
IW4Gqi8KwHLeEwgs1dz4J/Tb9Cm/Yg1SKqlJBErni0k2JPePiGKSjRExOl7kZ0IIW/Hh9JPeCBme
8x/s62Oit9IMoCtoUOraq+4D+9qKeTJpNTnTzlyjmXS/rDkjkMeFPIE4HPWQLDPZsNGIVz0Md8Tt
ImhpbHuPVZWatIY3ldqJF3n13UTG3LGlV41iR74Q27lJk8aml3I9SCnHH6/nkqgc6shKgzzMwPwT
HbqrSZw1nWQDJa7TFZ66qgBdfRgZ3G49QdNTISPDC0HirhmjpZP0BwJ1hcEpLFmAMbltZX7qDqya
ORKy22z09zTx/J+9rNKzK1x7Vo0GuRbgqjBJeX7RkEv7q9xC/4eDogwlXYmc+WEsZYQMazgU5h8Q
EKHIHx+dgzdfxKInwAeEHNas37UDX5tYUCuukppcDLUETos8Mv5HWsktKFUL41grlIToZqYUYo3M
1b4XWtMgi/9zqrsXULos5nGtAtajbrzBhdG9Eqasf+/ZsASqU7ky3IANULTSpxrRey3s5jYmX1gk
pZab0wlHz/xbWHRdwztm8yWKCp0FnyqZmRbqWk7agKbt6jHfy5qsPs45Gjroe0BOC5ux5FZbGteJ
PwO3g4V0h4SrVw5uglFgv9dmxr8OCmidfT1XxlLamjUWCMFRKV8NOte2wgciZ/kzeBRNbZz8aeQ5
aKqnWIzNbVCuxvVHR7RDOnPgpBxThn3NtIJL5bCMoBTe3DbHzL0qx7IdCh6i401iW87Joxuy1+lU
q2l5Hd0a420xffxMG7ISRPiaA+8wJFGbduVGvLNhA86Ye5SOg/tZw4sZ8vWwhzgLDbekGBeiKbka
ulQ4sal1rZLScsOvKKMs1cd9UmGBjTaIDKZ6u2ikies/+czxBVWFQm0bLvmIfxW4aDLcFw5dXuyH
gUE0siQrp1mZDfSFLALO8vWeNUXjOSCLCNRLT3fGG8Le8sjS36ZRVoSgceR83Udthmq/qxD0Rjic
cOrp4l6+6PzfuapYxrJNFdsMxB+3qR1e5dMMqqTH9tMqW8BLqicgvp6y2qY+fmjzWudeLxwj8sgR
TDNc8MRgjX9zXidGvrp4lcX849e/tzX46Ql7IdgqOrzRSAclm+z6Eenpuov41kbNPv81YxH3EFvs
QuxRaTnEogyO4GjT/H+Py6P6q1n//iNQF22Eqsin8FRfUeRZY0f0p1jMaKseHz1CnBE/gKcdEwg4
bFLdRP0UlofUpw6+LGg0vPbErJsaVQLgWIorvegBwa1wQt1xikzETnSfRFEhx7HTbCmYnIrcxlMm
apCQEU7ku8HVSoOLfjtq6zzeBpCFGt+AR8IY+94XNt8H/e+QzBaot+utC8t2zjJLbcjbO75w0t4Z
fvy3shlUSwx/Yr3ejhQV1U9nOcayYvSNDDzOyV0xmjDfq9rZDuM1Nyd/kkQb1fWVnjrr17E1RVyR
JA3QKAoXNP0eyLqVU6kWdRoHSNweT/FbQ4MnT4rmzFoZaPgdeblRmFJ6it9WWGmNvXV884qoVfq/
Dpau5aMwEJVARqSuk3Tsyv6i5dUmI1VFacrwpibBQL5mpRH2sHLd6wVTFGQT3FTvjQ/mVQN+rmyJ
M16rATMmJNlEj5BcQkgioREQKx50cKyjQ6rV5JXBTZokEidYi63tdObOR2eedar4ouOOC5NnwT1I
Bg1yrPV+nOJy8r1x4WkU35tHLHxsAGPb7nZB2mlLjo6KL6/Rde+TwTB+QMWyKMvgrycbgCmZaA14
t6vX54FI0aU5aNcYnQrIhkV0HLqoGAr4S61vhtar5HnoKRjd7MFjdOGkGE+ssYtg62fQLTdbfqHX
P3EKkzy5jB1KybocfDvzdwgNqJoxE2wFZn94mF403oMaKPW2bZbl1NrbtkSQ88qMjYVhTg+q+JMX
7+5Gj17hL96/el8jGscfJr1np+MhpBEdljeAKPZz+F8HK5sauqXKUvrUko9FY1lfUAb1Q0chZ4h4
oJd/t1j5BQfDRonRBRiWPrN+PG1LGCu//KaEz7T3ibweNQQxz23jM9XOMxzJDta/kKIX+RYYa/fV
biZWQVicPwxl+su8W4T+IOT28+hEE+GNgXseMuobliQcLCw3g8rDPoY5GSNYJ9Y94siWNK4qjgp6
uPtUVDjSnDtcrQR+/sHV81NK/cFp3Yg18O7ycnlHfjhXMNBvFOgp1946UmEPiT+26yhrU8+l4ZuD
7Ceu60zjkwwHnFXT3bmR0jG2EKo9tARVyXpSj7I2P4z+TZyE6ngyh4gPf7QxQlr/CjQ24zDia9Z2
SI3SwLrBU+9G5wZSi/VbGyNAfqoRPPTlMHfdKNzzv/CyK5L4KKa2VCGHvIgUWptDfyn91vHczEhR
O0xgnKAQveQvV33+/U08o/Qu0m6BFhYwihdCDqC8jNb2PXcqLSank/ENcAkJXGtGlWL94l/+pdWl
rA4nFQTvM5WIdCbkF6Gf6Zf2Rvh34RDzKwwWoP8/Le85GFTeVjWva6Ezomj0WUb8HZXkP5mQGrOh
whk88MbzfqN+nGXkaLSEj2e/LpCI5yFjgCdVxLnlj5MdGclJzEcftEdY/xdtQRs3kQchhPAYgxpv
BAf0D6Zu/xf40+LwnIZlbvVunqgwMY81Qa+8KdWiDzsXKTg/8rTlgRYN+bv8+LLQsqnBX+z+JJS5
rEg6buJ8brjTtw7rsHCClyNItbPBRnQCc/GMrHo4pg64/kpG+RBelvBYXV1r4eZgdIyF2LKVwndr
dL89eQo5/7PeXjGDAiibnGdCf6HWm66v5l+f83aKX1iwD/kXBg9MjA52MuS5/hCnpI2iEQB3GdeS
NCG8N3TiR72vG2qoLm73uhYqQAo5JM+wIq55Hfocl/eoq8G0vUi7QbEhrVNsjRs61BWd9J+lcJMj
2hmUy7I8QiImMwaUeSFkxy63XKV7fCb+0y6PvWSdWARsFzk1zpA4RE5ft6SdrcWjYg4jt9G3JPId
SWb1x4SFh/lPlc9MOnCaMHcFSj+5jJyKxfgnBMOMmNJAb39gVjBhsD+uYmhAN4wMpzVxQ0+4FZtQ
ij0OnBRmu97U6yYPRDFvuyyJRKE9yLPNQ8r59DhFku2fG4wB1eQi+tISTVPF9/Q6K7iuNGlqNQJ/
BddaPaJdcZO3dx5eBJSIlEt7Jy9dqah93F2h7TCtH9Vn7bBAckXQGcxKtY010fPijATzNbzNLmMC
BmjwXbK5/6rh+nC9BD9wZHmYwp0HLDaKCvNsizPyr9A3B0AH+g8pIaGolPhGIYcVD+kFCmBeq7Lw
57GgHLC71wcjI0oq8HuprpiKWMZDXQ6tLLgSWSQxdz6Hx/XA9eaf7a0bSJkNuR5gj/PzlHyVIv3Q
CJ6mvx1HsFyYWnBZM5SLpi0NgQqu5dppHTZEFlwTYp5iDoMJkAB3/xa6duSrcq9IpgWYVN1pI8qq
VyUaeuGqS5sjjudfodo0Wrqbv5c1Y3rOhG8i3OaNjlLI7ohvupmwe/FcahGPEvVZPlpfBiS+CaSb
CIgmo4TJRigxB3ihYzbSOJTgw9of8li1zx59vsbJVt9Hru8//SHhwbbbs6RjNMnPCVwsedLriooB
ZFvzBF/I0yNXCGWcUpy1gEJPbsm0a5OUWlzIUjmk0IxGR+HQUtHIORGAC6Qe78wscM7vv+X2FyQX
6n+SpnxuJkwqXttXhf3I7UaejgbCMNirVIUqu7sx0GiyNWYqVKQteZbo8+FNLSspUk2OStXYn7Wr
n5brJz62rna179WtY0OWzBA9Nl48xoY9OvzBuNze6byrRQV+WBc9DE9NTAhy6obo1mDSP3v7pNDY
+oe6D8A4n2dkZ9plsAOwGMjvfkomFXTCKX82u/DUP/igPlCxGaF8ipxEoFEtb+1Oog+AjWwDQ3RW
PLx9gnaOe1CqlzwsLKcB36xazVi1DcbX/3eaUwp2vfvWG4kESVEHa2aSTS+ArLRh7lQtWzLdlIwp
54anDmGTcx2I+5C5y0PIj5dZOb2gK4S5zEI4PVcONSRT0GLKuQo3dM7/c4QJTWE6ru2rr1WlVl9B
tXD661HHs1u82Q1u6yuruNeyOEpNtONVk9GhlPzinq8dEzV5mfF4nOLut8gfEAkOSlojo45ZoC60
dnX1dtUnHWfc53S/AMPa37SMOisX/s8trc+x20oLRXXuu96xwsdIQLgMJOn0xIgaNBrhCJmrBO3w
7ZXsDvdmvkUJ0CNHHrI+w7p4g8sqqAxkpsrUKZHLWWY37360ogEuid13XPqAuGlnvhg9UXNlTFw6
qiIGxtH4I9p1rPkpj2HzwO6d0k2meDvIRROy/lwACVkpnmhn8lwqC1538PPWgDknHesMXiOoCN4M
rzFSuxb1hbONxRqysFUQAWuf+TSU+MF7i7y0znpU/UCWttWwi/XKYjljukUTf1HNmc/aLXzMWyab
a51VoB8cfzfmSNA8XjCz0ZTYzJasLvsrWqt3unDjOv3S+PLKz3x0IOKjgayY0UKcDH0vpXcr3AoL
RhUMRuZpOVonAfhc5dWBWpJVdN/uL/Qbj+11STCL4ACAuoSQXUY9P1YTRH8QSUmmy8IlI+tqohHk
JnYt7Jzxkfdx6jjWAoOplfhuUDpjSbTtUZv/cQdxDYjT07wGus+MN8TNVxQFrcNAvKrEyE2w07XZ
s1KrIB49wI+FEBOW8KFHsLuOnfQSAyeh+hiQE9FUSFFGhbBoBmTPhaXiJXGo+kce4iF+07DP+Qf8
gjBAJLIgPQV19xed8Bna7ZGxw79oJCQIIQ4CsoevBRbHm/ubGFJlGXJirW0tnevsxi+YcbX6N3Xk
OuKL8CTMo7WX1wkwBu4O177D9dP9slAXfq8fe4InuQ8ABSw2we5eDOXGOK+twSSeO5wBsEPgrcLL
E9gINDRyNR2V7SEKEjBR2KUENv5ykAseF46+LR5v6XKau0kKifroscadhtOhybFMj0/En1HBzmvu
/Ee9rFIr14O1Fh4ThvNZOR/6ZALtPvLse/mz2O18fDzlYrc14gw9hKz9+PMZ9Z2Da3g6i9j8B9t8
yK1opyL2Vx9pKhCmwa7yAG/F0kc8GQqoKs/HXu2bizbgU/k0BmjgXXcCIFmc+izSw+ZXw96oESAI
pPpcMJ+KKq4YWGbR7SXRTutsO/lcNO10oi68eljGIZVSBRgYeAacHRURp11UWJ1aKceIrokbuuPL
Q6qpNprtcLtNc5wF+GqsySFqGYLohfNvZo6QBIXxODGbXHFkuYc85ghWKkRcfpzAhrnrEjnPL3v3
5YDOrgS+bxsqPV+0cgeB0+Qc0JqZtxJ3nOM/fWa8beANFEzVB01HI42oK0o+61Sa4H0KRCwHRpK1
xozlinj2swWUBDFqp1JsxZdxog2QKP6aAmiJfreWHNe3RyZ+8fXWF3zhYCt2Qp9BA2KMyxmoSDxd
khK1X0vEME+zeltsGzjS9bOkLw5bNx+j5Dna4ykC16RrhLnLaeCfZMZUL6W8Tr6WoaDPxxATsQgm
5HLHQrYyuvmV0qmk0uWi4MV6KAidTRuB1dQB3FNcqseXXnlIwTkeubct4YxyZIsHdAdoktt/QWq8
h1D92I0MESg3u+LIAm6ECtM7bzDe6HRvDfdDFWfsl7KPZ18VtfJMGVGlfhnLt3dkyArn+vrE8H/e
xOwp4rZagNgCUqrCymM/W+iu/O4FPoMYT8xzrOmxcKSN8/jd2MYTs5NF2nImAdX97gEE6+rlitdW
H8tYD+hqVQbQVGCOcxop5mFAu3L1aTWb9krlkxVB13R1fAFSTNbc8Mwcj+D5OGaRvAfrpQnCkUB1
j6DSM5iemmUkxWXpUjgiGsaLf0KNEsPU2GTmm6nkFLR6sF8+B1a42VVoJQ4jfbZpvH5VSQwnRgAJ
pm2QADg5b+upu3cvm5OnjyggzDazi8jeAjWx2vly5qJZsoi4l5WBQgU3RBNBk8YXUxv6N8tRg4/B
KPyLzqwzvBUzmstSkMeI6CNiUuBlQD6qrgBgzcYqBRCQ99u8XqsjBucQNZMDjbEf5kMlF+gNF1K7
0+JTbQG7dgJCm8NyWgwzhCx2HLz8QGLZprjxzqjwTeMuUqy8OC1E9H9L5aLpp1G7zYLrjU1ElfUL
SNw1oDPxXoFA6gSVOoX2dWGPXJSlcvQA3sg/pUJ4ugp+k4CC+KutdTrSzK4WgsMIJ9ezkqwENulG
OQD8WxTzU1qshp5P+l6aRCQmS8W76WJmGTBci7gi4vdVnzOu5zzuEoVpxTSrPOJk2UabXGuzZI8i
3plXnVrH7GIuUSt2VW3HNQgtOfq2AVg7WmYXsIy2TGe1OMHt/qNyyHS/fFmw1hlVqd2x0/CLagQQ
7+UBlOw2opMyEjIGGYV0vaWCD3raJm3ulJ+Wo4ZG92MRzv1yXsVBLID4sibyjlefjfWazshBNTsq
+0oRinPX1kgjpShLxB1wXaSm1CUdm0dzL+J6jh+ThiLUeLMOqcuVroyb5gBPh5f4AmE2hJvg9FO1
20RPoazVrbuq6no0PzaBPSQ6VRxg7W544IMscraTYSVuVkm8JM/E4lwnwFGahOZQlzJawZfW37+u
jCpXGCfQEeHgFbOXGy4NhOUQiAQotYYV0TSz1Aa40DAeSBn7ALYkljLoSKCPib+OZl3XEEgRYhph
j8k2FR2hW20i9YtxPo/0udmFsnjMPeSIzaVAOUm2AmAru4RwmWgJ3ihviaJ1+fDQQiGCDZRvk5Nc
IaHZutUan1EZ/GpqWo8zZhhugWowfbydFdmLPusDHViC28M+1KIGqCRANNqoyUm+cDKRlyHZ8k9P
/g1Ovu3rNov+m5ytYKVliWLpSv3O2d+2P80Q8shEBE6CzydWIiEl12miKyfM5+bNYHo3G1r869YH
tPcyy73bzOzOE8rNAhGV4EuxrZzXsOzwMbjxMfbYqXkpJy1y7lUF4ETfVRl8mKrmkV3X83gX2ARt
+qSbckRwSUiA6ULWkRiPAgTmR3mBt4XxKMvfG7fQb5eufDsV0J5yIYgoPu5tuv/EBywGRVABVrzY
gxdKLtNAFAp8rSIFTLwhtFbIqh6wfDO7lS/undfMt3ASs+zG9RHwcUFcqG8hbTOpSkQvqLjsDTxi
rCSQP+5dV1xEfTHjXWxfnf/k3r2rcWQ43upcUnUrdU+iaDQOCkEYQFU9Rsn2V4+a3ztYHpW7nIij
VWHte+c/PWADgB5+sGDtS5NRxvAop0q+R03eUEW8RzMA0WtZF2VoqCl/aqWkVGzpuR62erf7xq5l
S5CwmamfhHUJkuP5Q8gblkEt7zl7wF2+sAEdRoPAtKYz6S7dbojlVNJmEvUabX5I9sCB9AqOiozD
OqwwVikaZag/kCOfwRfyC1ADQPp7YLa2UBwtO0N8kBcMvfWGDzOimT5yEPuMJ63ZTFSC6ogKwBzw
LmgsdQrXVl2X00lBwd8kmBELIOamNbb4FhQngfiVbwU0CIpkhqvMVJDVhdafJD8LxkDSa+ZEBrB3
UixdNl0lTJZqQ0RyV4OP8BCgYlI0H/I99XuUBFg0lPX3wRmSXea6DUbkrbx2GsQiuwHcFcZAiFj5
7Qh422x0l5V6PuIPtOXIbw93IhSlsyQVz/H5rXSmOkSRm1pFUIKtosNWHDmi4wazjPGecjNQkSVS
XahQsH0nTwzmBGeW4Wau0O8boGppX+YmAMA9Yd5Cavg2Xx9EofBmFGnSTDSqqPIJSsDzAnXTsBDb
hBKDd1FmAK2uHllqpNSHBIbHpl0q+q1u2nJuXC/okv/+8CTkL5QQ4nXEdJyrSOEjptpmJn16aY3p
OtA/xUqFDCWa7yQ0eaMfP+3N2CBBpdkulTzj74kkjQsucbbtp4EV2QRtOVdaTGqkt9sBcE3K/fIY
fnOpEnI4oWeBZ6LnxS7c46vpQIxRbt24W5GELLXPFLGJi0ENcddeEymw5fE1LIqYCc+95T9H5tZf
kWVjufwzOJ7nKn/JjLFu89xnovGO/CauEaotZPXgCPxrB62lvrKvtr4pw8L4wGBSyVkwDOJ+cURs
VYr66pw/20IUCF/W2PggA8o2subq0oK0Zx2vcKPoF5kO3g19d3LT1eQfJF1qb1S8ccM6o7HT/Tc7
1+OwY0uVdIGfCctmLxPB8SH3+8QcV34HtMXdix7+pMaKCaDTKyfIvgw60O+JgU98YIwid8tf1yfD
BgY2yrHeRKXhPtszvZKCd7TXRcxqEZI/d6Q5heuOrRM0IDtcXkZGAm6IfA6DQat16zmTaiqk9G50
6wimWsDyMPmeRg99B2KuA58bqPr1w/8+QC3i2dMnXMwmLOz9cdb45zM5qsKTplk3cadnwbXaCHGs
BuAPCNf341OJ7evmpR1V11b2bODH5ew+uhvTHTU/aQvRhjYviaOxegHwWd4MPj+ZTHbC487GBPhJ
95qdiCZ6FobFBKcN3Kdmnrp5K/4BPgw8HTGvcPXjOArdBEWc2QzQscrf46FkR6ddZfFUIF5NRAZ7
fB92OyF2QZpZwPEgl25bkTg/higOsPnOSx9hsUhLhcW5I4diGXMlsKVgDkrsHywXwl/epj1j9g7C
QN7RGp8VoyRMD4c8eoEEjEH5cewujYzCF98+H7+1PvF+VSRpZLhH59VnxcoDRNjGW2nQvGVq5pIv
Le4G1+ffFDJNByH2oUCA6agAmgOzob+uu6jPf+qLcx5TGoZF66qxsm/+GBOWCizYByAMoW+1JtWN
IBhx0xNbz/5hGuX8rMQLFLcL5DY1b3hhzqDVE/FAc0DFerNDjYvv4BkyAdpPhn2LJCyyY2isVy8C
USXbji2dOwgoqX2LXbIp4A+cJvKTdg027oCbQ/4XbyrvVLcfGo2/OLOyHPqo9kDmtwOFPvZM3xh2
4gmZneHeYV2i5I7D/V1xZmhKA/M065mnVNqKES9/HxeEhDSuBzVoeSUPpV7sGJXamq4EVEA1t4FM
9LG5C092SkS3WW7B1jStgZVqxILnj3D96nzv3bpdQHMLtKnEFVxVIAviVxCs+mDT+vFgie17u0u5
98AlVHS2A8FLNqatW0/5vErvt0rgwOSRfZ2GnemQKbTJfIg0O2wCxF3V6deWYLBi1D2ajbJi41Kp
Yb7vHnBFnMy2NvHVfwV/c7XO/5oQcltknq69ftdkPWT0PiEu/efKt4rHdgTdcpIMV2xRS9u2WXJK
LKlCUF4FWlTHOtnis+3Dz5yxMS+JkrZ/8ADhZtzwo3bNNQ9y017PimeuIOwxdg/2k1cVZyKjtzMH
S/raP4LS7KIA7coz9+8jjk9vzw2HaLz38/sgg8ENePs4jfF7fwkh7bxUIymLnLBQMADtnGTZ9XBz
mLzFqaQnBjnwx7lcFeaujS2WFLu4N3plpqKQeqNDi4iz/WkCBvGnkRFOxGj+5/YD2vd7Utsrbpi5
LjgeJDihxocUTexelcEIKLd3NWuF4OZ2SuN3yziBW5VjtejVT1DVvyS0+hNNYtfGTdU7b7ce67xG
kKKpv5qyGwjRaHVC7HkNeKSmUMm/uwaxknrmqBtO2ZpcaMNiXu+GjzvxJ0JGDpykuREGunrbjdB2
H01Uo6WLZRCYNd1iDuoA7WYmWP72zu9ticPAKfRa6OIyFw74ayPv73oGL5iln9aDg7K8J9qHqKbj
DjAxtwRB7kOWkuFB2PhdUzeh+GW3mKroECA9V+jtDs/IKOk/SmGXo84wH8X/CuUAvXjDDFiztmDW
rBRRA9JSHe90Bhw0XDWaJlf2ABqkZylJO9cj0/Ke083NJINlPwJtMcJQOMjmFfpQ3ftynX/4++SO
gMSuLjHLzREyeLBK96HnP7uOACJQ/IRmtwNsm4Ukkoph1Wdu0gkVHU6e31rVxHI8ruZO/SmH8zGo
IsOW76kuL561hNDIVI740fhXenB+oOqgNRhbC1kqdYFKkUzFdgd5LQUBeGJaiOj5STFifERJ5rZm
gCZfomFBq19pymDV8R4mAQdK//oU13c3hqyuwT+EmegLEw83U0BnnQzdjnZcx7Sb3kISfMtMfaLq
NUBVDqtXZMYx6apaoMvZCLna9LqKj8/DBSXQP3fG3U/yDFKhE9cJ/MwP0TACy+tsImWK9H0kSrG/
dCLEnsNIQNeVMc+wd8KfAlkObCYdZ6OviUM2vzt6hP8y5RpnsLFIfs7GwTgWmMMRhdJaH8Yf87Il
Kxzc7TYrtO7OcFpzOBzT1bUBlzYgqB+YR29LzZYYRDRGKNyBoQIOw/u7UyMPUTAChsDYSwwvd1vD
xyzCPl8lIyA89wnwHDuYsZ8FlH1/5W6oQ1GqqNku+Ni6rjrIr9Tqe9PPtdnpqBGEkw7fguNnRlkw
bf83cxbkP4aEVDN3o2Vf88WbSXju2wbDLwgmNPUTMBPiHs8VbyjiwJtoMjsJnbjMR9kWs3AVf7gZ
XuTdZd2dwHR+wfOFls6XeqvCm42lbV8eQEhEZlmYsCOmUslfPcF6O9K7XKbnMI6ZLi/R/WSmXnGF
74Kh5f2XD1BrM0I+oS6RTeJb/4UPAx+ixjOklc7Aqm6EnMdv2TzOkmzkIYvemwtqCC4rLdLjkXHl
YAcoNoowsLt4fuIR8ytY9ApOyF9lcQ9UCwGrW+vS3KiE+bwqSJ7RYwns5iNaKxHv6QTdVvTaeUiQ
cJTADwgL95mogxCyaRJTXePJiYS6SkDbhEvk4wgSl7lh7f8Hd2STP1M2Y4DIIqQ38sOI2ZAbzHVR
6FCw3bU4/DWfr1PKn05QLhHcg/8Srwgir0fnuXejlfNSViT9y4MxtOkbmjbEZjigQIkTBZezuaAQ
w0LOJyOSpIlHl26LpEZeFfi7ytdZ0rJ/90lfdJ34kSKkOEmI26RBNJ/1lLAQUdINyktF/jWs0Bbe
Kgw7bXL6XtUY2p7iPtYpIzB513+1Rb/8Vqj1e6AbJWmB7QtmSHk3W1YDwHdcaF1pOVIGsTD25tTN
Rk7U1J9SnWTcHR5wcpEAn4n4PuJk+CCAP/7WiQNbrzUhWewLY9yvXcm0FB/b/sc0AsDwGfad1X5F
DXotXKXiXafeg0SiZxbfmu14Zl63zAXVmCcgWQ/J/D5d26O7yF/PRj2ggcku3jKJ6+H/HESnkCGt
5z6YXmfiW1fGqxVkYE2zqGTcExz1HPoUlnQmcA3LXNAXvZ9WRxAboWwFp8nb30mssjKQsmln2TcM
BKudu8KrBNEo70iBaDJqtLDjvGFd3WHPP/UBFESEjcQ31j+E56CXpov0pUAGVERv8cQGdP7MBNY6
ctBVcCcHeLC3O5EiIvvYmHZgLgW0tUiSJ94AwAI6bfSMl4ex2h+n5yaB+xx1TwwEw0q4c6u8HN1C
dFo6WoimGLRCjhNLaghSQo8i10pYWTq4qq8kN6Gx2IB9XL+Uzzf1vTGBhEwicZMjVJjmB1TwLwp2
nbraX9MgMaKkpgEnFR09F80GknYl/IvSJr1zMk8Ykaqs+YvKbZ7qKguOpg8AV5pDO1Hz4JJkjRan
LgwjpoFakIPdo09SLxQebtCuQi9NX8H1UsK0wkQ0DHl/JqN2CiGz0veLJQ8zWijlbYKgjVFMzhyc
sGNwxXcFzi8qlQ8FR/kjTRydJAiGlUmLg6fT9VNPlu0mk69GEnYS8CmVgNtIIRqfa+4AauUdomhw
NNnI4spcH+Tw8jo0TkFxDAzSQy4pi/+fTjwkCVORhp8PKI2/2xX0BYb+KyvrgthCqAcYg9UScBtt
XnLFJdEeFIvAZcrlSeHnnYMRiYouMxjKj+oSG/XUCLAu9SpDv/5IH3u/554dbAkO3eEmCMfL3WiS
3Thw/mP+KL24SzSRI6zqX985m1nvUeq2a2K7qZLYFiwNLjbhas3OlYlKMy047Q2P2E+x2FIgJkiN
/faiKCEdGTOsv3EpWBrcBZ7ChRviDK3FY8oBXQP5XMothu3cXUp1zGRNts2xQ3XxkgDFTBhRkXJa
BO55SNKUhScULUiXBVrBLLkRytXirA/3DdyVlRMXr1kOGa/RU9Yn3WwUMtI1c7xAv6Lqf68QwhlU
kgOfdy2E9is3aUT1UBtg+ZSCONx4Hwc5Ii9aj0VttIC9GGhtlTOAIW+3xn0xZjSimPDgv8OVyIyu
Ik0OVZcK2SojPWjY3QDvCSP2CbejzkDsbL+PcjVeLQbU5uZAMnLh1pI+dnQFlqTMB37fqS2ILMu5
BDDskKfe7u4xcadXF8OrrU5KFRKQMVN2vYcNLn22914E1pAVGgPbRbfVrLQpNqJHD82Kwpu10qVR
yiPhYUHlrl9uOACY7mvErI6Y/yiuU2mDmIw3EdCWYFGBbfXz435igGu7JsHrAI/o7rouvM+c/CHq
d0HiKfEX93oPWnF5j5QEisrL92UFmrPzuTiFM5i0WhlysC+Zshz8Mf7BV087dyqTP57mJKBFkDlH
MQ5bSL0Ous95c2JyhJDNee1qfdZ56d2+cEVvDOr8DPmercIsYD4pZdNLKWvABT1FtZuTJ0GGnQn7
zdMrerw3+5Mn5gfCt3kOKeDA4liqZNypaBGns0aiBVHrXV3xzBHIq4XkjFvZLU0lQhwEhl9RVzQY
yuqMqrtaaSq8IrmzbEnARswz9BwP2gJf9e0Ly75fzUOKPM3zlQYruStUguV+Lj2O+er6+rd7ovpi
2LuuNNCcStV3soufS/KBCOfppU5IA+zwL6CUb3J2WLkpayGrFcyFb9MhMyPcypknZAO2DGWAJb+I
Ng2vi0YEjj8zvkiAQ9m36KlCVjbY71xUkim1VO0VCLOCMVSSyo9+Kwpp95uzWzOfos+FnOpt8tjr
YicSG8YzY9dY300WHD+WElwmps4Ywt8WYYkuTDKy17a5yYyPAXllxwBAKnsIBt+nb/tFupw0z2Mh
avrp/4aSGIHyXBeFk0Ud5Wbvx2uyzsXCpoYu4UiTJlnb+6LVHwjxpxntxveiIgMdTU9UCQDxCnKP
k5Svnxi3ywYB4vufihdg1FdI064FoFCrQrBWv4KeAwnWD54h51uAPK1iQGpMCCosb8fji7+nVaJ2
C0Y56oxm1CzTu69Wu+1SOXo/x1cudOVaK1rZYzWm7Wqc7H8MCwOKGVgnampUjxAHwnxvsToIN26p
CUgXLiA0khFLiXPj37ZHXzsYGdBxajaIiC58ZUIpHjj/Sa3oHxphvQPPssVOp48KI4rcZKq5z7Zm
uuuJuqjdb1rY0KcL2SVqXwmZHrNdQ1iyL6TfXPnzu071EdLrakQ/Rqu5RGkIqEHe9D1jYVoCZU/B
iVQdAnJTDYkXGMeF06uJnA3bUIyqp6StrKrZDj8GzTviylwoyDYzfj5gY2YcNU1h993kpd8N6RF2
/uFq4qJMrbeVt/ESWWT5Ij5xEymTwV9fW8e9xCqMqcIPGIAvguliZz6kjpzsAtGIydhXuPfSfKHv
BCURdWnFYSOPfWhehZnnGUxh4LusbFZGJCtlGF3CgzTRG6BaQdsOOJ4fcfv3Q4sF/4m5xhwazELA
11C8lgjvi4QnkVTeG1g//hGkCG28iAuauTFtYoB5vj8CPF/DBHY961RzSjkWZEOFFx5MXqPhCthf
UXN4bbJmII3kTRY3qSs3zjtutzz1MfRoem8mEiWZKWiXcnX8xPWzXAcnNhXD/BH97KY81ufyXj2D
8I0+QvGFhd2L8dEKUDzvdS9r894S2ImsvY5f4PhpVbkWasCqeC9O7BHg2+//mdGfK7MQcSwR6zQL
F0E4nGDWxzHUWV34Wbg8mwiDGBMKCuBS1Tn2FuFcKcjKgfugmGPgxiCvB+rDR7tsVHWyY7gbWk9r
r0ObtVe+6wt9ZbjLKPXxi+Q8+CXWZdyGpD2E4wi7HbWN3xoEvEIMk+wNWA6pYNF+EIMm4PU/a+Tt
SLH+txYKaPJH8joJqht9JLxag8yN7m9Gkvy6MlxICy2b/wFl3PYmAeve8IuNmt1wC49wF/nPnpmy
0aGP89/nvS25IhFfriX6NwQ0Bu4DXYpZZ299fF7SIU8nje41uFI9R4oppAotCh8ZLVBG+XjZAd3H
LbIFIVw1QP7cDFO4hwv2YeDLdmLo1FEamxEqtxoHPPwMDy6FfL/qSGmGLIbiE31F0p9llX9P+8Px
yFW51XsK9pluHsLafXADOrKaSDdQDY0/UE0ByolpCnaE+g3Wwyq4DoRPxPa6Y/Mw14DWHr1KGx42
qS2HrqyOp1AM9mEuE+Cv8aJ4Y6DCfeozPq6vWkIRWgVOXttBHsRsJnsUwsw3X5U7Zjj24WLX3SUG
whBS8bLhQjClWjSvcOMgtRmAodk1006f5Fod3r+pGWgdQ8sRMzPX7zP33Z1zoLHls19Ls6uGkg3c
HISiOAjfYntO2dZQ7BHtb7CFmb0c+r/HACL/7euIGjAsziQXQZsPnAMJLGpl0DkBuJi6jmpPfkaH
ch3pgnHbW6WoW32NJ9GXawwmr8E8bbc6vLZg+NY6z3yN3hUJkGq7Rlx3NFQbtLQkAlkHV6TrHqYr
GqsFL71V/q7jaqIekGM+/1khYWIQM6ZzPl9fsEdzk3F5Rr7KFDDWPsUBWmBjv6R+sEeVgyzP3/00
YO1cMZlPWW9sfBrEAC0/JJR9uAZV+CrZ2587n/N6cbGw+sFHfxIW2WPJs2y5MbajUwTTCKBkT2sC
/KPEBoXhXnp67Vw9x6se8AWyeJq+2qe1DZxq/K8Mtftg49/GoT0EDSLXEB4Apuoh/RfJsA26vbaq
JtxsyVjT9kjJVGozu6CrG2PuVMbNtvZnsKxbp5U2ZZVzU0aCG5xaNbTzUjkF6ZvTcL/a/Z5BlMyw
9Za9LoEJWTJEn7nR4sqkFicSmXAdn0g0RmYNEMEJmv9x+Rqwq+201DWWPcj4W1w/TYToLtO1iu0i
NRSWTsLYJh4O8Frza65uPFOAN4Oua5ZNTLqKkmqz51Qz7+i8wRgE5NuSEA526+PGK2zkzkNbrR2l
2IHAvwS7b9wuEFkKCRfw2J5JmfbnA7bFjp6yf5Rwi75dBO3unRHw/JQEsGa6FJ4TMtxRVf+ejIPc
4F0QUwd+2iYmIWfPWB46CEUwZ2uTJ9zqwy4GisU99lKAs0M/DWUrIyOvJ2nxSMvsbJ8szXXD+Nc5
7IlATgpfyu9qkUN+UleSEUQJsaBtnJAt2OuJOmQAcBmA1g2nfv8vTaCG3WEm28cGGBJsy6jUD/wU
yqTn5hZnr0B1gv++vO7wtxUyJDK641VCd5dIXPo8bWlI8I65dHA4k/c6KreLL3wnlmMWOIxvqIsc
yqT6PmC2P5RH6mFt4aJnX7a6ykx066MGHnAK6lT2MiyOqA7Efp9RMNF9tE7tuh/SRf/Zy0yrOFQg
njmLyYXQx1AQCGcAE4hGFC0njXjKKNQWJFzR+XKKHuKo6+XSFvauqGaiOk0fQHxt2o1hh9p2nht/
dM3/YW4ploaNAedCmlNlLutTNtfLJ3nSnnIn63RAgbA2vOOonj6Plwj+ipQ1H091Rx1ZIVcikYeP
+Ior+2E8U3K+AKTmQurEVS18/oBiaU4YDoJGvmnWPp7x26k8YCu3mRD8j90/wfu79gudIfRm+31r
M4ZWQ/ysD0xWgNsDCVpYMXgswQdtoYBtUfwnkcT5Excq5ZeNxHim+9mXHhKWX+JkvT7thpvVoE5L
dpVSdOB4ngKRmcX2CSigkkrn+jeHO05yREGNtcJaagKIvz3eVdqvjrG70BK8FCDWm5MrZysYfIFn
pTM6SnDtHVz8WGnqbS1cpvhPVqa+SUPud2ugADupspFGnnZkQ+yLlLrYfdMTsX9Kg7/AtIy6XHQy
035QMRvLYeSftqM00mL2BfiSvAmULW2gW3D2i3c15g0iOdveAx0bUwsUu0ohSDvJPjdYCc0pFoQ4
ely4qrlHd/yQNhLQYvWefv/vpFBIYz92E7ztRFLPjpllG7ph/a+wJL3N5YwT1utnjr4DWh5sAZMq
t7ZYvhOeLqNNaiuElzsfjWE9LL8Weet9laDmMNNgwbBsTQqjAw6SuB0ScPJwzSspFq5dWoXnNjsb
J4YQg8u9lUxEiFmXK5/vRuzzCDVObUsanDoCLsnLsqZGgxJtYvb33FVOb1sedL7XOyL0Fco5b9nx
3mAj36+wJz1sd547lVtwiKxAkW8oZLk+ch6KGE5oKDzvG2+GPRDPVW3M35vxwTL7N3P17i0lg9iv
uJl0jptjGozSo5jA4m4S48q26DBftxxtRiztsmt1ZeO4Z4g/bK8miRx/Jrzw03g1ezEwmh5p4lmg
wxYxrnutey6kwYgnHnqOhbyIsIWha5m/Ty7WpdRAkENXywHoYbNqj+wTkiMrQ8dTaljcqRQXozu6
KyU62bTV2faSv2Onf6gmu3xpnnu/voFH4HK/lJ57CbZsmMXRouSc4RngvyvFcaP/umx+QkoSXyxK
bZzWpKc8J9L8AXOztZHCjKawm8mxgkbiy3+rzxR2GxxAelwMNfCtj74HPLeFkhhq1eQr8UIZn6kF
IwornwO0xXXkJH+piVF34eTgjFvA1XIxpkdM4tIh0SYhx02XqLO1cQL78wXx+z1AkOo3UozjkAvI
WLH74ojXR70SWSGxmvSs86iFGTVWmqhaIN2P7SWod3BeQ6onum4MaTIbbujMM1ixTaaEA6DbZzuP
bE20stxLEuc3VhxhYPWoO1m62dEbY/0VFNe7hv/hlftEvCMxp3O7xVLnqyzKTOy9ehDCREYjrHsL
rbFbFQzrkq+Zu+DIhOiMzAo05s1qJMsY6NS0w22kB/8z1qcSXsyChXLs4kYWxxjFjKCfseVcC04T
LsFR2UDxA1PkFVs09+4rzC8RnC13XU1vC5T687p90hVcVS7SFHFa5B/sPkBoqnQkILBQbbcdcXDh
4L1D7Tt3qmFZkAe0PEq7TbmmeMva+yhEw/igami8wBHIBh9npgz1Wpb9lInn7wsbIhbvfioWej7p
awZWHZcKL0C8V4PlN4I/kY0uwzBbSSlQltZAHhMtggFmOfXbHiKdMwlprMGDkv18kxsuMMDp1qrg
1DX2TyJs7aVjiVhqTk8PHzuSzut8sqrJF/r4YUYpbcxOs+3EbtYvUhsWxt9FX42cxdmP7V3bIvit
L0eoLlN1potaKlWuf5kLCMnJv1ACFc2SAMpmEbzSQG5K2U0o/qAvURy6cbS74UUFtgg391Px+gRY
AETQkcs3g/KWd9GniuGItBQVQGso8ZBHMmXb9YVeix3Yd3w75CNsqgdbeIS05rjJnzzYP7khp4p1
BV4hrOOSPqtqS0AI2EloK/WslZavcXuV8Ms3iJcVB5o93Sw+k6RZ+JTYeWCk95MdxKO1hH1nqK5C
unel2sK/ahDKnJcC5M7hjZ9YcACkDy+ZRTym4fdPn8KclxAmR0jRePjCg4gDVRkO24TlYsKI70Iq
0qYlh6ql5bh6MkGQx2qRMpTldS0Z+Im95QrjLNvoQMnxaKxS3p+COkE9jQ1BHXuqNLbJ12bTCsB8
QaNdOgD6b/AeOj7FKtTp/YI2jSRVZlXsA2gbPo6hXCftDLYg2q+wRlCIo4b0evYy6OoluGEwNz4H
2iC4gm2mO/nqndU6MkcNMh9LbSvCFP3lJZ7b3Np8mXRQKZUciq6BxHCbTXywgdcGHMlW2dhgF3wU
5uAFgSnLrLeFze46kAvpxXVufd0MnTxFxBhakYrocfXOKEGiSF7cC+yztzlFZQ47BDK7mmfCBVLc
58MAu0vzCbUph7HwXrl4/AMHaRBa9vHWZpSGgzk0lnpiLv759qGhjisp1rktkUwDvoGHkvIKCBQ6
nBEAVgkc/U7ncNDPBfdB9pYiGQ+5KIuIf8Unz8xmz3MYVWbn0TThFKuEZvCAV3AtROjM1zteBCcH
ZQnn5E5rE9v120tL5nwbN6TMEKOSGrm2xF34R1Jw6GFy9CY46h8VoQmtz0e3egNLMZglvUq7ut0k
5AMmDMLQRwEt/ozyaDcMK3QMhYfMCHe5/a4QlwND/aF5fa6qSq5bR0HxD/amrJ7w1Ysvb8EE6jRN
lqozWmmAX1Rv0HDMN++VNN1m7nKjDoYibfVCUbxLPpvDB5L/i6a4+9wIzNndgSgpTeHYzlt29GRA
EoPfdRBwA/C/+2d2RYpyDF2XV31tqIEiC0a9MNqCNAT7SoKmx15NBAIyFFmndGz3pmfiIK/sM1h/
O86Q7WXBDhNmuj6DB6QuVqXpg7FPqYjSMJC8qQCpsCacRuS6gWbT2QDm4JmB/gwWAVWscLJXdsRP
LjnMvwEE/MeL9ZaTufagpoiflqsgEz3BkNFejFUq4563YwGkQUTB+KsrJt90v0tq+oFb45N4JNWQ
TRIFC/r/o378t7wjNq/S0K33MJMAMy2zOC7XQW/nMsys/ndm+m2nOesx3Y8xRX2/YNXlRPqCpt/I
mwwXVcEKIbvsv9kLSWYdHb/GgLR7i3TYdez98DeQpdPmkRHz9sA9eKKdrmeAAkyuLo/Oyi+mZEkF
OR/iKyluWgV3EFTtPD42DSyV0HNURVfzJvNG/BK0lbbzbHgghdljjm7kzGrEPyj07xtULSMogy4R
N4Z1YWszf8GFS4vJxHzJ8TLdmvpmo9Oj+4E65villj6WQpJxukRHPPaloA6HdPMArT5UPBHmbuku
gyrgJcHkUON28JWanwSzz3mDkD3Tt3ODKrZq2y2oKj7T3tKQKreMzl0e8q3wvxklxHa4nRuZLoaz
SuCW5e1HNRQeojxBYjmA05F0xAH/yhr9CLPOdcUvRTHwWjwVyOVTLSji94rMh0yXPPtaCSLWeCxm
V1o/fIGUmYkKq0pNPT8LLeN9t/lOLljBSoEL+DsLsf5rvIpcQuYDwtbZxspxYI7gwvVYDrj82BJh
UWH+HkYT+JgWUdxF/N/KXKJjuejM3DvuZm0wMkM/UN6vYqMIGzWwY4NMuOIxNMO6Bmq4n/jLPwo7
pleE1RbS8JgmEBjGI9wGEVDYgwjY7LRpkdofDEMnIioWifqfxDis4F4ef1lzcRFsaexicfHEuN/I
rOkwdUFAY9jUMWBzRBtY+WUHHkc/idJLCV6rerUZl7osopQyxLhVX3r/aSPUhfis79iU+4gWfGlK
7LR3n7o5sxH4lC4Zq8cvKpNVO1fug7paRh6z3O836FsFt4eyB4vSYQr4midGq99D1Fs41EAAQ96G
RVcRNUiOvJNuN7aUpQ4qU5PbYlIgZGkrf1+61rX7vxErI0Sw0shQ5syBzaFg1DA3v5NNqLkNkI9p
BBW344vQkW4GaYvUmD0csNTGQaZ+niwlP6Y2EEgLZX/ija3TgfrJUV/OquVXNfFmSwHkjBrdnqp6
TkG/Hmxb+RP33KRtijVsyG1RFfkLLekOJ9YloDmtOAzyJWZudOmJ3+blw1lzNC4AqKxhGdndhlUW
HK0NFlcO6E6mX7TpAl22AjG2OoozB3vsc2H6tbvg+jZ2Z5fdL6x4jfVopSQ7QMgSsyHnmg/qFvRC
Ed5hUf12//veKOlmRsvbqjEvXTrO41mUL+Cc4iCsZT9kNKWQAPQ+zETSYM9FSZHuEeWQIXlk2+56
l3NyV2wvvN9T89HwFusrWB5iDAAiSnBT0eOYa20yepIWaRaVmYMNfoUc6zCsXp03XMIkbwETJu/9
mfcGB6kszhfTMoIWu0ECYfyvFhtvVbCaakErnl12CROZ3tMA5HpNZvkSwXHF3LjqG8Vc7hr0CTIm
IgS27lI0Z5B09aZ/CF/ORYAdK12KjUHnxmNtETlB6a5t8HnbYWziGLWvhxmqsDthLaqAJKCcP7Xr
T265YzBZbaG3H+DmUvDVdUFc1s51EeuzDUh5c454UsNp+54p0DZ63lfsRa35ksYha5Po8SpaRsEX
B5uqz7+VrNeCSqyKqn7NAHMk8OGQSal/sOQhM1T8pOXZUQekDK4nNETzmRYSFvUTwKtAVppVCh7P
YCT7UQlmnzZlDGHBc+2MC7kaDIFUPZo04gdu1a/mWPVB5ftOodyL9G5osfZEcr7H5VRWwcPvGSIp
giLmxKAxC7mMzVB6h0Y7i/xfb4xH6K/gwhoE4ZHBlr/7q4SNUmrYJIGoaF+3JE4kkPmJGwO4inlu
oolPBeGLB8UknjV5o3HfGs8vqlPUJLFMadnRg4uYsk2iCblRxaWsaD4JfRCgI7a/mcJgHdrkpWf1
FKKLcoGuabeE6ORQVuZQrSBXOPbTHn4/d/PK6SlgyZMkMcMre9IoGzNO4q8/zsi3xO9wLfLBXVpH
rLSjXZ3ZFvL7YeCTP6gFW85V2RNK1v1JHEWgIRavPZIqlndwySe2M2t5u8srGcQIAUtlkw7gsnSL
UKW3kkuiRn+bSZ7vXByo/mjmO/HHzaQPcHbSCxYdxxhVPoVDd8tyeFojrWtHN7iXuSwQhLzgmGzS
YC887JEV/sdfMVwZiQUgFnQ/lKofesOxdw53pzYO7w1swxFkoFoRJRI8VfP5AZqrInDb9WPKfKdp
AsX8smNkzlRbC0Gh3ZVY1b5B51DIb5JFFMfIITZnO977qjajfxM87Z0YN9FoeBQT6+z7Ylh2fNVO
5u2RWvyxM5nKLlIwB9/zfIV2d2DOkrfV2BGh5fJ4BXt8Bc1CIxD81LxC+9fli9nUlrav8t95W67X
L2HWn6tnaS6UlWjjfIGZU2j0YGovCVd3PzG5QL5l8UoVauORFkkUvrcwJcvWPy/fJXjCjxXTASmQ
UITYueVuC81v+I4rNZO9UM1ciPoMdeexprASdyRu3YeAXg6WFc+YTmmMlImDAIDg+fUiVpQliRpL
ifmWLVrJORxDqA638UxfryPF3C18CDurPQHby9JnBHkSRixB2DRpZE5kC8ARZFYetbQK2Z4uX3lA
VXlSXJOwqiNLQPBUiQpyAqmCcGmKLh7lfK5Js16mMXrYysXFksby/tVDuFJHzvKiEdEPQ1KqsRFH
2W1d202CR4EWcjGP7CN0qPomgR8OeoQD+xLbeOw0St4SauX/4caBht0wPXU9HZC8koLc56MSluyP
huoRJlDxWyVlNMVO+5v9DgD8ZOYXmWozJbv8h56RR616TAeMpdeE2dCMnD74bUCImBVlbNrT5ffM
NXMUjs1UYtiSvWVeVwM8/x/6WzVON5tQcob5j9n9FakBvXBD+07V2eqoUGJMvMHZK4zkSUpq94jb
L9KoTa9d3kESBAkuJDPi0Uk6FoLQ4onpp5fbuPpEKdNe/wl0z9j27sXeHbA39fwiBJ13BAGJgdCo
bnddAxPjf8NRimAA0Yvz/PTA3WVcCG82OxnG/7AtM42O6VoW5GbB/AQs/kbSTuH5dJxt63J9ucOe
r9Vm8+T10tj+MkdZG3KnEumRjAQtWvDIKyIXK4PlBUg8jzaFQ9gLvfd0yTEJ+AoqiJqa71Vee8pc
A+zYR42Mm7csBN3aEWKGTyIjQXHOm4M8TczWrJrMQ0Atl5ZqRnWRaqfZhpYn5X3dvAQLwK35KsJt
ECSSy1273gj5pqXg+vtBKng9QmkOpLZOmdX/51HG0hHxZ6956etp/v7jOFFoU2gSNBbCyyDFHFRB
qg2ixi9WJv8Ean+MXVnEiQPnQPIaV2ULW9dXhgeTd/iJh61lEIUncv63hmkiLo2B60VmKSu7HKEl
AY5VR9EZE1QN6p6LUGLj3Wtd4ZMH6krPQth+iuyeCyDoZl+bxsTk2bx3qfBGWf+ZSIJNpG0vIadY
WLcyaHKC6SGUBow0KbU5/FL3H0UsikB8AN/DvRuJQMlZXQzNa5r6LYoGdkp8pB4midnyldb6iEw6
6FrpdZEYPtOXPBcHrr7fD3pn1Pt14fUJldLU8t6E9Jc1YpqG1Y5JuAMXgfKoO2aL5Vy8EKLLHdzj
MFOTuPJjL8/zgN3KOb9Id1snnT9IRQ1vnvJHeOp6C4CHbc/zlEXYvS3l3HjCwG4+nSFSkh4tc5JG
tugG5bYSLFCRv4zaAT1ecMWkSIS6e+sBcfyxxqTiTcZFa24YnQWuu30qKoNo22MGWce5LfO/qk8G
tlS/Kk17y7P2yaLCvB6BXxmvymP70E8w4+He3BGw0PU1Cu2LbBToP5De76JZjGibp3R5JjQC+5sc
/iP0ny8fqGPZSs4LdpYxaSNTiNqlVfgN6+JYz5l83bqb5RrzbaXU2UWHzs+g0MLgTHGNm7ApdJXs
Y1n36MrQ6Z04v3y9k0InQRAxWpKEftAeKtn0o/DOWORmqNyaNShR/e7VzD5B4K4ofDlUqQGIRqNR
poCFpErLIukONy4f3oheksZxWOi1jrKrl4TtgpZZv7cesLvgdQDUVSfDsrbGm+1jYvBib4uHWDZU
ibSKm8R1SDPfWNAcHqEBzfdZOs5TXyNnE8j8CG2hkvOPtoovGOqKUv0U46x5AKHatTcTkOfdetNt
RmTHmrnizOzD8Slitl4cogJIQ2mwyhdQsQAzvkXqEl6fyZTlZ1KtMZcdy9KnZv+snFXif48nUTm4
cg6v0+mJmCl4025xpQ1M1yozfpGUg4r/QwQLD4XkIghTKnU1wAn9dQAz0fLZqslNmlY8p9laH9LW
fruWVaG7fIfhIv08cqLs0pWLuOFU12Y1kV6FGdweVCkxv8d1mnKIHGpuX8GOK1+gIGf4nGk+yThu
Cv10Brd+KlqBAx7SzIC7SZqA1GnhzFogMu9lCwIQXjK6DdnVsswdbh3tj9d3Sksjzmi4FuDHrWOe
7x0bSH01vkeEMuOIn0FyvwN40rt15JEbnxMFc5EIrOYZURjoac7p+4xKAuufmJJqznw20eCp6quY
WWqyVPm2ccmNp/1te0Xrn8KuogtN/bqe0JvAQ21OqZR6cjB6J/2r95rmznJUqQ6hksZf/p+gpn3h
YbcLjTNRljNRc1ACGdzONveA2qOsfeSymBHtfJofMEBQ0x/uf0NVgQryl5UmYGrSTt5aAs7iPJ5x
5Nwq+i2v+75DQ7l4lZOvkjuZstzarHnqGG641U6qcz6wMXfsgw8EESK34Ts9In5M6QXo5tL4Xq3Y
CIlk00roh8VTdRi0N+CqKKXw7bSJ3Xaq7gg9nhSDd2ROfs77/zy72dV/RITUfBU639tgSgjFdmob
zhcjFP8es1wF8PE+n2+Z1tAbY1PbwhZ5PeWltWdbM53iDYZu6Zc7vHNC+ykhvzTqrFxUu61NU36T
KrXYxCR7RNFu0S4YWu9fcP8ZKDxqXErdlkm5E3C6xufGUUQ167p70ExQOulhWUbFcHWykq9/KliF
fp6oz2Js79/s9qkJLbDgnePpgAW/B2FB/eEpwVyO4xBIP2MBgMPDtMw8BcrtNMpLB0UCqrq7ApX5
NFTxg8u/MruMjmiJ2f+UUO4P9wMbH/JBWs+YUwZ0x3SD2/J1v+Sj0OrBfPg1TF3YwrNTVhy8e1uk
8bKfHQbHhBvotVRSsvPPYbrQJYPLC3IKAHa0qX5SVmnX/WyvkjRA9vyO9KBsCu4orcCew169jRo+
AHtGy32RJd8vcv03INpF/dqrijhjpVr+L4oV1kOzS96PnIEl8ZzKBNJHm6I4VCTUn8sdw8ZTJDAl
sRQ3CUGWEeQ1Xreaqmfbi9r3/kRBpSVsBtup1n3IbE4WEWwOhMMW9oy1RMnkF0P1N7YvSFBpgXOw
GH6FMR9cG/nH1EgRf8PS5uLMGKSQL/8/+yhtcFSeRsAeRUcjzaAxfaAEzvY0CJ0WpBMw5MT6oM7p
FvT/NWoyIaoy/SmBAeTovjfvYo/CxSD54aQ/ipkcAK/d+7RDvHr2hN9Iz8grfyqXhG9XzJ7LnGln
ePyeihMywKghYy+bAkBRjy2dhQlMAJsnzw8cTF0cjn3/RMrCjq8KjwrYYRZRPZF1CWkIXaAB98KS
yf2iVzwi37eP5kry/eRqI14y/5CG9dGw0hPp6fs3b4tFloTFqfqCwD2fNHyGL4ZLQyE5Lhibuj/d
Sj0MwVqtRgp1QkUumIV3tNWJe6ZxxDg21hMg+sd/9RffP6SVWVMw4od2R+3mTmUfACHLQmcpf0M9
xRPLAxCgZftF68QzIonh5dfZq8y0GhkiXVV+IWEicOu1Q8Zt/qgLTpHglUMRLip0cKHMIu4FqgW1
IOHrANyW8vJ9KfwyNsJdxqOWvOgIU/dy3kUBnGX3oQcg/FuyZziyVEUcwsp/IKDCJx1u31ku1DOY
EYrIYW4Ksls/0qIpsu13F1ZTk/hGR4nxsir2GjqJMK/StJTYwkX7hUvQ/inPW5YwjwgvVup2MD+h
LyJxZV8cRBaF+xGypU29WU4Qo1XOXLXnz/UexsjNyhdUiH64P/6lIBQrwA+BCCosuC33bWi+jT3M
k/BMFqFp4W9TreoRw63V7kCyHxQBoGKNj7LltaQsQYVdAN5OutPbiV2cEJbJEyOXx6+1F++oqAHe
6Ek233MqNKfE50m+5i9H1JV7eT3vTmI31amA0KCrKNO8BMF+3UwN1CiZo7w4iiBJ7frwsgcWI46i
XAT5P0cKcOleZMzudQEWA11iDEEK5iIOztzLfvaySuCM5m2cF8riXtsr6/E51hL3HWBAaEelo0Ca
a38rUa+bh+M1nBEEOeeGxyogCnjj3kFJDpBwx75lDs60/USIGvirmmylL9/f2DZzD/GWHVbZyLxU
f0khRW5SQ6lduKRbPCjqThvCL6hoGVn6FQ+TjI49H0oS+cYIXXKQHjN1y/AirJ5rpMMvMMzqoN9u
GbdSjgVe2ThNEqqzLBvkoXJSDLwOEnt/jm7oLE+jxuj8YUYi/oM0uO9Sd9G+WtaNm1OP89c4euz/
IogwhWHrqJv39ZM5khZ+l6LNtdaDq7ZnpjCuEivmuWaSZHpEqfzrsSuQcu8tBW+PN8+g8aEhKZkR
t7fTBSXrPhxWgdX1sVNRM720y3gWh+RA5qd8nCGCD/WVC1TrPTygcnL+lKePNoMnF6kc7HwA6Hje
Kr+OG+bEueGqPz4r15peiYmi13qWckar4T99fezpH5Jj4LApu9HtjthDLR/TuMfOGkdW72sPnWQY
srKUtsrVnYXYeDkwNQ6MdxZKalvEWLnRuNOGvS4/TIWDDjWTmbdo2t7rfHh5PQIf2T5r6bs8eBAY
hLmp/0EsDaFeTsSQ1IdYEFvCbQ8hySuaE1+IbJmSHHSn3C9xNCrOjqLmQIh/z1kgijHu9ZIjEcVV
MnFtGWXvNBp5xsjsPneQfpZyH/wD1gG4kGil1+04Sf8/yFdM6gWd7KOiT3RL9328l6Y2S/JhfM0p
yuT3C0ROfpZa1y14Y4jwH+jk1FKSnAzUkrre2wWt58WiO0C2NW5UykpEEtwwe6ilfp1DCHSL+dbo
VwA5VQLcneVkub/u5MiytCq4HBjUKJ2IRnvQa+BD6JUUo30CKYnQmG6j+OLvJvN8lya4bkxOSL5s
znHXquJLzNd13Qr7bKHE97zF+IsDQd9kDkXWPBTQT2lSHCdMS8A/9PUrGAxbe/jUW2rcVGAik9RI
mBNfGlD9BCc5YrzMV6PxWPyiBcpmFX3scTrio/b789pKFPnI3R89wL7i0FOIrH3Ee+AEQG9B5gII
7kuC8WEgl6iX13aR/weiZXMYqH5gg9/JN8qcX6/BlIf9ijg7acKO8ckfCWpeqC/L2jAt5DZbm0gU
sDiUysfI0jfC8n3AULoad2Vm7ygRuaWsY9J1cTwLw0FHfOgEYEXspyj9HoSjwkauVXd1kmI0S/vo
GP/P8RLYgxHSikYmnPQPxZ6kJ3BiMAi3cvBb916Lj54Nge5e9hX7lcLHxDrmA4nHdpGrP+Vtl597
UmVEbCCLS8nEA7CLOlrG7LnlO70G9W9sHHRupobRXxJ/TTyQ0oxV5FwzS8cPxqbMXLmLWX4md8fL
uG/NLywNNFJDaPId79UkywZY+4c4GHC03dwjrvVenCBOr+qis3BfbAuYt5ZVk/IRzKJQX9+/jzda
m4W8kYk9Yz3SmD0u6adeJJhZ3H8GRM8rBZL+zaTq7LuY9aRY679OUtWOPQjOpHC+4GvBB/hoCvBq
pDEZ6P+D7Q2reBm0J4SKOIHNqFIsHDcU/ZjI5dwCmCgClpd8D/O9pa1BhBej35U7Jbh1QRbypNv6
YUmvp/aBt4QX1DYmgvtKqPy0FB+J7nnWzl+k3GT4q2mUKPK6LNVJuom61eyo95tmItcATcm+1eTD
cwdDG2ey9m7jxzuEXm2MX75eGdST/PpEwxrjB+lU3j9Zm+Vj7PNrt4+uUhWVZ0sqtD6NwprH1rQC
YPxG8tkTY0TCA/KYxO8dK7oJAp3hMdkoD25L6x2zLoqrDuMpHLzwTDfBB4QHMfNXjTACNnmt6j1m
9KuNFyavMFTeWqiAuQ7Y2D/rp4KLwV0hRzvCRyOPxr4m7QYXTyatfIGHLMu3YnSzpa7/aUhltz1i
8U5QvJfAxSJJCxltKmHkdW5oeI3gCCurzCVlwZnjKSJFmPsFLdayCVFtIOkmgc/60MNg8c88ZpiH
3ygapBjRGiE0pSDPlNT8r3yqTPSEd9rKZP0shMVfLDB/zBE281+aO63M8MW5hPHZLQCEHwI0kqRo
vtCEUkPPtIvV5aA0RFKx9MsuWDdKNHvcrBPo5wdy6QX3ra1OKYxZujRjBQimVvOUQP+EQeFuYSPb
vlNIrF+aqsy+MLT3hm94/zHtWF+gHkyWyisP3CSOA7XP/snoFgvko43TtQ67mtHOLj5HgOF1N7Af
gG21Zu/rA3je+e5K0EtbH+tuPlaC8V2/vaPCzmqOdCAI84U3Ebbs2oKa0bSbpVNnbg8qd5VVtqmv
NAaJUJoODkGVX5LldKunAhL7/niPJ7vTI5GIkQYOXnmGW9RaN0yzDbim78Debd34I2ZbZ9muFcTp
Ygzsnh3lDpTwXPzF4nGaIYzvgkCjGabTeNTepbC4sWRrbwpfvk7aOEmVX7B3pow8dfjsKvkjKTjE
7iwHNqFXlBxRgZDq15x7iR0zF5djElRqq/0K9UTEnNmFBNeNKdM2HEisge4axhyTFqCMcOS91wnW
ab1OoSzTUONLnFHUwft49h2RI8c9zN488yM0ofRlsriD38sIyNrSbpDwVIl7guSZvqWuLllFJ5ty
pMHF8ITlHz2+hYuSQKZA2FHlf5uRLLVqWWFEM9w9lnmjjytFFW/44SdIrWGxro7ZodfuwkYTIxre
EHykvb08k+3tJutNaVYxp8SB3hopFS6F13YBiICmsshcwpTA41/b7ZidH0Ib8ZqrwK5nQGrmao2i
00BrLxOZ4tZephgwcZeh2soQ3ul4PQ/Eh0yjIZHadtEjqwErTcXmWLH7kqheF1grOqNWePDwdazr
MMLRAe+m7e1jEd4FmFkadOD7f1UKn/EqUWKAZTGcPQDkdhUk5DpdzAojq4At7E5IpVRIpG+w9qO0
Octbywd7YmY4RNmUViPg70zjxx9E4UW2s82IP/5C1CslJ6dRqiTGRQYOMp4L8mRvoxaUch9dh/1a
cxeGA6JjdQP04QGZt/iychA530OhV1HPfmbr0Aba4GPbZfxHBz0EidVGG/sVfuG9znF3mLg2PcBT
zQUTHHSlHYMMpULSiwBK9MKmg7t0l9CRZqOJn6geMEH3/3dL5/WiGB34OZjG5FIUlLGSjRKCuW39
RBkGbpmpqjB3hv/kjfyqhLRdSaW3+HtXBhfQg4S6DyOsXAO3nBrXZVLOwniddxsZfr4H1XiZ2Uro
jmk2GmPodx4wefRA+9eR7mJGDoB9mP8/YoBqMLrBqStj/cSS+UtzeYUi+FUNQOl0aGT/pfK49Dsy
HRE6SaOU6wAW3kfVNSKRhCfepI5AtYvO7gvnpAVHZXFCzYm4URVx6KkOLu1GFbeqWxGhravHoleM
2Ai4n3GPuUP8y9HesYJO1fVLZuibH+wd/TxBlgFfQVuZEC6TTE4GR8mZVqAml60CX30j6NB51Mbo
+JHaKQz3Jpi+FWEoiqSXMqE3/oXjHQeSBpq8dfQlTfqTEdlQeYbMKMTCoQi5lNrAt7LC6nO7T+h5
c4qK70u3jc6SZirb1aeX2X9LO/5NcfBzhHr/Ai64wCHBGtnSZ3qk1VmLnhZ26NRSJ5xfwS6VZaXT
xurFrhvs5/BXKf/0qI8hdsHIHDRYU2nJTo3C6uTA2P9dt7zjSUk7XvsaykZzwouVsXQX7+OqBISS
pNKDMtOGvVkfHS8vTjizQnr60ONi0HUNM2TUFtQju31oD1jt+9A4E9Sdndg+ypN3Thw09vOSHdcY
g1MkwPr490vO0INvkQn8d9NlADXhJY9kTFiZbfVPDz+Wab51SzVUkQ7prR90f6OItd3SDuAbLP/Z
4Ae2fmTf6AkoW8v3qpdaE+68m/1Il0E+KB7AYPRCxepWtVkoVBdwClEqg/+nj+RZaVBSn1dyV/sR
t9wj9ueuiBxpjdA+ZXbd8wiP87pl97CroYBCBRhGX9gEw0sfKydR/5V1Mt4dcOWKrURB6d9twC6m
t8cOiMtEBRfkd2/MIOOyJp3D5hxZoGMaAmc/SuA+eJ/JO1rtzX+wgLSr8DCLXpVyAlwE67md9Rjo
rj5AIAng43zkZfolmYeFh9UzTVGvhA2DO27ApEEQk5xMT3esjtIZB1HgxxRC+K1G6bCcGLnzZ2LA
DOSoWrhqXtL0VH4atNus+JS6k7kS3jznaeKhII/qu15oS4Npi7rab8o+ee1PlDkjtrjZz7Ii3y9/
pfhOwM+akQ4/hfXexkVlGcdXnuKX4RSdfkasJ4NdgwW6pAf0EB3+IrOJ5FyUez4resSREL7MU2qr
KY8fpiCIgSgUT/2n0DK05RMO+kALPVz4rvuW9R/MeSDznUEUVRlvABYKh3S/qkT8r4Z6L5z7+le1
NCg+v3oa8+zu2DHhIt0ZMSp02P/6VVXU7ux1l+KWMvuQqEkR9OSu4Sm+t5o8QAT/qZG99JbGR9KR
SFdfw6+D0QI4pBvJJ/Akciosifegx5O/kDJtQtAU9YqapslVLbqDEhDzAgMp8Fgwrx8xhfTXfIQf
Hy3aFD8e81XcigIL3zYD/xp2qLrCGIvDIostYMxRQ4KOVc4x+w/WYf43Dd8Fs41z2OzK7tfIgriE
rJ/izdnNofgIAzWJqoShVfqrqtp5eLuTyIQIEfd43r8azT+lL17Szcn7pLp9rh2st374Zuo30MlC
1iRUeJ5uUvMmJmsrXlBq13aVORtoxNKT6Nu2bwS2TZVChaNemTHfUyyqpMH0QNNxgpN3cVD+JAVC
4EZJ5+0M/NGFRd4GrySvbZPbL4Unb9b2xXXZZpgnHC2wqWZdaadrYAT9VUDGUJXTqwuiLGnmKWLr
H2CC1e7ZYzwXoqoxlaVAdznNzZgZDZdwSy+/m3U3n+TGCeOhgzmg8mFtCiPjrC7y+JAvi/Uicojx
BSUa4DV3IcdfXYPZl8MZe29bYy/4gHcMc+rqBVOzKGlZFuqhNU0xvRJaEyMA0Qbv145DFcpR1kJ4
YurHsgOemWJmeiqwjITar1hLTxgdWFWpn+2AFAOmWeUddU28LXu9UNQTlXRyQEHe4q4Hz1ka/Z6D
Qb3GOujOW1dGxx30yCrxXWhEtMxsf6s9vVPz2+Z8dXCRFplEW7j4/ndet4iL/mw9Dx6pFyAAJUGO
NmVHW5U4r9NZ8SmCQ+5E+31e1cX0x12HkJEdbvmjl+rOIWSJmK1yIEOmm7W17bhwWy5MtkNCjlxS
+/Xvf2V88vXZGyD83/tnubKhWolt07zsHihAsgtzi8NunpVi6z1MiX28h6RzCdEWgeCUxH4S6x30
V5fY88rJ0cs2fFWZoVqDjkT16ebwr7JkG2X6C82UaIZEgBt/8QJLcbfHqvbBfbGkyI6pi7U8iQss
7fJxU7xZGWfzaL2UtQsoVStld67VIJRPtHhH6sjHm3MbjvQH4Raf8xiV7WDoGAFGSrryANV//Xnt
qR9ud1y5/gE4YUsgushaj1gilZ5TslmyJaBE68X4baGhqkGH7CJOdwalPX0otXFF8SACNZOdmlh6
zSBy6UIUGCztuOUtWiPaQQ0Us6RJOXai+2ejImlNSrm66v2mmpmv/P4+6/XpGNa8wjOQAMaCG46M
oobzEsIYFZpvSxXbvq7N9bkbmVPzOgWjiuZL0tCfgPD4R+JAHw/QNGUFShGXxqOTqpANpQ1UNaSz
g5kz6l6x3R7tenUS3XmSRkvBtqYgabEdIuhQH5kQpF52GeEwV54/w+TDdTGc69uf0+aesu6rvSVA
tkqu9cFLC5ohTRRPi/t2tMncAywOtQwBgJtU2tEb7KgwT7udkNO+L3qkSNe5CINGGtgK3lE3sRjg
C+N9tTlF4jBZFgb84JDVIig5rrPksYMebL1MAUZFFpxMGIf/TzT/jaL0XmVZz2ctxo/I+T/X210C
KONH5tc46yUcbO3brGciB9e4lNeh9Eimaw8ZyhEeVbO/kmVmpeErzywifOfccK+Ce/UZJyICHzec
bnOVn91sMnu9uJD81V0jUWWx7+qSOcQGlG/Z9GecOwR/GNbcd6bAGVj9vCFmlOhOlikVd2AMcpNQ
cmucFI32dJT0+Fy0VECUYNhWFoKM+Ru5adYAdtKocUNfj1OMoWhLVv4v7rnq/W6elRPG+XehO5b8
gbqg+ukQ6/UNKVGrRkxUbrVX2dlfnIYgKNAV/H2+iUPuJO1VaRu/n/4v+mfZsuQtWp7pByVvbUKa
uRSN8ymG/PdPtW1rywJahjrHBtcqEPe/PWysZPQxPleF9cYpOunnGzn56hibOKaqcR7sq1H47KKw
0aTlitUblPBE4GvNK2xgRtqGYb48UjxkSvxnZpfOb2lPh7sJ8BsVk1SL9UYHTZzkJ2DmwFJSLkUh
77kRtf1xAWto2U8n5QPzOHSuED1Td6fXMEqhm37zu9NxToOpRYkgRMlcE++lBPlCY9c0f99E3fnB
WXZVcNZg3vcsQiNoigJT86vjomsDGmQvMIL5iaK0GysbxbpOLGC3uDorlPTfu+C+ixg6dLNQVqFk
4gNEqQ942y6VY9JaQUrINd/rf/r+sVKo+7gm7I4c0P/qjEbCLJxzvuExnK8rF3hTseKwfqiyjxDR
BcUla4qSMGR22VcBKI80fGbeNsQ68WR1G74tWVxs2w6RCC6BEdixPjpTLFoWC2Lf0n1HS1yOOWdo
QcSeBLoTOmIfk7Hnqc90xsTV7EQqP4lcUofi+nELn3FJ9J+juDWOlCrlfldjSgDoVx40/8sUe2JD
5eXFPxGhO5UJdpgkj91D35wkT6DgjX6/xfw9QEBaaYLJdL4fIf9zXIuITtSlAYhOZzX6rICMvxpe
v+ZSxfaiaA/zNJgkKx9NDyTwOnzN2dlQjjacmH100xdRNEJYXgHvstUKAWcaIYtKpAhPypmBaX12
xTVekxD+008zBcgozc2CCYdpcn/6jay0nvszu9qoHMhuNwQwrOM3lsqGoptX2pUj+aofjZJUbINX
0j1kWQ2fu9LyP8v6kYDhPylFGz6/Lw62C2KcevpEOKa+QkEKtvnDSd5z9SWly5ahVxxgd1PQGbfP
3vpT4b2Jb3B6WFRmjsE+89fWvqKCysTTBLO6vuG4C28G9bALlb2FwSVcVPwoJsPCBHvKSCmKeNl4
N9t7blWjTDSH7htB5BgxTDLREueUzyJYnEuh02hbdvIiFtMu5JI2dAAbxznbndqvCCwz62llZELB
7q0hejO62zkbvF+oHThMWe624tZfHlrsuayXKxlxj86Ury+KC6d25KiaWU+ZKQH56I8zEwqRZTug
Kh7Bev6uXIEG3veKWLcx03cEge8bPk0Q3shG2hZVo1fEevxMQX4/QKZarXF4FrhZIZMHsetNLeny
csBygmKK8B/Kovxq+ZJHdXJxerddqsrXac67Yl+7U/zwnplI1/z2csIIbHdkeJousHyM2gUU9C3a
WYLMpy1UJ40DKtslWVksAsCDUunl9E9+wHjr1z60eBoyxvrY7aqLY6EY26MGkH7FbIEANNJJPB+q
cmRNZQU8UCKCnPSuOL8kKS1vQuuCbBSbh0oBakUPJoFz00+O9Y/mhr100wvplB5OKB4OVkogsrOW
anQMiNSJFy0NnAS4QYP1Qr+OzR4P+ReyLEYMihgIInMMHJ/ro+K63OZPyMSZqkH3onD1A4pfV32X
lDpe9xdbtNOdTsdb7RDRu8dZ0+Km/TnxHc2lBZureZY3cKp7gGwlPZycocaPTTgOSe2QuMiXHIiB
5EWT35iBavTazQqw66sek5l77pc75Qfp9x4XvfeyUeq+WLg8FZbPAR4hTTS10ZYTjznFKgJelrej
k5Xi5cP2OwuZ1iVWhFj23gJLyhRbwI7vKDKekFnjZ9AsBuWaGWCR7KEbx+d/slI2wH/bf8ky5pdb
uTBmpNT33O2TBavF+py4p/Q08+n2LTNE95SxJNZ0IJqXKKKbjn7GyTsjPqByBW7P1XkBUsOlMMaw
30Wrik1zvLjuspLrRBKFF413/s+uOvma01CIN5E4VRl6zHllnHZMFkWeqm9WsobuHhBzRvSrvEMZ
2an+380MTlmaqs+af6ztLJceXWEysjEWQ+RlnHOVr/AY7tY+WOkli9AL1azmFeuByv82vG8AA2sF
lANdxickgA549ubBmgcBVuXBshUH4PGKvjFB29jU5mVujTTgqsEWAMCWDxg0el38K+j5RyZY4jKI
DiV6bQR3G7XSDz9wF54G47S/NZyvRxaQQa5krmwhoctP/jnBAf/y1ZpdmIqCWqFb6XQy9j3Zvohj
ef+zh+dDvcrROoKJslzd7E6R2ZZ6WgGwUKm/eSCLUaVnL7cjod7cAOzBPSfvl/fOaEGZkEs8PdZ0
mXKeBp1igWX2z8wiBL8OV/ysSwPqRiWRIQgdEQPaipE/9az5bND6aOKfdLy4ZtGdg/vXpGy9xl9R
S4PJ1t5aCsNsv71LAJISWgMwI15P/oOMXsjJTD/12QcvAVL1yxcRI3Gftglh+N/IyGOvvmW67Qa7
lJDuYzPjElQ5KPQnsR7DT+fxBlCOnlmHtV80RgMe2tKE7cfX4v6wVqUUrUeKtD/2QkJ4A3TVIYbr
RZZJlwYzvQlV5W8LGnNOLwyW6L7FM+/AmbxRykbNKSdVxz77RTxBqZNV0WCYbz2VRMU988310Bn3
5NcYgCIZ1EwEUDTv77pNF6Z4gRC++L+0c+KweNQwX0H32WXdO1CG2bLZq8zSQSWcIn4Z3kc6hoYj
8baDbr9OUZo9ViH8/ocimo/gVD0v4riThDBYUAynUfWUHOtEzVIBUrTiUy3iQMYBt9CFWckouxqg
XQhqQcgiwQH+vKaV0bS/QDRP/+xZC+NTwv5xvRRkCZ3fH5ucjU8VVegFUCDZqogBVpGSuYpqweWv
3q3vCZZS0nggM2cligX9h4B1Rhm5d1xVNyOJmaWbbtk3i/NLNQMP3yF8YLQng5srq1BicfTHlFKp
7O/ymoy/p+DrHx+GpEce4iDuVMyFyKkUH6+iXFE9DJFgGuBW2jtFC4xU0hvfNS7emieRAt9aAJX9
XA2oRurW1QA16bTinjB4ZNzOw33eeYnrSRw4OSJ439kU6IjroDjkMkrAi5eYh4wBifHr7D7DwQKp
F/fHbvMIJkgZ2ErV3GcyUTwydusMFQdoQ0tBrV9tXryCi/24z9YtjeBSNnZFXdpsAbgJt2YLISDM
tn9rMG8Trr0QHA4ZajbQAhqIKn6e8NWATPgOKSO3ZhotceNWPPzYf5D5YUWdlO1sfKbgKIeN01E2
uAeRjZ/eihOZEc4qemnFLqd33i7ETah8YJUym28Nzg3lBqLkWgINMYXXnWzMoBPforqtONN3cwLK
K8LEogE/TmFdLD9T19IjE2TW15Can2dnKwV6vp3IgIkCwQzohG30ReTuSz4QSg8aPtCc4wbreTrb
WgAVNGCxQiVHDwP7Z5M+uDwIyUjpyhk48sS59gJ0pe+7F57A/WRi4AneB5CuWzl2E+wk6+xBX7zw
gSVvyWfhIRCYg7LeFLJCVEN/zwrfKPceKzQZ09MsBwJlq+yhJgRaXuHAWReiGVMveU3h9fhcCvFP
8zMy2WnTLZfKSJmXCz0o9r2Mcgh4CDKKsoOeX1hmr9uClfDP4pAYGgv2cCv7xUa1PzW8xIjzwtJI
9RuIBQ57U89ZZ2aWxy/yBWr7AYzANWaT8RYChq3Dm/TGBWdRFiYMlNQTU6s8AOyl88AJleCC0U5j
fM6iX3ufASSUgO55yLWtzSErU2Ft1JdLQYwLI/u69NUCPZBUTjJInJam0rQvhezzdGhFirK0tEMV
hQGUUHc3k2uEKI9ncuq5HjuUywV6WmL4Ztgaw7IT0ZJfty4Rd5YEshIxqso18cMtvh2ODUZVuO34
RP3DAgYc32jO3kZA29dIn3z4q2rpkaMvBQvzjAXP2tocM54EHWj5LQJf2N4OwkTRn5Q6GRjCfqTo
rEE/LOCgjsgxH7upcy+lmOSYxR785orcvP9b+RLY5epNiY3kRoow0/vzRnBxs6OjZ2RIJ8qchwKS
UNEEuYdw8qQ9b8bas/8EiB/Wt1AT6DEtoCO8MB/m5hFvKeJjTXrY4SD4ODjQ2vVpHhtV+nM5WSr0
Huicj/egn5eIDB9lnWp817r9gHBwe7DF5sJ/N0w3s7CIEPtn8itgIOm+PczsCQE1U0gjA6eBmmBx
Ql5EzAThdns8bR+X5Wg2U2ndRqjzmjv7TJVkew9IM7j0O+e2PdDbfVp0H9DShmJP6NVUG3K0MrSd
J22pRfcTetRQ0FKM48tGDjkxfTixvtCe/WoK5IjbJTaLcXVIdwo1dZwDcTVEgRDFbYZVJCljGhCM
UtsJQTL364zbJO1Mr/7llV2D2xrIgyHXtpz0FI8LjtlAAQ6g4mmqS3g2/DnHMfaRGvT48szcujXm
bis4PYl776W4nE7NmZQkGUHi6wikx2drxso2bMe+H4v8tmEhyxXE8jHqadno/GGmNZ7D2Gloyc5x
zuQYPWLcmb5Efu1q9B5J3IA2VhN9WjsMmO1Cy2YbMnnH43S9SicGUv5VncgDw8R1uEcyb/jiWDL4
eIb2W+ybX8KKyebM6P2fX7x1kgTza9BCfwoVM/3j7LR34N/h8G1e6KUcDlv1KIr8ueOQ0ZsRcWPd
YkBxJyLXD4J5j6iKWDpU+A/lIMy899/+b9SUdwGDH17gl4L2pe+EMB48Spdh2pqTz0j4NIFnIrKV
IrilzuycwdIN7OunOz8/dTPNrOjuPwSIVkiphYSklAoXPINFbGr+mHYloPTT8/cV4FyyYvsod9He
Qa4lFl2GEl+4ABpgpidN6mny432uhjdBa9siWA8AVEB6U6Caha1Sl+UUFwDL9AUhU6UI/dqu8FZY
q9XHetlSMVHqwj8x5kzL3CopLz/CAAl404S11n7y7DIxfNaWny+5ZhV3IdsF6qe9J8KyBvNOONB+
RchAnQgvNOO2d2FZNVq5hCyPldOeCZf9Y8Jzea9oKsSmdtNPTADBSfegN2QL/+PYdr+68H72w6Pv
YBIQsGz9plOXwBLoCGwKsHy4Y0T6HvQXi0ysKj3+B8fZXvhYWIBrk1NlMWe84CJTgDxTiVsAuocw
sagdmQ8GN4GX1pKA/MLozz5F1hCxo7uHn0RSHv25B5UKWs+RCm3Zb+v+G6XdagrhyjvVAy6sWng5
aVhht668FaeYXFA2Jcg7+ZK1eh//ib/6nUt6SGnyOdWEREJSK0Ui4i2zhIs2BaCfERUmDh4UBSOU
yFHcwoHC6CzSdRRoKlWAw4YfyuJbETraJ9ua+fuwUGpo1Zl31rEXbJJNKkdliQBIpq0Ywwo8Pjs1
rbnxwCMxhXPlJVEl/8Lz5ds+Z4XvTGM94G6epnadsuEwA5o41F9LvVqFASHWvoSeBXB4scVV+Jtk
LIgqAuTFuucB8BplWl5M38Q/pdPTlwHimaZ4HFbeatki0s3LP2MYnRdAJ8Ox6TpbKNtGEx105q53
m18+FOFn+PMt+WMh/TdebwQ3xShhZs/ntPMLasmwGPLEe9FhNQRp1GDdDoiWF97k9AAUHMBrxRP9
3dM5lB3LAOYLU8I+BXMKfE394BpazVptyA5SNbkEDXGtXcAMURGN4xfn7G+dGeXAjBVaaAErZapV
qS5Flwz/OhsuJKTjuXlvmUtFzF1Us4YSHmdxtBBth2AJketg0ACTU/vUjpUUV62XIKTNG+l6hcBU
ma+Byq0o3peGz7Ks7FtHWlGpUaAL1DMQEr+yef9Fs92U167eTySanV9EJkZKoVvnRTj/qGq7KXuL
yG4gExZVRYZOJDOrWKDGMgxw5IsTCisdg02xaVZXXuvQ5UZDXJJ+fuj+GWIUNg2JnOTJJLQtH/IL
/doFbcDqxQAwj1Qlen3IX49WJu900wC+Z0D22TYeLLtSYhdIGABBq70rlER8u4zKCJIqZbNEMIaS
rcblczGnDZAvdnF6gsMmnvNg/v3mNW8Dii2sAJhqumF98ikWX95fAIdiw58+qsmxped4KW7zSYEL
l7ycMzyhFxS/CkZrkLjpGE6gukzGmudt7zXrBdGuaW3h5nCf+BLLLK1XavMd8uxq+2Vi+c784Z76
guEIhitoiK3wbIvgdEj9RT5CNIQHWGGwcijQppLfmHk/mb/iigONWK/3rgw/j5uNcZwPjbKP3j/Y
y38t2O9CSmGBbN3SLPMtYSdRwCRxhhMImiHK8ADhE8fl4IuUb8Bq7/PZCUbCGnXt7k1yRJTFYSFR
O03iL2DsAx2QCOx0cVh5brTosSLaIHlgK96EhptEdqYP8Ug8RAxM2Wzr4kbnG7cgGibU2qh86rnt
qJz8dPbg7FwT5293UhVBu5SPEyXv1o4JYyk0LY95z6RwRedXYEjD87cVKXZg6lwGqt2aaXsAhFGB
7rWZ/J2+0KBTmqIfk5Ro4DdTmZuRf6vxwRExf1KuatLP72i5w7Hj0bogfWcdI8msZAklC4UfLq3b
Jnhv8oMM2BN+ZM5Izv4pwdR75cnCCTKoA2RXqvW8q9f/TAw4nfQ1fJfDoh8x75TaCnNT3ZmVxOm+
NWijadDeiH4xpDSaRQu2PWXyJspNuOhSR+bg5Ra7BYmgWalIHR3ZPoZxCycCZusUmp1wk0C9E/yU
mBMdGUu56NkIX2qCNw+02hqq+mDQymMh4Pz+WyL4FFj9qMEj7fT/w0g4YPcAbc0gO8Nwnt5wUS3D
CHKP5pIQWc9h4Ho0unFBiFIG7yzbQttjb75lNFFV3uTNLK9cAQ7GkWp9OGANDpcZpoZ3qVrNqZkr
nh8v4pOWS7FTIcOnM51PgL86rmtdMpSmHMD4Cm7TuOH5GFl57huaJSYUTC7EBMr9OCFIHA56HBKg
N1KpjbnJ4MedOeaudEcbajpJQph2/e4VaAsscxyQpX/SPL3Y/25yiwdYIAQhJqXNPtIRTj/tCKul
+UQWcPpHGRsU4d7PKzBu0Jx1J6DgLh3GnChFYeEdyufXSUlcaXvRGZQ1oEQYN/SF7/aw7nA34dZo
h1M2mHoISyDl2u5lwrep2WZq8YORFUZ/MfUoETG2ojSp0eAhc9LgRB+vzZUozXLE0x2UN7qxIjtx
n3UL9y55J/IK8tgY1fnQW3uxWZZ07r4YfGmWiuDo2Djm5f3WNfVsDYgHEzSfYNAx5k9kghna5MA4
H8ZteFEUGl9neZXMXz+SxQZXWuumso09vvg0wAJQhILc0xd5v9J2LCmMKSK1m2MaNh/CrI9tnERb
UCenmMmuR9L4xSilQoo70og8RYrIVJZjYRnfE2xfPKQA9a3kBqHo3bKuRbsRVUzYVgZ6dwlw+FN5
BxgcRkt/iCUL0xv9VxUBT5BmL7cTZR7m66IQQPBAjOwdCPLBvpdnc3EG3ivfO5wyeyTc7C551xq0
hUtVUrD7toCzRme9YvVvs5JF1WbL7Z0gnHa6LdPJmBjslQMuYwIbvbSgegTBgkXXRYj+XUnFhn8p
CRD7JbYofpKJbnt5nDqOmdPycuT7go4O48efo+J2dWiEqDay1e2A2t8mEpjJnqpShjVxCL1Ms1/b
UQo9aLlR1iFeYlvVhEaTZctR0qM7/WhI9UxV1QBsw6yeCFz55KsAepjQ2gBKRkOHedEW0HSxkEmv
0dbStakBMC6Q+g342pRipCn+5Ua4LiCWjUuEMN1qfs878AjqhmJnZbgCzwh9KMogKbgQqbjT94rw
n7I1gZdLXQXma0d2xzIbikoVSly0udd/gz9lGgK/wwL3wH5/LXoze9tsoXSVhJxn0//MwTMEE2Q7
6nuEIU1FJ5sA9ax6Z5uKBxlhWZCtOWdUHSZlL2K+ZxekpWbn0AijuNKFY7yWxjbq83y5QwDC3Z8N
nHIYVJPc2+/0Cdm9yeDKmRMkNrvUEj0h+OrqfskZgN0NbrdwvV7efqXvi3j+GLSAR1FBS9G/EZxM
8EgQoMzAz/D7FN37Muvuli7GYHRxSsqYwK46h6n5Z7bsvInAj5ESmLBCxNGxqhiZAAMdYlOmYc+Z
dO47s5hKzviDRS8VNWYQB8Ddmlox2Ps+b4P9zSoezTyNKJWjlBxwSYI109Z8zzvf1LX67fNm5QCo
XiMyUkJjA596M58mIJOnZUXAEBLlLWXDvTjLEGm/OVNigX1PH2YsMqyE3tLVkuXqzkNkyIMF1jb+
PULo2NEB7d3zFHW0tZaT6oABUzlNifXMFATtMJUr/xVuh/HENNVU6sBShOeSKqzVuOZjDsvR6h4z
g2RSUEwg9JnX+PTL0eUyC0g/oZX4QrvDBktXnP94uYiiLMzQSrUyMVszsc3hKQg4bHIzI2F0Uqs+
wjw0HxqJZW7XepqEOXKeuTyxuPnJagD2/ENdohIx6LQmgKh2EUp6J4e/a7pABI4yiG2j/2kF6B+m
gb8jKu1JIn7AOYYSFwR1WmSaMWDupz7Zvbxop2Ma6BGqxOhXACFjt+izwoV2b8kUWepGCmpr/l0V
kpgqBef12uyUjOdCWTDlRDIzqmgDNbOjZW+9caM/zyGA61cF75CwOiGQ2b8f6PtpytUpamafKqJf
CoO8W1zLH1AbZZGvWJ0RqXqDep00TME1uMPnEwP8Nv2JNNCbTQW69dQ7VtUO42ssXc0/eEfwg2C6
c3QInHxb+KofUpuCG8ecooBCAFPxGHk6n2eglL2IjbnPrnixvlSvw4JeuDppAyeKZkY6WQxZqGJf
54kl65YhlobUkYyjndKGhMFH2WXVo0M5vJk0fJDjQWcGXS7rNEIGruj+DDyelItZvu0mCqNRaT0o
JuI8/6/4ducOgqKEvWuk2REPR5LJLjAFEsgxGl5mIh4lGVCFtceJRhlVy2ZIHaxk6OxgXGZZoMzp
CJWEKZf94cH0ocU++kiSZATN7MVuiKGWzWTdtsYe10aGy7vEeQTyRSIhEjozglVsyEqyTIy3Iag0
p79gYodOJrez2JeprdNddmdjjg2WCtY5XlTxkqj6zhGtx6+m4i3x+ND5wljoZDqvhwGJ20W0PjVG
jepyu8fY/z53LJmRBGfPwvmCquzvmrSTLamV61s+r0w5sFzviYkAaTBfAlbZyrjYJORp2mbw2Sl7
MuWSOoneoj9y4FlnCEuIuoAREuOa960LdObirIB8ZhEaG3H2CDxT307h8A3z3UUJZ39EtFxI1UWe
eQWBXrJGLQTEh7G+yvixze7l0Gb135IMjZHAtAs6qSggz9ydh1ht62CU5fFRHeztzvFWwHQKwAlB
67SIUZPzZj4ln0i7G69AOpIH6fCBvcRo3r5azxzX/NaZVIdthFDiSl3N8u25QLGpu5klF7Ys7q4m
ce6iXblwVKQTV+96QLFhMlfjJi95DEPB+s3wauG60yJUMldlh5nBgPz+6XUuq0bwZh8fqxhTxz6T
P9Yx9Lq1mU3dMYNVDh6WyC2qrFArXPqylnHEOUc0SlDbdJq+XeTJtAm5jCvTwMktp2DsYBFdUiDj
EfhQxjz77IDXoTaVWa/90pard8Nq1uOA3Iajr00E6PXVEaMTQEJSupe7A1KpnngKI+o3yLFeJp3K
bffsx4zW1yu0VYjGfrBC7LT8UpoV/fVJ+OxX1ABPxYtf6ZNLsWZxqKHd5QNkwT+aGXpmlnRBTwRK
0RW10+TgiENWB5GPQ2QkxFnSl6pW7wHxahl860twRRsl+H24QMPTaiXSIE+BugliigvJnNGXCu+N
1WSpiZRUeDPDU5An0qSVLAYmh6KJBLLH6KgioATl2392iiGJuKv2Hx6+GagBN34gAhCOdZebCMMz
h18W1eD8VZINcS+0tuDJ3KRE/txLA1YI/7TqyEHbzmhwj8wQGN1e8jbg99+FcXtcsl9h3ICPoXKr
Al0inP4nEoSv5Y8t5AHpkZGRHbXzSqgrQW/KvC6FKO89t2TjpESBAjs8J3GWQiK9NNXprmBL47K/
LLfzK3J1WSNTUXO5uFcvNB2/YU9oKcX5POAmvWD/e96DOz41Q/t4bhQzwA2qt0sgvTj1iGRmApsj
me7RiCHRqph9K+QiMkR796QckAFEUavAIp1S2Gi+q9gCIk7EwyShMXRx58BmntOvGTKJbl0H99eT
vVqgLYG6hji+9dDxNTOEgPjVzU+L+bzAyWVvYkgUdRW9S5+cvIcAuthYZHNBTMEEcDB6gxr59G3L
eedivTHxK4l6rtY8Z5W/JP+E15UbopmSolEpQIrqaVj330Wf6Bof7hnLxkx+2a5qItJExLl7hqFa
tkLw2ANw+e468YBlkSGNs+6ZxtKjbZGh2TFA45Ry6jTR1OEUVudXahmN3C0WVLgaNVpW1Aq3hhJG
oDUK+07HjVVAAYPRrirToVJGSNrbJEM7LqexXnuE0VO6Z8wuAUJ5HhtM9LOqpXtg0LnhfuztV/kX
QwtHtlxL3zVy9yF1CU3IJ1ygz+O1YEePrKjNIWycoIv35Yy2EHG7PmAW57wF+FXIYHdKR9EQrcr9
Jr5bcxTzwLAxxTmvrRnDHqKPu4oAZs1IDtrg2HeV8RsBydpBaaxfH1zPiDEiN5lhg7sZ/QIQWrPT
yXfhT0UmltbfCf0n4lY5Z4Mnrrpm8iz0J2b+yFk8jnrRwmg4UO3jsFP+PCib5xBYkYbgndMkm83F
XBHHHH+tDCtUF/w2RYSBoT4zV29nukRCaxjohsawqp5p/bzI9jQ7ZkKqScc1ww84E4atScP+SMoB
9WBgDKdrPN57HvU6VIc7Gdl8ojjH22klUR1v4LLfJKsEh8KVvqwfhXr2Ldg31I0xr4m4oR8qqL+t
L9siOGKmzZUadb/rrvDeaM8WXQYzftVER3GRJrmrqC3yKPZg467DlmBykNjKLelgzVwWhR2IvDBJ
rEUOt9sx/3dVm91WaojEAjvpUwkCvkebH2TYq/ZN1SYpEDyh3e6Ig9Iw6EKoWyIcxf4tHR9SVys/
GSB9+s8GUGE96s1pYQ5PxPqdN0dvgrxOqK5u+9fKPvLuofkFy0CK5khNRoKvcD/8pLSjn7wVaNiI
+MtImDf/ImJznr8h5vIbR03IXoXkOprG710P2pxUB5pHNGXuVUvG8TGhKSJuaThn5zHWuJDK7eiI
jtuB42p0uNxiITwX9PJVGmn14h7VMyFIL2kQ+diwS/u6cBaWTzEOqcq478Dndol5QpAbM52YU44U
ALU9NEx6QV1oki3H81pGDp32VHf8cR08MDshCIz83dFhmo19hnH+oJu9xpXi2zA7aufExntHALZ5
wMDblyXftfoWE07QCPK5Yn3sINjhNsyqvXDCuxosHHbzKRu3aqRBTJtj2x66G1NKi+qx7yLUAMxo
hVtBDvryBsIRQIchJp+sU5AwWPcgGthG1ZP5yJZ0sPxFbewmzqsZUPWpX2C/maau8qP8jIqO0yAl
IBhBovKmUiYrnxwYRcXHJmNZzgkyNDs0D1WFI6DubMdEtedUoaKMSEDBxkH5re/+A9FZ7QJdyOZR
pPjGYYBlF9sfQVY2/r5Cc12wF9pR3bQhkltDzKBblu6x3jyYvFhGqnChaqFxChGYUlSn06GxroLG
nd99iBbISB0zw0xk9983ZpNt+AUMpb+7qFNhTocRo36o8T/TuXhHLosefMMGR/AXiv2W12sU03BA
YiX06dq+r5HEKDd00rh7Z2ozG1yjfXBZMKRT1UwO7CQ+zagFY56n67/1WOm0iiBF1PIa/RNuiQ0T
dkD9geBp+XtIeLNR45VTs2MmW40TP3Ahtb9ioErV+GxdNqTwyznP+bxlB5y88ouebody7802MvTg
tNgrjBJtaoPazaq+6XKvv0cxZv9q6Piolvw5MV9whpQsmvxRspVwN+Z8K5QAdtb5xusgg4KA/bVV
JRlpjfEroYXrtgwao52UG/UJbGIHGhfevZk0dZ5jvsKuGsjzbNiDYS5KtX5PI5e1KNpMYwiZv/FE
zle1cZ2aOUyIi6eiicP+1Gf+3i0Mvb2HkzX1te+J/O0BWCngMKiJ88HWsiPnobgpLnjquAJEIpDC
Yys/VQPKAM2EfMTStY9RA3krt9wk+N7SczzTJqr1tCecchAu+uDFd9djv1IixWOVifxxgKSF9KT7
4/qAJK04HQYxE2sMETasEwgUWmY1jkWiZ1GJ66Zt2o+x/O6NzudGuAMRpW3SH3HZexWTheEqcMqZ
5ZGCfIuQSJdtg0ljPPgBpd8KdD/HvG0GT4S0+DRtmNrcGWeoOfZ5wuzw43E+JfaCqE1jZEy82k+5
9dpJ/2ISD+m51LQ5EJ2lrpui3Cj6sjwZlhNbMp8kcG6aMnkPY2yOd5Hy9Wjd7iIZQD7o8l2m/QHh
N/KeS44fKJGLdDB0hlb8QnBk1c6Bmm/oxir++Udx3tu1lJnzbzPPIR1Uyvkr2PKbl1ru1jMZZVOK
+CTA6WIRSHyIkTK1H1K3puw4DjyvozQiE0qkA4O8qQeGZi5x105eF0kWR4WOcPfK3QugVCwMpoTk
gMM2mn7lhlflYYOS1ROd0Vvkcc57I3WQ0nC0YpgeQPcB6c334HDpHIBo+I5xmb3pPTszluwq2X4P
sbiX7WO4LvdB6NkCadPCEcu4sOg6bVfBL6J+tqIyREZXZ+Jm6NDqxxhiT5a76I3XbAFBrAFroY7q
eV0fYEiv62hFLPVUyCViuB5W1lfUrFnG7ZmH88gG3tv1hLnC7m+EsgnS7uFYNo/h58r1x6CePqTZ
xSHIPj25koFuVvJixc/CuomlnoC4y8TdnIz0s2mxZjqno9NCQ09WIjLRCj97ZcJypdpNhsFEPlm7
4gh+KGhDUnsNZG1SkNGbKp5IosB+pb4tacwAf5VZpCfooPgbDKWR+ms5VUpK73yc6UXWD8koxSun
Dai5kHBmTLaHPYBJbKEHAeHCXw2glJ/RmdQBs8eUfCvrxWj9cPe/eVU1WYDdCaVnCVf7sjRF5zsZ
p0vkbgxaKGCLaiUOFsffJMicafVFM5qZGRVSk4SenZ7rMy4GeOH/lvemfKGxmEtSFNUuafkDNiB9
OAJmqjjRowVLqtvCxUBAHr+MhSm7Q0WmafOvc2NHCnyyJszRat4mQ69vCe/cwKdXuYXgYvUhEcAg
0I6kMgXTkimqYn8Q+Hps991rYI/Mxd7cmA2tojnmYVDI8hQZcRfPEBv4da/6NiL1Y1vTbgK+MH6J
7fcR4a8Qlwzw9E0jXheH/IMyTnSoYgDaq0ytIiMSKAJMZyW/UfrbbU+k7x7dAisBjUm7IPcOZ2sU
9DGVUCp598b1Z0mPJ+vkvMnU6IvjqUiia9ebZF4rvzB+vSSp8iPSM5rCD52lHfAhI9OrUdH1v+Ax
8fRNrlDhAyGfPNYwfBk/gsxntJnQ36v45AqO2fWK4LF/JkIgodSZiEDbZnNTEs8s6eYSLeFsMQHW
ydNvo9AgxXM07zTDS5YAUuq8EfwYjArpJQJGot6NsaBSqaBO69DsppCTGepehSAqKI8Vly1xV0Fn
FcZeCTODhL59EQg4jiWhrneC9zCsNvlvyovJ5N9HdvCLluHUUVV90ICFOwVWlEKnO7oxaV+EujiI
AlknEhFwu12G72f3rSAzo11K2yILbStxfk04UlIecEgLbszibvaSUg1JtGP9xeHpvK06gKMJntDe
cCerkEwvJ+G7nkkMp/fjlyFnir6jTOat9WYX6Dw6PNKPsDkFmiPQqtXsHQDUd1C/A7a63yTuwlpz
yEXsiF9XwID/YS+M02mWCH/jNu2QHAyFg3wqzYbVwdnJZ5evCWl1nEFd+vkQdBCfw0BW+7orqwwp
6s8Ntks+nrrY3amh/xDE/nzW+a9otOVr895L1fCnTqAr9lizGrhZa81iuEy5evKokqC6ccnUWowa
ruXgPIEjsltorks8Lw7F7eMIPyvlFWN41Sq8YegBbbeWIKqPG9bqyPwfjqIfKrZEajbgeK3vKSRg
5RgtlJCgWDTQ/lWUPnojErAmpqy2DN+95Qgkfzt2Ob2FwqYyiq40+qj5c754jLxoMRsqllLIx+ri
4CyHdVYKLYK7r8SYH7ka/j3g2fpU7Wt62OvERsr8/rvYH5HTwlwBwBFf11teURXcoXkggw33rtOf
hR2uFzHgeDRzFMBGZrBm/Oj2I+MDYfn2KqCBq62/TZg6elDz+DaJ6smGzpG1n/dpAOWtGx9XsesJ
PpQhysaXuzr/x7TaJ3FpEHLsc8xOEIzPnhmHTcKm0omV7LX7PgJI8xdswOfRcPIwuBNI7HDfcutL
VaC3Y0vqC6880o3GOOVexB3A9ZUooJpRqvCZ2LKaqLmKXFXnfzSIc8aRUPgRXCAW6aj/MvllHWa7
GHoVjEXL8Atx/2TOdnSQpfiuKBcA1K+K/UFH29qD1oCKXw/xuwkJWQnYtXXM6w2GZuOYl5wLoEio
UQDXwI/bnh9USylTzDrsnV27Uv2GnXYp8YAjj5ma3jR3yRt2J22kUEgizrapgwjI5o/5EA0yOBGJ
3u8FAX+1tBGTScs46eadJ5ksYORaCXaDvSqTtTmfmWiL7GlkU804+o+S1L1a1TGwX0LA2GfH4AYd
mFFKi90qN9JspDb4INT9F96dp96LzYFPXYbpAB7I50s0Qir4hkSxClysdiUvuEIvRmcBPZObHRjR
zDnyz+fE5G/rGw42E/RQmAaRg8F2k4ihwuAj2Uez0haojibcK0d0d0EzDGDexnNbAFhG8LUY/5CF
fisjpTvk4B+SVaC6r9pASC3dPqG5gmlryRTbt5Tkq6lNocUYqA3w8tbvz/FMOnj0gOUmy1VTfI92
Et+lc5aEomSZqNPhE3EeSBUNBuUIS6AmHqRSj4TRB8RpxcGNIx0SQ5HdXXNgbniGG9kqpFg0JjQ8
43Ck9o35QBTMaHJtTcG0l9Jod74408iwYRP98CN1lXlxGynhCoeERtd4xkSmkl/W9VUun0fpnfiD
Beep85JAqD8PsLAKZxfvTXhzmA2Ach1GXEBFMDQWMJb7MhwLwHeYKWY2mPWW7GwE0/oKl781G+E3
gAbotyvwPFgNng+GbwA1KE2JuB2y366+xbnx6ftbLVOpFrDyhxeS5zaSxvXcwi9Ao9hu1T2kn+6G
KPVxvgeItwvNAjq/9ocFc/CrSMy5k88P2YPj8Vtt9SIHFCso+/gcaEgLWbzaNH065/pr0wc92nbU
KBRH6RF1vdJ23DolS3yVcx/EPFkU+C/xTvmnan1KUYN63yUIrDp+/pnjSUSCvco3qVKMrr6hLBPP
aN0J4XM8y0UB2fKJh9lD/2ZaxvSJiQYa0vExHEMtMM3w4eVAjOR8mYGQD46U3wmQGYqj96V7HO5K
FZwYxPrLQnAFtgZu/xW8T/hry8dU9hIYv/VPWOUa0o4y2bZ9nzrPTkB+oLBUHL1wWzi96l2k0IQG
bwN7WR7IlfHhHEu1lTmnsSP2KhRWwT/h0XkK0LUgPlGulsmZPMWz002RmjsTNPiOweVN2ZXTb3A3
jXkaTTM9jlZXa5i4/mQ8xNo9w8FOdzOVdcp/0zXvn2/c3EorOP+lTEFTIZ9NIm1A/CBTSdW/Lk6E
G0BmyWpPDORLaeSShB5qqfPAzxvPph1iqifJ0Z2xCAqIfbiahGC79L/Rawgy31m1hTdVjeqJSh0A
3gjEZhW0z1XbhCNoeOMvmprmHlaRByvjXOVT7RHMg3Gnw2VboobLhAKJJT8ozm1cBlng3J0kcRoE
ESv9HMvtLUy8cH8BL2B3w/tkk8ex5+zrIFKk/PQaowKF8NE2SQ+YSKI2YZMaWxLG414kSV+Jeg1L
s6QHofcpmsBxXyyXKeKgJ9bNPCFBcHBcBwG1IdyFXMsqpSORAaWzmHH4KcfMrY5iz5XGBFL/fgR1
E9WFM9YMUM+K091pcDKFOpqNY2kQau+/PqsUusfAaIpHXGyeozGtwf99QFPEgInwjUxZpYdx/vBu
ZhBiWfwhKryoq9CnKY5gFGrRwGcB64s7G9lEJmqVgFTGMD3WajiUBdBUb+mjk0gniH40b4c/ec45
iBJCjcMM5v2ewGTcGDBfZXwmz9+LLWpho8jr1rGTbd+4EmVRa62UL/dWhrD/B0dwCri7wH85UVuh
x6bh4qLI1Xct1a1cKIQApo7vddUAuKQZF0m1n2j9tmQXVP8aO2ibYsURUcISp+72D5fpZcOgXMme
RwnZtMYb6hj3g0eoNSg1/aqzSVx+fGM92MxYNKOu+Yp32uWqAbi7NVWSM2tc48aZqtn51wJsTfzI
WnxRPU9jsxKJTIiJvrgb/DKSO47PPPZFfp8hRAoG2y51bcm7Kv7deodaeqjqFFSqbNPKwSkAJrOU
OOFILgJWWhePNcE0zghUHgpyf4wUqXIsAa5hyA2ja5fya6PTOUTUzHw1cktuQrEfGY7Q1JxV5EgT
NkctFCtHlRrfmfjrhYnmJ0HAGJ8UHJ5W4BupzyhPONuB6LmDvDUQmJz9Pi0uZaglAdchJVvsTquy
OEqgVUp5a3erOMKZg6GRnjiWQqKzUm76f+uOXbMxIToOqho9msrXljLMffxqwDLICahKIPT0eEcw
F/kU2YTCV1A7Vcu/CTS4wWsJ+dEGZ5BcCrK8Z2XYsAbvNt/EzIV+yCoK/VjkQ1ZZRiHzKLjWYxi6
tj/lpf1N/0A91k6xN024ApDQt5uezENrIARDHBEDBZebIlyIUvzP+lRV6D7AGrq50S27zcpzxNiI
/XwbtUfYmRouEn5CECEEUO8NkM+wyPNjq61VquskCliiAh43uCocBkGtJeQb2PEb0F++uy4aTcAK
NKBrWX80Bh77eiFhaOP1qvdUwMxR25rHjCd/rikhMrpjyaSCXPDGEmHjy396U5p9c55hA5bpV3M1
fcCOOPjtJ8bSHQ5AYccnNZaZBLpqbNg0hkGExf3VRw+4tLr5JMCMq3bOq1qI8zgKYY4PCNE3dLD8
vuW1L3c6thfYnIcdQBHEnnD7oKi80uZUt4pnEvi5SKh9d43oZVJ2yfA/oIz/7H7uJnWVmR61Q7yM
cFIGjnF8BarNi3XkCdND4YLrfLTu2KT31DBSHHIck41TBHBWDghmHAH0DqTqKDJjc8/jfAYuWJoc
Nh4IttA3A6e0VbTJ2VN/6W2OjTg98JJul8uzGE/XJJy08hI6pk64wGKl33+X+YkUBgau5MJxdmMp
tpDA0MJyA+zMtbsJ+TEkcuMvIa54EAQ5XsZ4i91TQtnYgyB5GunFsnqUTpCMa3NMvzzKVyY/4lF8
0L1EGkscxUWC+uRV35ziLIdjWcJTQtxDI7Dm+OrISCUZIJ4GcdthIU+3cFJNhtErhv4+nXpY/eVj
dUfPLn49mLdyy3OJi/CgK0zCIpe0IvyWL2yi8A3cO2McmQPntQRu186ZoQHAkhNy4HVKKmO4Ptzf
fXWS4c3wzrwQmOkuZTfTb8Y/f6ivfJcB2uv6aXjHB8ncr8SckuyNyjtX2PvrlwLeQuU2zFeFs/ha
u/LS2mU/4FqnbvqTT2bB7quj9BEtbVXSjsng7YhuMHDN+znbxBxxI35DkuyARtctANZv2UkFi9nF
UmbFSsapwBfmDouR5LF50En61h7EPyb1KcmAW2QAGve1BHiJgMkRA9S/PykHYulvBAZ2rVTHYi35
tUUP9uRT8PWrbKrXip8gMt1Y0i/v5NlccfKx9Kr2vMLjDYpfH6NTP2zYaGvODAMqeUsWYmfVzEaJ
JIYIMIcIEzNwQ4vPPrvFb9wbjyy8DA6ueiNe2jxabhlfofvH4NTKJfhEUfWV+5f9uxRwnuoZuJ+5
PoCSFFFytBp2ppwjzm8OsreiHHG0dIho48hnmdcyMOIZgoV4ebJxLX3VhIi2uXoDTA2Ibumodx5O
Rw4nIOzvnsp2ovnl5J4Gz39AJnkU/E/kQVeN5D9+3Rdk5MTU+2lbuNQvn6xlGzYZjJBaDH+SUKxg
0YOl8Hsmbgg3liq+c+UuCnCRdCxM8bBaSLlUGePYBJIQcq6PTVzNdTQ//JxKRviFrMh91S6Jh3W4
kMzop7qgaLAhztR7V+5wvCwV6FZapY/eutaTmXYBKsf0Ven5B2SpHEzwycDIOMZkOsNAZz5U5N/M
9t+6t5kD67c0kmdo3IzbolxkIdJayB+UYaO+CjHQ4I0qiucVJ6Mdrf9Vbub154ObTi4NadGAPFNP
YXzscpM+3XwUi2Iyp8h2O8/tRtX1IAdz6P5sYclZnNWe0rOwWN9Uecm4VMnhwc8xnJjpxrGusMKE
Het8w7LN7bbHvNXutspTDlQhbdzsbS0vRv0T27ivwOphbobEUbGzRdM4ECaXub/ZBgS49yrt/cnG
dQDGVU4xracy1Fqjf5AYXij0CK3b6fdEbFgrvZeTrCoGli1frZOxUtjJwwwqFgJEN5ITbI/kcy67
KWve1Yjg+zfMLkAWiB1DA0zdvUN5QNcH9fjqq/Lb8FmAOeNt0b3HI/1qjAFA1bkemfrmH57EOeo7
sEztwIjlgkJh4Skw8v3NSzEoh5fObYxecl1GZ9vb8g2aGuMXBBzrEO65ftxxfZmLOBzy34446dP0
lXTc/nRZXQyD+pC4U+mEywQQRw31u183at7pa2+fRxHdGBpYGJQFXvZSF/4Z8k6TMXZVoTGX/EOF
oSwVUprGp+Pu6iRAOhEW6dZlaHsvUk7bJCnR+AI0f2iaiK4GzV12bgP+QFInar/BW62MUbiJ5V5n
yO6n3wWjtNnl1uY3tbn9aTp8+UG3yB+0KTGiUDMSIFJZrqSVPOlfeHo1djhWhAPl5B2Uw7LKiPsc
L/65xmv5eWHPq5WULU9Xj5deFbBGLsEgcZKVBxhYLYLBH81vbgyV7sLyZoOw9hmKrQYvmiWa084C
FDEgN5q2eYKCfXTBhu4osqNPlb+jWfyCDkjp5BIuygyrwnjJNczODfFOqG95AEzmcq8GoL0Lm0aP
7EhMCmU0DFvv25/FegLJdG5HY7lHFPETIEPLM4BOPC4Rkxskl0JZ/JSX46OmH2jd55NrisgUBarp
pIc2ZcZ5VirHn7FXlTuODfzHmo3DcuoNVfMLKkdBV0E1cdeFGOpajmHdhu2EpnxqokvdEGyxqRTk
o0ynYCpqQ7WU8V4crSSI+t6v667EWcctIFxz7sQRjfuY2g5NHpZlMKaI8t0JTO4B03ILllvojiYa
9mY8FatcNPWRvreTLsUOws2Pq9UjFJG+F+6XBfh0FQAOw0X29WNTnA/aczCG5GTtumSsLWtfd3bz
rQ12KX0Tt02Gkxc6O7c0pGwdEAdCwkGzc1SuWCWdtFplJ/bZtu4+Iz8wgyBRsHhowVf53chyuT0C
8de2XjNVbm+RxRyMiGt1XJTj7S4VGw9Z9sOoj1589uRwLWhUCXFwsYFY8ySLvXIyoX+236kPM+X9
yokx/0EGLA7o5fOKrrPSjhDRSv8c3claHY9HZFA1Ipvr7eLLhJ3lF/KGYEKCkDz2SnVc6Vxt5Pw8
xNdgLt2QCoFWQ4H0j5VVNHQwh51mZV+JzE5QjTGE9bqubk7dfDKKTe8tJ5Inot22LqRU/tvbluW9
E1ZbkBYRA+6DSCdm5eJdawrc5yOUQiogrmUMXmuzNx0/BEuX2fMPpWcMgaAclyFBrZwflJkecr5v
JCejG9JA109Z1AhOO2PqPUs3+BB69V7pEoWMlehUyIy5T0lj0ttt+LkvIPVoE9EjefLNIvYcnyPH
w5s3cTpbkVMeHi+AG/FduMUBHtTLsYyItp6sG+5h7u5gyHsdKqb1heC7MO620qNpoQZxydDEvdry
/eC/ouroTW+cRu/ysbgn/B9qf7fYUIbENaYk8H8oPfMuuib/DxDs58KzPXPSr39kriTrjH9+dV66
NM7dqrlMhbfwPuWPw2oEkq+uIllDjSodG04PaKxttM9e+mjd0FxAopZPLO6ahWOn06WtYB0yUunI
p76vMyP/u2zu5gBelOgWzu5U8t/dymnFSZDHwUzkoTGpWcYVOid3bR8WX9fDsTZpVhTOKeSyX+lW
NkuDuovQ7sl5mVfa0ZGTEC9YwEu4KjAcK7FemtU0GtUEN7HhqL3SI5v/jQRBevd9Z+HoztlMj0mx
kFGmEEVVq3mtFqykd4lCcywEs6O0hLZbjlpDL902bRHah9EfkhaspfUcwRlKLuRsqzRNtQE4OxHr
RJTpMChE8l4G1R5xdZ5338RTruqGy/JLVS+2QL1w9apf5mnjjbMh8ia0EffhteEnfgu6B3YOiyEY
h3kPE5REdDBHZbcnxDH6sj3iSdi68hKBNL6cKjqyhjRnnZ+vbbOkwBdvIiBbt7vtqwZri1c0tJ8G
/u/iEJq+zAMqnppi8oxBW+RddqHUJi8hc7NCM5LRZOFXGvy+2Q8yU2yFWaP/ECNNn3rzJ312xaaz
r6gpmfK93BAJH/nbFfIWqQAwcGiaC8i2YxQTqYqEnrir/VlMW5ak3cQIsnUC8G1i5R1w/923Hp10
MC5/mjBYlcs/DKoGC0hBloWOO5wgIRpIhVP/HcT0yRUXUR909v0Ag1ldKtFzD4/zLVrsn9wqRonW
lg3DgzKWUOLaTklLW5Cg9I9ENBXDNs4LwjMWvcBwwM52LZ4OKgbMHjDUZ5Ey/8QOZL1cAPCfpEiz
WhkSTeuQEEQsgmIuEOjCmjgU28F2n/OwmPK4i3wFVypot/9DssJu23sgnIzblSR+yAfHBSuy4IdW
6Waqg6wBiKQG54ypIFFgZeUwZZsGXh0rim9QiyWQIqn70jq2++3UAhTL6bihNbSlzMSgZEC+beHX
onJDe1NhAQtuB3RAG+IhlhZvzg9RybQn4kCnkhII3eprmxQYZOcqujJM44WqibZ9nPkwUUa+UeRk
FCyaqFIA2iOt4u30uahuyRuqJTx/ELhwRC0Qj8eLAJf8niPCpN76Ah7WE83bu5ibseDM4tv2iKMj
l2RLseUrJW35WsIsk2qrHBap0vabLQrx9QrVsN+sEMmYE8hPdOTPqsDi8iwDVoBuNOexYANvSBgs
PuGoLY7JBpvDmVhdu5squLGsVFTYTJm24eKQyZaR4BirX+yWsrRoe8GoHCGc3hE9oVyZbFk29BJS
UWjYZrf0GwVU02Ks+QdNGK5bHFiLnsJDSpUKkh7qP8zw4Dx3Hvp439AruTDEnLbKL/eXHPBYgpG4
Lwyi+uCOSI9W7jCskuBn1FHGUTIAhomOz+nG23EoHBv/bM62QhuytnxA7VfpTOJFzTNWvauu+imd
vvPsY+o0PNRYyQOcKzH9h8QGo0MxFNA2fczm+BMGOpD37ksckE3zqFWXTyrcOjw65NqsmZYVf//H
nw2U32GEnKxGSsqYrw0D4ci44rQ+ze7hfHG+WqW2gPlKZnFIZCDsO57zhhuB/xQPePTQTphf7DUw
4ATuXtwak6ngcjUDr/5DDlXc1pxaGY16DpglE3plxj0kMVi9vfyr+yLf9C16f3XcoDTOMCpVCaBo
0uKWzU59KIqAb4MFAt8P1kcypaZqqKhJV5VRJDyVkH2ZKoFN2geHR+UOKEhujM7fgMBxSYewX9dp
/7IwsDFRsFMD4ls0sttgswk9N/JEleRqjL1x6FIqz/qVehPTHfuwRt3NOWDNqMk3eL7BgbFdaGFn
WXQxoqqCPDWB9qelbcJTOLSHS0Mzpre5dEcTtINQAJvfkKP4qEqzUAHEoSOgsIxJCN03k301x18Q
C2pKDAJTRlO9ZvGgCFVAmh9tib6k+o8luranEiY5eF++6og5lQYcB2B57T9xusWr3PoChHsDjRPJ
33XP95M1ls4zSVpWStVjG+4X9nuY2nt46NFZgu8mBjJpZxUJ78+1/Ztk9HX7SCFxBK+TZpg41sMn
SO+G2NR4zKFpPjzRA5vrt9foH48LHkux3xlLZiluE8Nelt0eOuzpkmBgRq8hLl/7x+ywXTA/G7wu
OmXUi76zlgxDacQGw97UKv2MzulHH4qXucp1ive3z1bqv7spVBhs6RwpLGo7WxvZxT+Ogn9c5Goc
2D7KsBm38qZZjNUf/tBLHlv4BuJNV9oDBcA7yr5cXoQLLRdhAhq35kM99aNJRJqskazxBhTRZulf
k39SmdviH941Pj1+Czl0UOG4kY9K0r5TH9eL6tCZsHJOQEJtWC3KzssQSnAvN7qBQsyx5wOol6JY
k07QXKcXLTKhY8AcnjANrOm/ZxB9Ju0jtH+qa5jx3ONd81KBasz06YAMEm2vJYYhcwigFEoUH6mf
bz+YY+tdGk/Re8iLbu1PLEQ7r+CZFf2IKzZxUgR8FO7XYh4polw8mjlLyOo/mjVty/oeIqNPJf2e
Jx5aOWWWJNF8u5U+qzEBOrRWDch38+Q0Gn5m7wf8u78wixdJfaTzL1bVexPc5tW/YVhyyOElcc4+
U3ctid4rLqqIKrv1YR8uoMHzACYzlR1tHqjfIzlQq1VvCvSzhkckx8eiCdDPhpb5RwdhQp5nuqmU
5rp+DBQwgPOb/hJAEqb2467q/aHtD+oex2+6WoeOc5NTP+Lf5VWfy7RMZdUJf1G1V8jzl5f9R9H2
9xeD5Imt5eA8Ozy5E5zTkUVg5QJSDinbAbe1h/+cBSkcLVb/289G40XSKqjsr8eONHk5Gk0dJmlQ
6vYIpHSxoYVE+Wq24KReeFwoiIIxqu2FCYb/3cWzoy8MoJvdHWdPkZlxL3V8gqXUmIIsFsKhoAH0
TPzvfY05YCorl8RHUjEEw/9/QRV/BY4XwmhNNW+P1cFfAJXE3QX9ofpI3s4GXSvTJf7WcfsOMYPp
lXsi/DDOA7VbN8Hz26IVI5ZeEXjKtOzMIKD3NH9qcCNHQ/M4bQAGKdaKigTlw4aUoQt+a8MUXv1q
b+zKdrlTWJsCln9dl/t4uFMEtRGo/+FPZTuNJWW5g25TU1GaXMV3ypDUUYx+Rf/i7Vmn0/NCpcm0
1h2UNv17emGhqqXL7Ewx4gDjMe0fRkM5yp2nLcGVEbEpFQhiLyaG1ju9QcDTMcpYZsjtZrXZj2To
2mqiOfb91xxW4Z8HtKtCmb9wfb1y6PvDOjESajmB7vWIRbvVImQHUqOftVkYkxSquBy3kKMLmkGl
UC1vsavzg4UqyfPExkuQTJ7zhUfiJOvaGwJoFsUK23s0PI3CXL504a8YxsZitDRrypGbxHwUh0sR
o8fDvYOVtOAW/INcmjtx8y5sFRqq2tP3gbfXqHiIiqHyDygdPqhZ+eUymIHteojOmh8ngfJQCeEY
2CXpBQjaW0zc37oETY4fKct017llxqM4IumcZRoXE+ZVAA1gWN9YXf4MX9ULQ65YY33Xwp62gXGb
ActMNYPlpvRHkL6edZUsLcusN4H5egQhmR0S/SuAeFnugIkbPRu7bcd50gq3OQu6XWDlgLVr/aPg
B35ssMQ7fcW0GvO0I5Z6yzVRLzfIVgjFwmAwTXkurmx5sW1KFSE8zCpCPjA0JdmUJLhEdyYuHDFs
/NzZc5NzLgsZXD3pCfPOXhxmreuC+8kwc+9yvivwTYhVOs+Cw11Aez2rsZdsot3AOWzejiTnE564
5IceiwRWyMi/S0moFZZ8mzptnv8DUtp607LGe/ISDFCN9/JY+fORqwDkzN2Vjf5ZMny7NhQhpfhy
qybAh1hYNsshlwCYqCUnIjtXadoSb0rbUNmo8exZLQK0lBy9H+/v4G3BLh9BedYZEW2HVzMtIzQW
IJn9+1+avtov1v8FsfTWnqWWaxgERePRWHyYySxpYc7GlnJ3/4Cj94PMyN9nabJ/0GUvof+h4fBM
2GaM1Wc65gR0GDV8McedyLy+tL1ndjBV3KmU0W79/HxOUtrgXB8GNx9omKxpS3XKkPq2JVrXhl8a
kEVxwqeLgpAsxfTF5HEu8d9LqLKanvogkZ9hr1Y3ABW0dEU8i+3kuyb9T/BuWIZVk1UETmjnIw0P
I0haDno2LZIFKthB6I7C9nw7D2kfuGcJoG4gEpuZDyTDONG2fnozTHQmsGJMEjd8YrALuQHx8N/C
ffH5+NtEOBzPc5WHhIIjicU5I5Mw6baxMDveMo+vuMoX8P1RCRMmZ4ipdzULd1OMbqJgJ/hzJMNq
S47SHwOHISwRGoH5G4YsP4loAZGGl/hUbgXBNQ2ElQNOroAVS1kM+INt7vSCuQKyF3KeeX3+TCBv
jDUy+AL1181wDCTpybrpskPa+lbaCux6OoHI4BcWGiVpv+rkghRYaP2gx6wlS93ImdlN8tFw76ec
KB4fpzKTs8zFbzLMgoIUZGytT5MY8RN8qoUUJ7L5Kh1yjUGS2vU8ZmcPe9CStsC3WY00XkN8E/N9
QUxJdHH1eA+g+6Ag5vYBFtqNUGXiSVQfPtXJL2F1fL9wTYhHBB6czpLMt3wztBSO8cEmTN3V27OR
It+oBUVAJloiJ2imCxXgsjZiFR5lcB9OBJft+FcrpQ1S4ytjpXSu2mPC50cZel4KNuHhodofx8AE
n9mdKaG6EZOLFsShtctstB066be0i3wwrEUkRLWnXR25FEJPlgfJj1tdp5T4iZEBACVHCkymYdy7
1rsuFcT2D3DYWgY3amavmTY1T2MfQb4KZreRKxSjAeJQyZUp1WMGl9EXBAf8MPU145yel+L6pG6S
uAJxwsC1QoGLW/d1iDZYECatEtu2Hcp3jRqFvQqfLYrPGbpZfg4TLi9vFRoTC/PC4/zL5xF59aoD
gUeMkkj85Tn7kMkEL1+CDV/tCVQyqehbrIEUcLYHAuSuSzVAFHLHBVpfB0CK3Lfiy7jStp0hePms
qbVkUSvFDt4rqTaHmmtyEPzU4iS2vOv2FNBFvrlBMm0DAhdLW2ESFVr7XGgRSbAds5xx9tHnELaB
VVnTGUcUJ0AFIAkFxcCy+9JiPh24YpF8yM3fan6P1W+rLktU5zb/R+Yl85WqsOtzTs9m9oZI9le7
9d9KWL1mBSaQoe3lWPxEjrKG0nfvUZFRoyi2gMin8Z1Lx74aXXlazabNtHe+J7gkQN/SkA0+7kK+
P1yHduPkRG9JBGJumw7dFYu6KAN+y9vQxLk21C/hJBIJQ1kyGSDDrZ8CltS+qbjbmgOBFlzVrtsb
Y93MQWpeMD0zas0+i5H5nOiBaurxskRMMRUwcWeQ5RQDp5GE95rmVNumSNhDa81sYbQCd1j8eh37
onzneQ4q5bnuOozv8ez6g+Q21MOQ1AgKcdQPEjHIsykuVbRb0fVt0DLouGcOYRHAg37X0GuvNWJW
uW/B1zjfsxnfHsB3YNUprdlz8xTzP8qBjyYfXhMjaF97ttrmCjQctntfZjz/Nx6qKtb6vRdDY3G+
gL0FWP9vkPYMWJjart+v/Tt9K/U4T+A6SjPIXQ2cnBsArZjU5tlKIRzywoxf8CCxQ20Qmn87bKQ8
+Ad5SpXZ6iZ3+WQDi09MAQeIJdOH9nmy75xUau3yn/5QKkBIrsw03AnmsH++A8Cja8qQU/15tqBT
PhSe7tiSO8PNkoub6fyZugOsqApSEVFUF5hnN6qIgU0dGpuYWjoVn35lsWVJn4Bj5sRTIAFyM/vN
4EGzc93GKt0+0CNrABUVWkllRDMhyD0B0Kipl2Xl+PKdL9uvgbgZSMChoqC1Q95eFfyFPHIBkon8
ja5D+i++c1PBI49VWw64zJxx2fatv5jxafUT5iK1PPcAIHeLQFGMZZlL4YdAbmWFBiyfpC9HivWk
iyO4/2uSos8iL4f6Ua0vMZpKCsAIMs8s22g4jeNxoXwWwmJ7PsowOAAZsHOIAvdfWqXuNqzVj3zL
1xm8du7QVEAV1RnLdbJDxSdCLa7WAtc9RaKVx+p6v/45yzS9a5NOkNn8WE+HLkXtOjJ1/qvGpvK8
V2rHGQMJaBGZOBJSncwsOeghYDT1YoZnj+0Vc2BSZmAwmm3UgXXTxBoa+9BQ0isZPCBqspDdtXZ1
X4fAif+b4nwLUOkujlJnoa6a3LpNkWvNVzzsniE1g0uys+H2Vn4wAfg8g2EPKCJ+WitA6gW249HB
hUBIPtKvqsUu1j2zOQvLJgxLuN9QSRFBk8P8/SqMKJ8S5hIJk6Do6v91DG4oRUw/jZ8L8QGxjs+o
RyzQQYH5N7nD/Lnm7hKEJghsyeTqMmm/7Iee7+K3N7UsDWwYjs9mMQ1VRBXwNeUDvuWZLkNEFEr1
cMDis4DqF76F9yDQB8DFOX2UTLSjl7AC0dE0k0+WCao4frs0DgZOHhh7imYpSNWdF+i1GoA9oMkf
9pgRVv4AipgWNBd7Y66XNfRxXTQWdWn9XsYUoJOLYolvryy6yMFaZONoO3+IQynlKLjU5B/jILbl
Kr1ExMC59BFLDzUtz6ZVEe8sjFb/hIfNPvOOclLqojjE8fe5bg7thXixNEmJdsdJo+IwUHqgBxVz
rW6nE9kyKaE9f5aKCMrA70A64szfunajh4fb38RBz2kQ06j+8RxQZVabrHIdwO/z2jVqOV9i5j5x
DL5NnZG+T5sARPodf3JG1j77RNV74Zbw5KrdBjIr1igafmB2QkpMETPPKb2t9i5prAGOyXla/3/0
s+XP19PbQodQuZRtuZZJI7H6NMHCGA5hAwinMLUDLGvhqvsrCypxBVUcn9OEXWwD90bJ2qbmL3q4
eOX17s0Bl1/k7O0Uzn1uMLEBgdiOPsM4CArYFlmoZMbaNaJ6VD+4I//cJ+1MZCpS/JWLigxNuc+7
G3ATq2YPUDlt7RfiJifq/pc5lepdWxaRr7bD0Gszw3Z7Lzwe1TiOwWwmF60fOIu8Bb2kSoeRla6X
t746DeiV0XqWSsc5tx1DduBJ+p+jSRRzGQwpwIfygJZ4EzGXVy/E44wohUlUWUUYXOUFikZOpd0d
X0xnorLJCU5vMnT4OqdeefAPtlma7IEDbTpazh0Mko2TzxsWW0HIVYoXLtwov2gYwSPxAX2TMetY
PfjC2ZlloVyraG3SvORJ6sET0JkI/svzPFKMwkS3fSxIfORDDuThAx9rHfch2/3ttnqhf2FqnBjv
Ud335svzNgtv+v29JJ2dncdMAjLcBDIwKPd4u1fZWaQy4AfwJNKbZKfo2fqNqtsmMilPWkfyzWKc
Jc1XVgyULm2SKnd26sNwQh4fLh9s7oz168s+fd21E/k+dL77ldd60R1yXCmDxb16MO1s0Rc1Gewz
VcheJKw4+Ud/M3/uZgnrua/kEbw16NEBIRxyk+a8DziMPC9F5Buk03xs3s2XkENI+q82ERhp6FDT
B7fcO9tDvtv8F5/hMqYNifzkC/6lqDbLHAdit3UB2e3xpuTMCGcnHTiu//qUGD/qtLUEhmcP8JNS
XKcgLzk5SSgbSffTFvegUMfFROkwa17swGijUefnlsv3ItlBQhZ54rok9GcWhr5zDwJQ5LqLG+pm
UF2AJ0SykdALb/jCuynKTUPFR0yZYU3SXbTdxhqbivFGDoSouQ58PplZZu0b5IRlaLmN0kmAQHmC
u99VRkvh58zQXTu6pZXHzu+5uCdUNJqSMMrUmjr8qYkL2CiBCe5+d6jWfgM6/ankpOmoJc1cS9Jq
WRcUBcedPv9OWCaU5s8YxNgwxWhnL8IvgTkZ3HngkShkwloMtCx0LCr2VgT6TCXPlP2f+6X6Cwwh
aaIFdfUEwB9FeocvlyjCWX4stoUKdzA6ZPf7PnIxd87t9mKgK3Yilr1PCoG88NC4CfCUJf+RyIkm
RK7bbVv3aTJhG1VPa7Ij9AqMLzne761a5OMuLz9I1v+tD9NMLlknE5qs+ZKyy3yYNa0C1Y4wpyGT
Mgm3jH7n0HuLyIKGJY2x3CdoJC+y0c0e73ijhOXvwvaYdJLGkxQUIyj8luImyVHSbPJVtXhPYyEf
vUlaG2Cgi/UwHMUoQVgiTOYKl6aczNPLG1ikwUozy7EQ5IO5AtA3pRmVbqAFPfSxWMD2+wOcU+hF
nKEO55lauuUx+um6q5rWpzkdxbdxAaJ5hkmJx+2rWldZERIqJlpdtjawya1Cvc1WYW0dxXrzvgFt
ZCqyvYXIAHYvfb2xyA3czpLQdVfRc5WfDj4nTPOrvGw2Nq/Yaw+7dkS/mmtDFSc4OMEcc0b13OvM
D3hfKk3TiVCA1AAQeyuCeiKvgedPy8fvCD0fLSPQO+nxeTzQ7F9rdq/3r9lY8EDLKTnHhVNet+Ae
c6zWXnqXegh8sx2Kpa/VOebK7qrHDmwgPiB8bBM38Urf4n3fxOaiuXBs/Lzo5JHb8q6g0dVKR37g
bBTfRKWWQPSFc8LwfDfEQYMy7AgiI2ewrjqdflGSieuTzP8whNRwF1lXJ+MSF49pjE4qIgtxS6ff
Aj/g1UhQu1TwmTuKOd1kHdmMnD5lj/9mjVrGGPMN3qoRyexQj/ptAOC2Be/uZmp7JXNEIxoMgXBQ
cHlCnmMJeMALC9iP0JMHrTkplU7J64CY/fZ70UL4fc3PSdPi9jSrF8l46z6Ynl7IZcb+tvrnXhns
3egN3FhriDxKkAbmz16IH/JDwPl9SMFJNbMUc5ZGFB2YUuU5TIy0x1sQm9ALzkcUsg9CRDsghMBH
GwAICo9Rz2nF5EifCRO/Jjosp4pfB0ZFdzjl9jC0kPF95G1O55TgNBoT1k3cQWa1W4E6VcUdBA3c
HC27bvHU5G9PMFyDbX41ygm70W3Z1s2z5m8s6Y+pxsLd1Fw3H4fFjEpU6p0cOS/Wtl0wU9LtoBXz
uFFuUQZEoGh7xH9xIT/JaQUns72J2WSRz35tXaMTNtG+S8bPmIfnyB207KY57ebD278pspEJyb6T
OrUpxDhxrw6IoR8X787rDlDMq5kH/X4VWETMfDqifsietW5dVGRAXFGEZuIMm9eeND8G7xneDhpi
gL/OJkkxupul32Kc42yl5B3rVVcDjQdDto+9yPkOWZtd3eHG0jCQMPqXWpR3ZAz2X0KrVf/vRcAr
FtHNWJYUbP+eCnHJXjqAj4H25Gh2FFfTHi+6n0X+YEBa1KLNXuVcZo+6/lVBJBK4/8ZVJyIP4KrY
Cmh/s2c5buI8lm2lZQgtBuV8fvlRuBMv1l7ZCs4QAGC0GHAmqwCwFP455UmripYg1CSkbEoj0fQN
v5l12e8r6oQYFTdxejR22TeouOk+BRBMrdWCm0HPfbs6kt/i4lBYytH4GY4mGPtgtDLcGUTBSCAj
ORHQrnHhvG0/KVidqEx6+WbVF8DJcmW0xCcSdmJhV+6nX3lH//jVeQOOK1MmVs2YKocezmYasQ+o
6jZl6X5pX924dW4QKW1Z/grGxeBHXx/BAiz2yt0Zo24UiozTtmwXfm77oOnWg1HDj/SHL22Vtb87
Nip7n+Aono+0yjMV5wI7k7X2XcQA9TFXmIxXb8WPpzolNxgHG6fojXhr7pHheO9DIDmbT5IL05jI
JZyW4SOyyAh91SN5GK7FeCQmGmwXskGL/kapQTbZVNC1GK2MTjotQiBE1rQqNoW55zQi1VAjv9S8
Zx8Wpjzk0EsZeOAGQGKXczr8r0hwgjfom3M+ShZ9WrHQ+AEKKhep/nvXiy+zuq9TCO6WBvEx5ZyL
GOjzt5C9i2ZSBGAi5XQB6jE2D4cq8H7+O1efVK0EipFB//DIu0jguh1t3i1ri8JVASAjyfCFn8IA
EsJfxYf3Cf9OQ76hQJXGYq9GVEfWYbFpbRZZKysfiEiGbj6o46pufQBFos1/Ueq5+1Exkld4dsEz
ayf32+X6k4W7xS0kb3HkXF9+fJtKMXXpLljyz/GQULvTqeqCBh+Tr4VHly/nJLfDhqWRq/41PYRM
79mMXFZUFlJ7ROl1Pnon6gDoMB1ZKcludAkG5p2LWhQ2cLk96cczyhwJBC5QAmK6/QtNid7j/dH6
d0qGemvpQVttwVPw3Rc42t7UHCuT6ckmCHb/ubTeQts4fskmslZ19zQjMzuSKiiw8bm3X7WYkhJP
hVwe+Wikles1kB3ZNBpsIRe8rktoIwjid8jj7m674c7w7UsH4NSuF7u1fHiV1TAI8tgzJ1WWwy15
gYdfdMIBLR92T+fHbocqSR7QFC4UhJKHj09X3Q82fEVvlGzyJ31m34e41nMb3mNQ/Ng4r2CyVeLh
gbHvFcBxI+W3hh63oWJca96CI1xbQ8Vi7eHh7qmpfUpfAQR1XqMmnRV4NLqJFDhCDrUJicwvq6Su
3eeVhakSmtTqB4aPwGrDNL5HgVIRkSnwf0nmRBQkqMSpFJ/RX2YKQq8OthO7CLJFlr5cQoq6vVMU
WQzE4LciuAu3Smnsc9CmGlKYoh5ttAQh59AU1PvE+iHvRLlDEFf7S/2v1IGxRAVpNbxHA6tBbykU
V8DZiJCTNs0cccl2IX2dhAWWil95868o4hIFCmRNmcFYjEs7PsyVckNKDfzrCa9dQ2cKj+IW8dR2
s6gT3QxxWnYdRY1TnfNxrWvOfYJFPy4seEJ8T3Yz15aMXh9l13bsseXDhmOdgBqqJwZ01KLeZ8jF
61snPtUOuShIXW/iXWLt7CgRU3bA+8mpDA7FT/ckCnBhtU1is7jHqJvtXPH225WTICj+ZfhAA6k5
FoTy3DiZ/j89OKODgy3a/v9+C/kLXCTn0PzMmAIYsgesACeWH3PWMu76wTbcj5pscrFLZeTjUKS+
4PnObz6RltVul/+2RiVWRPj/2A0qIJIXKlZwjr/rg9AcuNPlip0G+h6OcB8SkgFKf0oxAlc/+TOy
/TLo4Lnor23R7xt4SXFKTHYNOJ2eC37sMx5rUCB/bkx4EkPVGxkSDY+d0645fsCirdkG6bGf5LW/
/c44G42p58L9yJXc7AB49TxY0hjrNMVYO5HC/qzep/RTqycrD2YmDjKFOTT0Yn9Arup/U6awYppe
frAU1ZFXbcqI3MB9Uhwgh12oFdcBj3pmRHwgctH63CpIzB4U9yzYPlBlBxvJdwT4IGYOD+BoEld2
Ih4F6zMfOMhSaBIiGsNl2bk9KYfvMjNt6eRq5L+aAIPkC0OwKfZTH8yaxWg7oCSeXD+wZBkQbjDY
tBHU/mKyiPt9GpTD3CyYT+FbvQpDtPN1arcj4Xf7icz/C4j8pKNgDSME+PP6958kLoeQrpVNExGA
xBNi7RQ8ZEdIi8r9jsU6hbgnZtPlGomgUzIW7JouOFiYQt1O1mOjguiYSGN8ZhqdOVrG56VbMnDU
xY41/Kk09izOSjan7BMYpMHLtwcknAkYvMqK68MdOD9c/lXzDHq4OtGv7Cm4rhhGL/3fWDX5rDlf
1ef9QDskvfl4qqf3D1Ur5I1Hrse1UdTSZPISsh0UNRgzvELgOhxTsSX3lbT804l87NNWcbSizxL8
PouUd/UWW3oJH1OHMFhI2Em9IuRqMdiU/Exl6xVcCTO1sFvPQ/eYFCsJM45QpWIdeGLBXUckusAx
302MUo8QspqOUHb8HYBftzspMEJA8w/0ZyDiZl5/fMNqAEjCG7x5dtmuajfl0t0mxZcKXSesIXaw
ejgBctfZQiMH7ip72XQXM4i6JzQw0pPsRBiQEj6Pv7/Ax203oE4ftkosiJFDwcrgVQuPEj5RoRKZ
qMU9U1Jz32tlK5pS0hvBNnJt+HHdoxzGFXTUkiUO6ipbmJDJ13BZQKp0HVI58n57BREuJWFTZOQA
2wkXOz26XKii9zJXiPUBOMZqcDTdal5CfybU655b0oHoFn4ouJEOga7v7mUpLyAAX89g8/oT/jcq
hmEor9V2B9EgDZKkbLP1SAUbdEEnwV7HBE5LeSbJW8lAg8vGh5V3yjidRvQgzUKkKWt3fPedFOzY
HTDu/qlTawH9Eq6kghWOlXMjSkqxsDjQNQOvcjon6wCGnAw9aI/+m/ordwHev4SincX4DZIpJeeh
sSd77WxZUy0eyhwpgCBBmw0pcG7zImRvVb/lTxaM6j88gdrqkURU0wuf0XaRL9LU10Kszr4PLOTN
BxdcSSIE39M1dUmBBSOBkGfs9tsEqtareAiFE55JkiANfoo5BqwOYa1rl/O3zPIUxKmOHfiC50M0
SlYkVruxpV/4lmjpfhOsnWIdkhwmjyw9/yOKDirWOkdj/Zx4gJzRIBgi4VEVs+rHo9YGoJVSYdnk
1KLSpTPnKD40uTvtgE/GbFv+Sr6pyJQkXMWwAodkrovXanN7gYWlZVytYGwPnIeMWzwXYrIJcFEo
KhjtvAarib0/watKR//AccMZoEpAqIUMbjcJ3QW57Cr6lHmSrLez7Rd6YUUGpsmcWx9LW4WBiUL+
F6G0rhfd5pfydVIE4YZk3YDEob9Y9MNLhngj9G+f5N1U83NcVhl1aLB6tj80tKr2fS9RQowvIrPr
MJHFCjtByXWXOJWhZlSdP7CbZizJaEd0MaZX6dI4q5BgTWLDfYEHFwcUQu8vLDjZS7Qlp/Hf0l0r
60nti/mTxJ4o/bIxtz2QPa62wF4tTEMR7lXFnYeWWl8ZeSl7MVUfkwExbsVcAC278RCYPWNBlTNT
CfOsIhcJtmodA0GFl6m3OV97exZHoI9W14p3WXtXLKAtch8nJXlsTSEadziAYSlN+zErVbKHSTlX
0L9Wm+5211OoT3uPwDdN2wDDRu3cD/VE5rRdboqc2m2fMAhFl/NaIqMkKfvZIdF8PZg01t4igNKC
cbHHrTKsQnN9C/W86q5vQGgvBOMZpyM73SD9NxQotU74MmRP+36av/O3z9P34anUQdt1TBZn13Z0
JsBRpy4Rr95kXliq448tlP5dbF1pApR9dnNqHRZyZ/xZ4XFH2E59lLDZQ7zwBqxTHA2mTE7BGJhm
FeFarDRKkwoWfPzO90xWtS/TED455Wm0kX2C0X4FObJLNWIZwRNLHehDwxBrirovXPATJ85bMOQW
gUa9v4yo680xqcPtxSPolbS8QL3ak2OsDSFvqVvMr5uGXQ+pgTJ+u8pK15lw7HIS1eCSTSrFRJto
AJ1oTtBv1He+d9A6zQFT4Xzwqeem1nT+a5sfEg4OSXgRgth8/AwJRZrLeQWjcPCpIv9HXk0a1bNu
ioZJZqYvW6C2ubfYia8zV+rnciHEMu6x6IPFfMVd5G3XFkdpglSb81aEctbl5MIZKc9aEaHlUb86
N7/uzTN8YsEFZhTrEG/s1uTjWUE7Ps0taCZgDaQiap2rxMOiL7PPnWe/BZScNBGEIC78RRq0KTx7
oWWpK248mK1fdH++K/RurbkcWGKOpPWg4p3x2263c7smgFpvC7nHKsbMUGwKif6wj8Ef8outV543
1UV3f23v4t44/lwQoHBGNG74OuYiWTzAFWNFs5NQ0nHo1owIMnyUzEFlfRRjHqAYxL81oX8YLtGb
VIaE7YtiMqCpxF9Qw5OORNSMXtP6wetRT801BvjhP3Hc2PjPw/XaIFQKlW6T0XFEjCDFNVOdH7Cz
aEm19P8Vv6XaoRaNB2IU//XPZi/pGnTfdxgRm3XIjUMnlbcAIV7njEQKRola6V8ikfcGZGajxp0I
yLu+A91u4OWpJofphfmr9CS7m9L3oRUWSxzw+ShEUVqwsPb/MPaGitHD00PPMNA862JtZgt8+RJ1
6YjzOQYRDiGOorpsdOCvtj5qAUDDe9DVjhs/arcGPTfh2YQDVBERpBWppYfv9JLwYweT7pa3hxGz
AabPyI+giLZWWUBLwPPC0fXb9G8EFBxLOfdyugQGXMQH3JFNOAfVq4PQdTeT0cX219194eQm9OWW
olAttqC1vNGwYqJKh1IcWlyvDymy2rpOD2yrls3K8IkOj1fYOwr/l/e1U19J5EVaJdIX+uBvrLCk
DZO22jbxRONj0cUkZ+3g2mGXZDKNvnvO1tjQicI4Q1kABUH9N5niHVfZCpLXr/9Fp0DNohTpvVpi
n1TYBKZthNnn0/R3CT/wvZbbX0MUuCJAypanM/CshMmRnQmIn3Nig+haiCs0gie0d+dOpgNCVt1c
MNt0nj6qfPobbImVlGGH37TElGjd6lnzsnNRLC7qiLSNH8wH2sfMzcykOlRScu5KY4Q504xC/OJ7
VpB5lG/a5ujLmkrRf8PkCA9HIWqseqnm5ME5KvtrIViAPbbqOp46T8UcqEgnkH082vM7KoZMXKUb
ZiNf+pRT/XiE/IY5vW1mFk9XpgPZLmQ1zdLgdT8SfbmI8Rg9LlzW8wEUafg7ZCwai/wT0LDc/Z5+
KuD8qVIMSPHefhzBSKx/bIeWIvLz6FDsmOBnBZrXTzdOlnjpEXVXpIzOfyv1ZBODq+QqgIifk5AT
Q3a81SL+MqMCPzFvjImXZs6vOq4SVK84nq1JvyndYXRWt8vYkmnxMDjqFinJhZbxiR2t3ykl+W7e
OcWA6IU1pZDptQ7HCvgu63YtFoK3vs+SMfjNiCtEN4ilKfeO6jVUtGujFVlNIDenxrRvyFUPZca0
L++fpuE9Et4gVrMdFQ/4wMWGIr/A+4IkmtpRxhV7tKZK0EUfM7ZsgI+7HVBmq0tm+i1R2LyjrgIr
/6jKsKz6pG1Oayp1U3JHUUzQH4Njj7lHmdbIvEnbNqzpIsRf8SgTL55zGp35no8vHgcDW1+8AOTl
46WAqJ9e4zEogC3P4KYQTAqNbi2s6qV3JH9x1SvOGjD7EjLWoIJ30P1owX5jGmeXhsK83aKvYi22
NXOU5B2BRT8bQ868AhT+c/CWPWs1jPuRkdbRZDFt5k9ufjH5aLkUXhjLtQ3jThfA74NZG4MeLN8F
naqmy7wk48rv/2vnvJYGk5NfT/+DVxe/hIQ4wsJW84U31p1Hq/fCQTsA9UfGaKfHKE+ISRoQ6k7k
uBonv6od95HCfIamlJBWujAVGCFMwmbujIFDYtCBps+5csMy/SjZ/MPctqR2tIjUqxwXUtcTdU8a
re4Hq2ZQehg7/2HawNr9Yi1oJbpdPIxdh+QPetoUC5ZKL3ZRiqi/c1LmZ1S7uQ/DN9morFyz4/ww
Ew7/B2vUfev8tVwDeL26NkdmUSawqadD8gQ8LwF2s4aXBwBtvcyAcKs+nARLS5Fu5M4AYW/UxeKg
rZ4/4jJT6uPyTB4LuKNSqyxKiFKPW8Iiz1yC5pXtJ3cLHrd1KOWf7iLQyqHm/CZElviMGBLDZRpo
oVLVJhKIW3CqNOQ3RjBjYTyFLLLki3jvHwC89lcODeGUUlLcU7mcI2Lxm41v5CmMOO1HTNOBpC3L
7ilJoJIorOvFGf8sPVaKjlQ3oLtra/+sEUtbT0Y8lG4dQ3I6lrRnfoRgx+7PgQ5H52lHqKP+MtPO
V8cUDvUemeryzgc77mNaLfyFw9ZK+7CfaPSv2ndVugsvCrw33oniMPp6uz+08F/wicPlN9hXNe/j
cs64o+HmoEWEIRDmbKuVRtTY8eJ2CYOKWMI1O0Hb5ovCP9OM/DX/w3upz96F3Jb0WMtWV538zVkX
0SejvbFnCUP3lsH+sIXsSUPkXnmAsSCWN4kq8BIDVGgfF25oca4/mBaqfKxM1Ptt8iQYyQCWq5Ws
kF6z5F5fIdQQKjXa4nrR4rwx9ARG+kM8Gg8m5Pl2PV0+NYY2Te8j660ueqpJANvVA7FMS0MpbmzR
Gxm8p930sydtLrjLhKfVDO9AFOWY5EQUKsU+ca13DOPXuAzVnDENXD281KiSSQiJoMz07BOY6Gjn
0C4ZcAY3JriAVj8Ur4oZfs6TvVIqnOA0Id5EAguNK9lMSH7zZZcWA0smafJxeudPJyLQM86yk4u5
cK3ns5H3Ro+ZkdC1KwixUf4uqVPpjj/TfQtEdxojrZix1S8yPE3rOC0oLf+W2vRjHwhvjtZ6xIbg
/szK3yA+Cw2IqsNKLFI2c+U+pK8l+HpUyW46rO3d1sxpMunDHQC1qL7dcaxYk+ObThrmJznviRuY
q4D6PPepMoA7kVeObvIz3ixOYsTtJPMDdXan8KwhXPEVXg4oyValyQH81JdriXiC00YIdIWbsbH9
eqb5M1gpddGRSXLeCCOp84sOjEa2K3JPlbLtMpvSNlTx9BX5kC5Kyl6o+9zxrDPd6qCIyHvB4ng9
RYsQABSc4zBIfQuSmNwTGZK053O8FqDeNLEKm+9ENyVZVLYvsfis+TdPdAkCtIfiBHWA/zF62EHM
xc/1IlS7cisc7JHWadt9b1RBccvvkwDZUKTcRdXUxs9CyjBpe15W5R7CXgpf8Ba0FqwCzkVRqn7L
nDWhkv99q/MK0VCYqrY06Vr35SmNUkWb0WezvSuok8REKQdJJ+aWDVvsEq/y4LxNe1USWI2LPh4g
m8sLHUdm2TcWe5h0AnvClmCP3P0Md1SzfNX0uSUBu21/7x2Xx5FlBRqnnibn3ds7QU7TMPAyhWR1
tj57j34fEK3z8DElOWQcKfln86DVULPz/H3ZKFus8cGQUyUyNGQcILeOg2JdNjBBH4NuLW1VumvS
rO0Q0hA2qe8ohKtgjPCVgfgDJ5Fd+d20b3V5L+D91Vzfj6oksOhI7ohNbqnhW6QPXbf72MPqUBN9
6n4gKpeOhNNbXbmbtmkrftOqZLL/BB2GRzePP2Dllyh4xrYOsDXVKuTAO7bxJztshFjZtyBamlXI
fmNc0gyFKlArzP+UpaRcxNnAceBdd34U01WGed/jp4hfmwCDFkqqXvtaEELOXKmhHeFQflPyc2E1
amu0EChKaCmXik1rtoUSlm1GpF0a8z+U+dKeWFRoY/UMiCNXiLqNJx9IsSQdol06y9usm+RRtzBm
4EDXefIx2Q9iAcqHAwNWCWepvE3sxI55lUas4p5Vg0a0WSPNMP9x6jvedZ/AJjjd/0x/YHn/fstj
3mU65WxqUGuNJScLZ6isduByhvmY9HJ7dwaGDwTCAOdag3WmMaANMt+quTs5uIzn09yXQs1FisiP
V2o1wgJ1dyYGHBZZWS0MO3LU5VLTFplNlajZTR9E5gmlYIswoGSpaSa9LeNRDZaxJ0J9+6nHApsh
Ds4rWkURcUdpOxgDYivEpPbgcSI+e/L/o2DqTbJlDQUYBr3vr3MMdNesOiYreT8EJrdt3R8qsrVw
Rviv3VVB39SZbbZmB0wk3d6Ok378HA5dl7s9odEWy1agmHmrqzVK5A/xAG5umGZmeCQ/r6plzugS
+iuIJf0N4Ig8uWB3W76I4hj9nLFEFmLL9V0Xy1fCG3GpglDw5c4v/uUOnW0+sGodXsSs2DXeqjMT
+xU4UKrU9SbusyUEDPfL39VK0WfQwGvM49GsKVAP7SQfGdXc1Lqv85Ll6NqbKtR99QVsrtdCM4Mm
Twt+yULqfa0JUswuy0DnX3sbtgzPaDzMIleaSmtWfLpbasAkxthE/EmF9FDKpRWhGhu+pE68rVrQ
LrhZiBwXTIciWnbkxqSSN5Vlux1tfDGTwYFbRtCYH2dTL/kmaqukw0Me3B/s1KLcHcs2uxTp53qw
Cf9eXzjwZNZnb+hEIKQuKJHl8xRgCJcIMh+V9oKnXsAlirgXoTPSb1kNvvWeSanvlgS1OArVFvY+
Bd2LPi/lZaWpveluV5PC908GEylU9X8AziQbkspjLjrvY6KpA7Z6p0jZSAtbct2M40p0uPEHHzHs
CKUfbm8rwxcOysfAckuVkIYCIjr/OyKNLNEqMAdCx98+v0xEkk8DIbpEzM3M1Uvzh9oMHdeibStW
Rh7hhSIhoDZxe0NHeoc5gHzLwKMRcBRKz8yvaRr0WwKUmxixvmLNEQbu4UwO7yKQgyRXH9B9SIa6
yoauqQO3VQ6iMQecH4NXuihrQ8sPXQdorb2lfNkr1IB8BupfQ1slCbKK1r7SkmBRDEjH8DwUnI0t
xpVpmrtPvDZsCNFM1g1MLAxm+W3yI5kLdiB6ubfYlbLtrNLBzI9CbMbw50GTocWFTj7S7uS2+S7q
Ucwm38kwNSaTv7ctPYRbULokhWdDLXVMiV8oIHJ7jhxDPlcU/VI1HtgCQ/C3niyhCKBKmIdMUvWq
Wx8RPVLqAug1Aa4XsYoS9iovQoQhgNeiq5NJhhjtPi5+0Yl5f/uaI0hQB8tIRjSX5jY1+Rh7OIAb
e9XQiYE4tei5dFnJMncK/B3BCoP8FuD+nrQ9NRsMgJalAPEPUR2nnSilzUv5VQ0HXqOSAOVxMHDF
YrD3Adb2ysrbcj//7WtKsRRRA8RCJOat5KBnp2HU2NsV1155zXoAjh85Xd8sR8I92h+WcUx/LuD/
JNlS3TMPI9QO57DyecgD5JkysLCnj9rN2d6mdKXkYbmoA5AZd6D8KwC1dEvmojkzS4d0K9nID/hI
hZvfm8SqVxzAw/IjjzSy173UQ2jawIHoYZ5VechFMzubuIqdFAzW949UAC/BqRrCJKo4Q5UWoqVX
IWfnw9HkCYOQ9r8BUC7cS0voUG0KQPs/p+EUmfWHchou2rOdTbC/NSE/+d7fJgIaFdFqM9/40sEm
Eb5k/eyq9MCx/NiG4O5cPJxhU0hNzRioAaKKk+twKhni1r0xrfZsOOUHqL0V12IbzAUROIgkF3DC
vzXGb8P8ZIJP251GVRUVTHE4ARX0ZSnaQujjOP9/NSFNKIb74EuMNXopqtRORDjMH4eUpNBqtyEw
fBKGL4Op96ofQNBRhoxc0vVMXfqnADFIG01aNGdEa7RnGFFSh52/fi9muqNsCV+stMKecF5NHT4H
GAcGN9OaW/8TKu2AKK9eH7Ku2XsI/qEYnrfPiOqycZ8iGwKMsi4UnNmcvhiHhU7NMpUuS5Qqeebz
awRa1+OxWtgN3j5zNDhpqUGt8lO89rspck6JJggJcaZQwuhEHnsZSEeDxxK7gf9G37JYpoTezEnF
7atmGpvOGLKnf0lxWrjpNNo50f2yyQRmpSFDqoNAOHk4qE9z8eS8CPGP+f+WM/QOstSSdE6t94U3
Z3MbeRTz0R3ZcYx/Fes02P1tf8olgHe+Zr234UhiTYXmxgqM+l1/yN6v+X9WOnMF9N8TUPY1q5fl
S5emdoKHjHP9ceIPw6Kz795U5PRwILBWeKPU3Da/en09uNULJEbRgHNUzi2mbhketszQcafAd7u6
aCv7l7Pka8vfjsy/fLRmoT+u/J4gc5eYV10aKkhuUoXdyNtqGEsuefx5LxmCejoJbB3LFvKu6EKd
QLoEQEXaw6MoD4DMizepY7Rn8Q1j8FvpeR1Blmynp8tnUM0PLhYQsNhDlLKP46ri6jMF5hYxNJxq
PaRKtuFYFMwPGImpglD/5aGssHwW+xrwEIVipJUdD/kwqYC3HYcsx494I3aaC13MDSSpSXmOlBLX
fPH2p25OSDy7fljP7tEZYpY+HkZqgkRpQIzLhjporoix4qaquFg0wVjyg1ztUV1NTu+Bv/BCKkqb
9CxVs1FjyDokbyS+D/vYh0cmfvPR/HFuklGPHWrov90degz73CiBUqbazDj6S+IlwDqjRlv9QQG6
G5/56jiDK1LJsuHXk4fsfgJnVM9tZo7jDbU2NBoh/gKLyUK5P6Wq5Uxdr+z6XBILMMeQAQ+E/pUb
Kt376tZk6z/gQ1CE+uVXsA95vL/AdMZQHvBeCTPx86v6lFFWBJecx/o4aAkIXph9qYObP4nWhdnx
fU0fE6l90+qjrKb5gzMP29LjR55c51bEyQJJc/zO3kl5FThT7DIJKbQe+luQKrt4JP9J3pSW4k03
qR6mOKQFeclgHkDoJYLuNov5SqrSEwu/qoaZZ8x3PRN01WFXBgz1vuMVzsvBMMtcvy7QkS/wbvDk
dwlvFLWeY2i9hrZAQzaa7DH5687NWWljurUa7AXlPB3kJpEjKvi2dnAAnGRE+fjfWbLowpFtYbY6
0OWZC2Gia2PVC9jiz+CqsXCGxXRqZLT9w6kDRLshnWStf9BcSkxtGx63OpOq8DnGsC+ughTb5BlG
CSZCwJx+Vqbylyp10iS7OXNOhSHy2blF9y0RXRDKG0vKQXpS+Ixd0s1hIEpzJG3WtMv8TUduUXDi
St6zsdLJ05OJ0tCLmoOwKuwKYnyRLrpnuWeEaQbW7zWMYIEz8oHGCIdCEFWh8mWRNrra8jp1JQyN
yTW5oyJN1uHp2Kmdx1IW2+LSyp4ohZDaTC1hdioOcI+Bbhph1AvRfwT27bQNGqVLKu750Kd8h0x5
5fsCTttuKUoZusZrJoCkW+7Dtnlcb1P/pl3WbhJiffdcocIHDPlzigdK6x0nGnvEiF0m5FACsQS1
dJ7iShFoqcqjbuECnxuaHgBeMrSD3BRE9BIEothZy3+d7CQLn+J4BXBPhBgAsA+BPwCTkHj/fG/k
0BiTNsNCCfGgbS1GvKjlIH/syA4ptvjFiPeYzrLHtyBUNc8SIM2y500zvbQsr+UPteC5/XOz7w7k
jX8Iknmh84ad05LAdu2On/2NRq3CW5Z3kiz6Et6AHY1bcL7/fkFTvPUoyVH3DHKp08Xu+4cz1QXM
FZJJvG0xKdl7cIhhqkCw8jd4wMz5BwhCYwhF8t/Og3nL9Ih6R8A5+LqYKYm5Aco177LclAnR/x2F
NiB39ZBzJfFkCYdOetLd++GSiNgVm7XNSotL4xQuTLRMZqdLRKdYJ96ukMZs1mN4EJqILyzMHWY9
Xn/Bl/hK1zCk9SD4kkEI3c50JTrERMpWsEOlvUV4EWrSPeLSeazH8Bt+ultY0NA79tuA519l02Ki
b7fdsMi0h5E109S/1mMusyJ9kMZb+Kw4auJCqngK8S6VDYtCuktjwjN/JWKVB3llTRTDDMD3bJFg
gqHA9jPFbt5VxhAIQBMoEZSDpEXjVd61cGkM2qC6gwA+XK4UdDuVTtWwxuCuY6M9GebC4UVdGjga
Az0P+yvNfAzfSQad0w3mfrpAoXZqzJLj+54YR88fLCw/ag2vnc08FfpnwIq5N5rBb7keriyM8OQT
Ga6KKroCq7Ze4ztHx0F9FnIfosWeWroJGk4udUM9JYf1POohEAZI0sLuDEKvOeyoJ6eqlMmZ9SKS
xmynjVm7APR6ZAzdOvSMz5kUbW5CUfldAS+k2jPwgGJ9TtmDBqarZfqk/hIl7/iVtNIyEc3vItaO
AycvpVtnkPGP9HaY/3uoCMSBRdXiACsHX5nym5bsnjxt41GEazHSLsTXTBNpIdHoVj69IuEbbhZu
e2kIgZnwl9sr6bdksyhCYPYrOFmO3gxNnK89Lx8UN0SMFXcBAVPQQFij9HDMmtbFh/cEIdk9BBIN
y0u4d8OoG9l7YbUv3LPoTSq8tJDf4tNsurEIRn/XnYbhCOd2zVYZgrrrJT/AXqjIr/9Zs3q6ECPx
Mpt5ynz7vcNCBEqYzj5jUdkaGU3ZTsBkuXO+UN1b6VU1paL5Pm2lWFVHmih3VSyQM+QlvKX2hVel
f0Q0rkl3MiNSZN93ZMVuLchuPSQnzejU8wkdRPcLXKcO3SVf7P5fk07Ycrjv1QoI76JnxB6FJohe
ftT+BKHaEWVAjwSB+cKonOxBpWVyZ/8aZ2fwY8X0EMbnV1B4pACSgdMbDVCBh44J6BTFYQc0MD/g
CMYkXDpFLFySaL0AWrnwPab880kEy037L/5em1ua+YyU/2d1u8CYaOKde7r0iGYdBYrIDXCF4z21
DSd3eSzzbPFT8G2DyHMWP6rv9JiFjrillKHIoBd50vLlRNqVOZbcwaEjNPiy12IcMEEwLehPUmyP
wkepHnv4MrOHMLlAr2jJXLU1dK7ueXLIIO0agOJUlCpa7/rmH+NbckIx1Vgu9Z4mxhXXwVMdEQQ6
tRqs+Aydh+fiHunxLx848Y7a6Vos0VbV2auulorG/ElaNzb8RK9GZJr+4tPEVF61fpkTI1qIBQ2S
En3K64ezyDizbYsIkXXpWFy/2rqrXdzVyXv7S3aPLjGKwiyOLB2e2djbTSYKEsAOWkKDA7Zi8R17
Ergv0bXjM8PZ4w20gZmFB3ijQ7hOYXUYSBeHWwG7RLQ2LoFsfw/H5/dI/DSI2CIaMEQcT5RkHnwo
mBz2FRQBD3e0EOxmJdVTq2Lnqv+R9ptO5m2XL4QYyhpS0rJPbn/jqLb+qbfYFiZISIb0OZw1AFZ1
F/ryNpBAbDcFjMxVt9k88/2zhgFrdor44fTnF2jvX7WzKx+xf6wQVZs2XQ+8nFSA/nP8mQ8cGdMy
O0sQAEMOkEoVCXHc4bUp1wAtLtOyEAsb0L6nQoMUxm1/V+9KN3TrzXdPGFuzxmGgaGFqlzWbRQC9
65Fkw39YQW9D1XS5Az7lbKPSqztOGsCUJhyB74Cn9frVFZ6+vV1Bi+RERTE2j+3MonYho3eIkjol
1EH6u28wrUQRiUpTYiaSuT70pk0/gmokDe1C1JPakn9PhZO9Op5+dvQNhGbUo/K+X9DhjukPywii
pqkHVXgFLzLWmjHJ/XRFJVGwE1RX3/wfec/uKm89X4YXGkQ0tcpn1VmOvxjtpVRycmyA4mrzZH+1
tpOmHGa+L8HVJMJYNartiqnzIi/tnEJ7etztIzuKkDtbnG+FetnlSuGft6Mmcn/zeiC6Xd17Z1Hu
zHHlrUrSgztTQrXvOwpwzSgmQC5q705WrBwegFV6obipOsNe3YQmgKEDoRCggBwfyiar1Yy24dE9
5PZlmDZx8ufnxCew3tAl5MvhiETjac3DT2aHy8SD4rxVK4TEs93Dl0v/8lW3Y6LhneFvEeKqD4V3
MHRBrR0lku7svDjKa63a3uRpULD0/KCc0j9OzYfhb4EC4vh/74vTfYVnf/4ThWZEDNuPSnALFXGN
Pxw1NJdfpHfm5c1D8eqGpO5oMKTrBSCHWw5gHI8lHb7j1vUnwMd64JENcYLE/dGaynBHGgUsYq/a
LZBCY6gNY8bbpdf4KZs2PsvuqO3aHw0++v6yNxLRB8jRdZZI3PRfGzouy2fo5LlKyTSpBQW/bC6g
4wNsamcfhZnjZG96OQqBcA0FfB6g6rDkIFxLWpwK8rF71WrJ2yKlTjKKelk4LFfBKM5KGAkUP8Bo
di3Degg4uU09Jf+7FLPfk8XmjTnmtoH1ibU3fe5X0sSHSlqNklI1KK15nYMKTwJqUp/bkqlVqpcj
Uu0KGO4P7oWVY4ycaulXDIw6DUlS2LOAL6TLqgTePwgiXxiRGldYm2lINY1MDtl8El3JJFmK03tZ
X2dXUk+1vtWZ3N84c+YiqzjDwIjBbCjF41aHZ/3XjKr6aXJj/1Kso4SmIF7d/6RkhDvZ/i9jTIbX
IuluQX4Q8EalO75QGX7ZQjS+y7kgilRaY8k72JS7G25fyKM9ZS0llmTYO9PnHBBbDNv2tmzvDmzw
Y3scwU/d9e3ce9wWOqYrrQbrDjP4FtrQG9ljTMOjeSDxcO9QEgOhGZ62S48/LKyIS4sf3bvKp0dR
zy/q+TZv9zt3zrRbg/otRk6oKx2mX6REJqIsgbJYAJAMGrxm1Wwblutuffqq6QIF8ruMwklv2fBq
AC2PeTfpX/aaguxl+W+8v/vZsRzsk22wFAVKpM63fkvctCHmf0kW0jSBx1ZH8ViARcdC4fH73Slw
oagVvr036SskovUM8WyLyZ5TCbPSxPySNBFxUcm109VPehV3dN0zmWZXgOYEo2zhajQXtBbpc8CM
Nut55u9OEMcSS1FcsTxuf0OCjvLbGq97ajY3xjKXTmbiYm58SNaIQLUZCtwEyWJMm7crA/9fi8yL
/7nAtq8f9KtTfwJIHxdABHIOH6sN3xkyN01W+omj5DN+rjzJaoUSc7JkBazlenfDGlLjyMaGyQqQ
MGNQKgJlmezFtsX4wLXwBNE8zBRUWaMKE0Ni9XvvAf25TzYkAzdhzL7/NJhCzy/7+43fQtkPmnjj
DxoGroi4ta2QBzoDV+5YofjhVrqazLadEOYcc5iEvJnLag8NDp3IiyK4H+IhOtcNRBqZPPFSZZXy
SP60NC5p39UzSgvoK9RM59zQEQasCAXEpxtbxuHK+ASR4bH/N7qFaIIBzRvIxLN2wZpAc7m7qlsZ
O6L+/vsAqBvMO+KZ2Z595MlRlYU/Z9iJMi8sbtApuq7PvGWYsQaMe5RxGZe1jucJz2/9bDtX6RdZ
VA/VeDS3C6XFbAIaTS9JBdR+nR85fJCu378guopCzEB/xdvCF44tbuXohcLHd8EDskDOpJKiFo3w
VJbYi+JBZAdMK6O80LC1W+GNWoKuxyMV7/CxF2Pi5ah6N9HlWjImGwtkTVifPyOpkPSrZf/brrog
3F8pc63xuS/U3n6DxtzrYjzwCCrv6p3Hw4E9HoITpy09e9AN1XysylVOjnBNcPkRBU5q55g2qCkk
6oUNsj4mMt1M0hdthmUogDC5dim8Er6HlKa6T1P97WBrQx2OqZwxJ65WvFVFpOmZZ4srLW2+JwKc
2QGwfgMOk3cVv4+Emg7xkeF/f6G3eUI1SJ8EXqHRtfEQnptdW5rTR0s/Gs/Rz5HRK6+p365w2Lpi
h929ixA+nRbG7HfmtW0QFrI1D2bj0JouIpUIH5tj+lUt/XCy2oCVcLR8RMiRvmCaXdpXuFlKs2bk
5T4S/m48ORZWZvkbSU/Vin+8uldPvMq33nK7cmwdSCkLMk5lwZ5bZsf3lFwrjwaiUe8m694raSMX
G49B5NL7kcJlpY2oF2b86Gngzy8lcqYHgXQvxVy+L3BZPT+RQgVVslhhUYvtL/nFfumXiHBNmY2K
OF3iCAVxxUz4iA9ak+/xYZvMVz+HZ85Ae1GWK5ofP/QJFmrQQ3/QOhtBwcHTM1nQzmsGq1DdsVRI
IM0Ej4Aw51/QverEOWRFm7I7RQFr4EjlQSwc5IK45pnVK/JVS3O62+P6VXQrEvBrLfpWNXjZfcRM
kOcqq7ug2yEB0F2Tl8BDO5xFp0/Wdsn47Fi4WeYvUhif7DtMlOwSt8yi7q6/YZfuN4LNQKcF5/P0
fHzDAWyTDKjAzFiMUXup/K2rOrNcC5u2ZwZiOHTMBJBW99iSTpNpzRcPJUy8ucbfkoFrNeiDWSeC
jSr9mUefJ0g78Gi2KsscGvoxouxz2LLyDTMTIRKGZBzWHF+vaDBsEcS64/NVxAmSyJvVgli4XQyc
hM1OKEYEdcQmrGlRGHS5ay9c707DBERNzjJvZ3lGVdKNxzRCGtz/RvoQxwtFyMBhJ67P4AyUnte+
29R6FGCiY7xCu1M9TwBIaErq/jOLpJ1oIK4VWKSQUUvrfXS4bFmnzJrRPEcHOF7w37Nagmdjznb4
1LldOoo6YxlAaS3j5vIIDTrLRrChpgKkp/MfRwgy11c4GVjo86Sfn3HHHx2H/yuDlHvB4D7aOhXR
EiUP208lOj/GKarWpcZkTJcewWtYOXirvagNPxqC6jCbwqePfiAklLErMwHVtBqaMSnKw+2S1no2
cpzq5c/GMUyt/PXNEp5A3ckys2B+Vyvn7oyYnkBuIOuLOxYL9otbEgqsKtMf74kg+BhzvMgO5dzJ
4t0erRQkjg+rzrhMtYfjOLdsDi32kiAySGVn9D3z3IhsTliGFqGFwZrCiXwkbCZxQqvAqape0zUp
m1XAcBsYkiH3A+9wYWXti892zErIR3wFTQf050Wc2BOghXByPjOuPoXy5q57GyqG8ER0cI/zrGu8
vXFl70szvoXikN8Y7NLY96/5ewkHmz/0PPewJPCRqenQMc1HuSkiHDO/dSjYwHcqZujsLvKqbHbv
rYtE1g9xMXRVS0mf2GRio+F08U/PHEdms/5C9L4Q8hyHdZwH2nfxqOyZDpZspwJlhfpVWxAmbjT0
8syaRdjfFVRhqotaJEBsK5YZX4tmk5ZuHnQe/7djfUA9PhnfDTvs0QDcUoqfcNwCc+YpFEsCwYcY
DpPIdtmEpEfF+ArOWtQuD4HUW2sxLt1zgKIu+mwNpcPwZ4FBggGD6YyP+hQQ6XE/Fspxb8uMEgVY
CYzAwlozW1RQGYli/L+N8YzbzARQq2pSp9nu5f5L68zqk62INKKFyOwlG00Cw6YDD57j+o2/LKRS
Bjc5MPxxMrEkQP0X8gqdMke0Pvf9KCyLxO3spg/6LYINwos+lzfYokXVRfoYeZeUEGh7Xot1g7sJ
KuqNeWD7gBTm97gWaXyhhxWET966lh0ljks241dHnJ1mTd1M7cr/ixoXgJm+aIzS5Zoha8OqC9qN
QN1JrZeYJbJ2RRlaJpMDtBJgOOP5EgI/yr65HbJg4KtSg9aNPEBsv50t4lWO/xyHlLjimYMTH1ns
nSumPz263PKOClUUhbgk5riMj71md5lLLbp/xO7488ge3dPxAIYWvyMBAKvaJ+0hdA/qz49tJFt3
g019zGj0zpjIxN6OWu3sfnNHKhCYRTfuFJvihcZCDlS1QIvvhiQY2MOSqScgrRqGyRFG4FaEOIWZ
cWfGoiOc9CIMe9dvXB5zN4z/UuQlovhl5Z1wvFHi4kKTh/eEcp7zfj4J1Wz4rz75SGa4pFgiIXmN
ccKvuRnc9DrFlXjaBNMY5cTbMnkmXrNetB8GKFo8f2cAuVeNjeO4EB2WQf5YxhIiKKzu4L226EDO
et5osJEclx/onTWxzRXHDX/Kma7uhAvA5QcaSh3JJSmt7StweDKh6EgIXP/3nzSaplCecXlVa90t
ulYVczkufIce/cAI9+Wj1eIWCtpph7ux8l6NCRFJWZ7lYn9EjTXOynTLeTFnj3Cpf/zwRWw49W1I
dY3GMFZ1j8DxySqfrP8/7woYe/RvXKLNIL1V7FLFskrf8m5j5Ehi453/0tLxnuimKjHK602iq0q5
DhiLeB7iNhMGYf+KyesuPGWUiV7C/E+dpFS0M90P3fMeEtDPkv1m3WunO6zqhMQM4ceq4XdSQN+a
l0F+HUGgnCuT40WsG5jvGsZcmTX1vBMyZJ0SiyOLXxDr+vppGS1dIOh9q5LafbLLJCU9OFwxxjn3
ugugfmyKeWlTDzDhswnloguWdPpCPEkZRgTFTrUlgx0W5nWDbAa5YHlOlMtO0teUIce9d7Yqm8yC
d8PTUKxPa9f68vUGvSlhxPrKJ8iyMgnzamKHy4y/iQl9GaoACCDoAZKLbol+v0nqioUbhmjrxMCK
+ya+7AIR50luwVq0me6QGBzbsieCCN/1FM3wcAbOl/h3gJEW8RafKA3FZUzclgrQxw3D2q/3t7Qr
EGbm4s7E/jUokQHXJGWYkLOtJUZDrNeDpHmShSrkF/p20DpSM1bJ2QomkOzGfOi/TTDxgZL55r3e
RNMKMIW54rGsNLZJKG8W25ikuntBovc7wDi4WeuwYGdvUIVENeilsECWnLgWM8MifKgXQcJ4Gheb
RgB2RlhRMptTbyC4EjfdxjmTEKctqqtPlLs6Z+LT8miaM/Lt3vZVj9wevgDcSAMHwp3AEpG7EyJE
OR9WUURgon2unQLCHULTG0OfqxeUA8xgt3R+bbQCZabxQaJKb6KG4uxpsdpRF5b3ZyhcBHCLJSPx
KAmFPZlF8P3lX+Qx6mTDVNHxfSSHPhLRTaV/ZbrTf4ns1v2qhVU1fSBl8Kbhm4We5lGe0CumlBXo
Bk/CRCCAMJv6ZeMLUL86U8wz9PQnZmasF0JO06znkA2LBJ4v+WxgLZeAFW2D6OpvdwZkWmNrBNvX
Y5TiiFBp22RJ2XRWOeYjXzdqfs9DAoSB8KSuGGoxViKfrl2ZFRUH834e9C1eA/a3YwRhFd01RMP0
m8VkmSB+mw/5SgytUgGJBFBtlUjfpa9cUEpisAhD6uSwFeXx0/mKUL26rj9i1aDlTEXoifUJXxKP
nsVyy7MEVxYRDYVAoc88phDcCIoqcVN60q6TMTSW5X5sg8PHLjME3Uu6t+y3Fa66yIfcAPcyb2YI
m9RFWMcHxO21gDe2jH2HyL8Y5bRmyTUvrAZASzQUG/MOYc0XsDowcdWhaHy+6dUNMoeYdbDqhph+
bpzJWsiF4Qh4q0LD828Tg54TX7hcCJnb/3R/5C/GsPoUU5I+jWjPSZOWjvpKWIa3YoBEot8tuMzI
fbDwCH1m52GpkH/Z0G+2vuuyuYbJIuwN/mfxHMz2lorLGd8p6SnK3s7ZZ6XWtupLiyAjzrWmvuKj
J5Fk+uZTVAcy9js85VSkcu/jibdUngo2Xbc9smnQncjBU1A4sCNMzLtjEhtW0Zyj8IP9EJoOIP07
UzrBkkTnv0kGKVBe4Uy983/05icdqm5JFr+VJt5bfo3M4o+a2O8XyAlk7cbKtpMG9u6Sv4INv8Hc
WFiQWfwq75HB/kFQfwx+ChxQdu53mSNa49TfWxS8NtOSy4c79Xa/sEtzgM3TvpnPNENOZZ4f9CLC
xD4DWFWlPbn6xMHROAMv1NmZKiUK63wHEavoKEUASrGjZfQ75c/M1ITwz6qcD76e6GbsDuNrWP6A
2Ffcg1NxpVsEBdftW8Cuujl4pbZzAf5M0nGTKZ843cukR/4IMwvrjnCK6Bpw9MC6A3uTlTzQ8JM1
tH6TquuzqzTZPvW6bY4w9XVn+/8F/laqwb1OxmaNRQuoWXiDB5CpNZR7HJY2AXrVHgqGtdezJJgg
gVCGSq0FtTeoC+cR3ygSt+kJQSye1/TiKLWAW1L9FTC6nA4ZhuP8sz6uGFUI/xnOo/qLlbaFTemi
O25KwjjXcb0lmdvw52FMvDlvq3XufW+UQ93eQInZAHIiRCkzcr5FNDew6AWN2iCZQDfmSROBpwfh
n88jMuvfDS0NLmVLsdf17jprxTrMRyVKE0pAUTeRK45++mgbnYb9QZWTrcSOZnueZTQ3/69DHaiY
gKw+LCFJKo7DM1BiC8BZ912xmwQDDtlo+bFRnordmq747Fem8uhRMaemlgTDAAJvdJhr4NR8chb8
MS7xel1mxrNp5TcybdYZF+VXK8u9isFrKBQMISN86tkSgYIAJas5taDM5GmE+vlJF2+c9tj6s9y4
EsVGmzbrNw2CgVf0ZzYvebQQjwRSx161VXSMaIrzRdGIBvzYA/4izFB6JbGHemAtTcWO1qa3khBp
qQOxFLq2rI1uM2Bie/ym0vLL2nQcdO5KyYDJWI9BwW2ITvvxaroNmHc2CCKLyoXnv2CREQ2x2WgU
PQiX535W6phTnyHqMtnjn3Q8eBy0bFkMrcnAoJsSD2f8SjZiWDItQbKASx17UhI/ssNrIxOfykSi
JSPCoXmS9nLolozbEp3nTfQuDEFbo1azIOPw+VoDcFlVWCDFp85jlkmCWOMsWOv/fwlk6xpJGrf6
5EOrEArTWPwiEPposavSTslYazGMkfBN51V+ReOjpYrz3+fkOTdeOsWXyoOLbV3FrLy+THnHw28Y
kVInM5l2ryp5OfGyHMLMtWaouitpJdWAWaTjwIi5htc6uNwBXq1PphbaiEKLX/t90ZgVjLbgAmnE
qdRAZLcU2j/D7iwmhM9Se3BcMPLkKY0So7Duzis8G7bS+Xw4TCLn1GQsm573rNhLg/pEOIGtdVK4
k4yhjLN3VdWtcbZTKsS+jPSdPeR+LaqkkfceuCuXBRFap/pvZ1Qk60XdFBykHFiCFnUouy84zZ61
elef2wbCASDeqtQllzTqNgwPwomxXngxyInsrlLwr1xJPYFeMxLtFWr9jf1UsP+p/7dvum1KiZU5
3Xo9QNlKROTp8X+hqk/hf1W7my3yppG750WJ7KQ/zmdwn31rFd2VU5F1sdp6TL0NFLuhlB4j+/bw
j44xBZC3rixYYRBNE3vPzkqOHgVMkvsQehPrSMLWl+N8bxh401jmcnxJ77xaFMMPE3+jBcC7a7Cz
grIccgRsvFo5Riq+fEDlRigwTmz1HUbNawLOajEoph1XQBGV6HIZsePPkDyzRl8LnXT9xsMJLEgH
aQs6wm9nsi6X5CxiIDUxjEpg3NHqy8JWEcsjcNf+gtf7qY4PazuCtjGiNl2sV7uwFgepLbEWkKss
mXZr18ggIyO4AMimxbCPchico00tD+FstvZxrraHL4O05Kaw6OEU7dAHMN3vjnxlCeJvm7hnRaDA
wbcFQ6OHWGax78QHw8MceuGaY1TxTRizZimEa8+HJRu8x0GANFzcEsb+tn8E6yg0WXfZcM2ipWDF
CnQzIb5HuGHgPUkSAmrvK2DJyJN4XIz4ln6OwuLNgoDPdv2WWSK4cLiCZAo0akXW9f8CDbWk9+Dw
ZjeazDNAnP9qCmRLIHEMpiPdfjUtRD3KtSoBIO0Vsgv5RyIY6XW192n0ZOQeuBZJEqLNt6i1B2RZ
mcce14O3xaMKRrzoTU/CYI8c63vtXdMhmTeOc8exkMZT1QBNwEruqOLgfE2c2mSvuPlhO1P1yOfb
NOjwUB7WqCTkwjXfHYGsugiC3kykxAWVh+N35z2kKhOyZXvpA2CLH2ELQ7s5KRxe60O85LTglNGe
RhMIC8pDz7ZawDurvkCADg9tN6gpdStlFc6AUTfHBxz3IjGx4Epmz9kwu3Kq4kWo6MS/ED6RxsAw
MYL8WnXHgyfCItvLjBr5++DZ+UepN+ebPi3wjZrTzmSSJ/fOJFKExHsKiXMTIaOeOOL5+nkjLAFI
fmE+gpokqZgEehWfeE+8q/Xt07fodwoojilkzT3aFgIGx5s2j4tG6PT2wQ13AX7mr3EKClhLtrCw
UG1Sww9X5qzhwMZz00JgPrCBeslDF2z8InDy9wmeXwcgA2RA06O73ZPQ0reUf+EpeK9y5poJYzht
mZuB+e30Ju+/6C7BlI/avi1iYXuUgHQz5N2LRsgd1jCKsoCTBFtPcLM07CsVRPjsMgleQlA+EOKf
m2ONCBiIxRBorazVQbDX4nzANimRxz2RRA14gXBO0MAqpoIL3f0BqEg2o1nP4kfFskgFjIOIQFeI
Ld352vOvkwrdYN35iEHiYOw3pe9OYtJGwVmHnnYBqWNz3NiPhciNq+W/uPNkda2ukxGJYjYe4Pd4
px1ijHXfeUezvEkte0ZV2iATVST1bBDg5pWf5FtEwcg1R95h1bmetzLGCmy1blADSxwfS4/UEwuu
T7JwpvhSgBlBKAs2Ju0rshHfN24pqCd9HhMlp1L+Py/tz4kdHQ50Yr/Bxgl+HMImx5IpRmHxumYz
q0ugA7XOtryNwG4Y1GxMI/o9HwYUdWW6T88XVEDH1vBpnkzasESCWl4mpJvjoKwYft7YfDoMToWZ
U1eg9NkwO+jmQnCAmGgLFnpRrRDCMuxnWAtMF+ZpS6xqxT9GB5ZjuLFEcKLJPJpTvx5RnTokwDBw
9cwc5Nhfmqb1A3YdKsayOCeiwEyNex2ZuSjTBvIzBas4xOKqZP2ApWMZAtG78vIomfz4A4wtOtDB
hVbrUZ7qobveJyPc0jPvUU7dlzjuL49sgo4tSuT/r5GefJrVCU3yOIccCe3TJJey5vhk6MBSH1UM
scBEfaJqOXq7z8k+UcV4Qjx0QXB7msVzHEDSJ8Oa/byLgb4Nlcla7xGcSV9ogNNYuzumTLpuz48G
xoNPbjUUkClzhhQLsdvvLBsfDzT0LzopAVdZVjin9yudWW36cD/EMLvF0w53shC3YMuzqb+EYbU3
WLhR3g56zv/RmL7NKVRvsS/P+hRLCYlkuNCfgsMV6+L8/X+We35YOfWWZpEdbqxzrgzSIAIHqYtg
fvsO4BNDCzM6kzaBYlDfQ25ej8fUjN3/SxJH9nXbxn0tUz1qUyBxtbLD1xZSOrS7itrqcWj7aJE2
CtuCcLPgXEC8LLD1e1PmFy/76S33IfKYyWQq/S+UNZPalP4dOEth0C1FVH+eLE47sz2dqF82GO1q
97JAefANHMRZAKA+90nhvl0CVkESmmVlC31a44iJtcc4r7nnjitF/TSMfCJyNKEc+P0LVAUVd1+M
N+gFlpf8kWTB4szOQXkg8GqMy2dk67L514DJKBdS9dMrKIC9EwoULpy9gcxlGkk22fYChK7tCJN7
et2SifuCEM+OEUIO/iYaQHuAm5QCMyIt/ytwAZ6rgPoy1Pt00gAK2HGfVv+jUWra4HbOz4sLx9wK
f3DvAqmpMoWixIOye/lfXx/u3+bzQEJ5yW3vFuWGtvEXU7uktgZ8eoGOeVxlMR+F7Q1prFQYo3qX
CwvuWfhlEJz8Taswo0N3XSVjsDZTDQAMGDBGafUElOackzby1ePPR4Imv3Gp8+KLk1D87bCF0yPE
VLidtLsmBnzzJH//ZHFy1KzKJBWS08yIudkrVyuS2Di+AWC13fP/JvfNHuTIu4s+CULF0O1G54VR
zotVdj/rykEVe1wqUaSmL1OxhPzdxCHTH+MiVYwL9NmtWeFxwyGC8YAqwa7VLHbHWgXsQlnKNC3w
u4ZlgnOZd2O66ZfdCwfCC7SdlJtwYIJjpw78xT4d5J9rOOXAi0jLa4nPg+c2FOtujeqfFsrEykVE
W37AxOXpx4Sez+3uNaDwBlPmKbwWhf6hdcT50GnD6pXRMaPy+yi2RPyOfr/9c4smlnf/yBkC30Js
SEHHhgSuvZd44cSg4Uf0ejOvMcTJ7/2PxU2V1mTRnn4gU1/FXYoZXHcILjlsGv63JWhvovBy7ka9
HgQvbqh+Df8fb5jMFK6zFDH8vmpFbF6VfvP7fpa77fgOLX8lVRgl3OiX2xZndFp6HcZhSxch1LzM
FIXP6OR+H9MtoQQOI11SCVgB2a6bVNskgrhGDoYPWdH/liBYgAl7auAgIdfbZaDpENIsU6Wm6v7q
dMw2VNA4mDxvSWKj2jiMeHzv5suCPAdJX4XVJPdS4Byxe8RJM7fTA3N9wQc1NHvThLLi/pDuBBfb
XbkMqCw6vlJrEDsebi1jUtVYyYhUR164s9R5l5hYSoyFRK8JFf9jt8kU7msCUMCsGFlf69IZR9y5
5DGUY/YCNkNry8gtOnFD3KBaJ8M3TFCFXW2TxyHwftD0nMWO5Mtj2LeRMEUh8+J/YyN5pQWnC+ps
8RES35F3BpBb6XA5pOmMpg6R+W78yejYzTk2Wbm3q78mx8orj1ZO5pb1vJsZVuvbn3h8zLVGV1wf
qgm350drSjxvMxcgHDLxeRxQ9A7Vm/eJDjqnp/C/1P/t2ENOfINOqcZVEGBFWtUBpbNVwY4Rpa7C
Fb1WHKOvpjxGRZ0/z3dOOjcb1KPJHlvQVfFjqIZrLgjVrRlCc42hPmisg1yYAwT1U9xHMzK5ivb/
wF4ujU3srj3QYvRuRrpS8wTipyqQ6lRig8g/+ptVynllsWB3n1IRxElq0P1PspfHxaeDr/wSMGLx
5ftJzmRdzJLRVRtMt7DGfrnfYCaM8Wjgx/5We3XEukzxcb3jBzh34rz6/HCtUAE6vWfNcHksSHo+
AcURlCuFeiQMfYiQIllP1ylWq98n5UfVbGCnmn1N456yz27VAdF0damOZF3MCtOa3YM727bVc0jm
DdKNXK4Lvluub77mYC3jaS1ySvCLQGWiPE/nx/e8YUCjfT2MGTeIj6Pc2Pm3aUCqSDfKQvgCdFv/
wECBnjkWbA1UdnF+vHQbfg/k+VABn/00WP4riSHg0R3M5P8rZ5rjNrgYdWc0TnYNqvELtKtoXcF9
nzdN1wmjoOmuBz3CjBKNt7etdHtP/2tRESlcug7xaQ9HENVWoFjQQY3GD1DefvzQinB1EqOiiWBH
1NLLzXGgl4xSiJJU/Gh0STDtTz07mucKG0ujJoEwDE43VKDG+jQwdfXBJaksygl5uLmVY4z5kcJn
25X2B0koeCujPzSS9tlL2ucAS5JBgsLlgbz6Ibm+GoEOkiBU8F9azJi0xHMbDiLBmhiYgNgowge2
LVlon+UGVKTB0a6s6EbM2WgB4ZaYelXFV1mDIliZIgUHidzf4sAGmqosUsNl4R1GyO2+FMtmsgU5
rTdkM+qwDwTQ0ZelAA7ovwk8/h/MfyBbxVWiIsNelyl5HwzVNzQbyj8QMuN9p8yP4eOQpxgME+Q6
oCgp+eP5Sm+TTnyKiRRr20MoDRuJWIjcB8Kqf0RoywfFNfE2yhFd8U9jWDlDMxvfqnx4dtFfI52i
ulnq6IhrtnAvwqbc3giKy7kKQqv6TXDINOz5ccgH762HsSf5WpqCZpA+5wEny1UttLK2rjl8oidJ
21buLq42b3WDmjXMnkwVMmH2syHUkiJwGIVvIdL2r1SrLFwDp/Zk4pnexc4zLBiEA9oOBvdKsQiq
EIVEGgs/+6gSIEkGURo/MrlidM3atwJz7Bq6yiZIAONxxzw+csswcDHD90tUYUWdVyvqfSLOtwHa
bkQQijpU07OM9zY/wC1V/b2rYNG1wfcKVPKks+Z/R2U6ypATc+MoLps+/HlYvDZ4otwZ9a+Betqq
ICGnca1ocRssa6UslsYMjrMEAQQmJ8MzS6VtrqXnzuSmAsCeHM6cxh646ovrIo1ZAiuBXV4Tv+EA
plrxDcL9i/n76DU52dF6N4i5yOKkG6LXnYHb4v31TE6k2bWsuV7cxvkUYq8rikTvJmhKbE++U4EA
j3K3+mfEqgzyvIwb1DB8f/0xaDXEeKlxakKCUOBl7TECmVBpe16Ybkb43Qcx49LVi9MzSI6o0u0/
pQUNXRPfSaVBKY63GdWavDDuicum/mbXlOp0IUqgUuvCSP80XzJitgL7hc4cloFeFQ1wlbVYFbw2
c/Cs97v8JtXEDGqeRdAgHt4P9Dwz+uqx0ya9JqZVfTvHD8O2E2tw+z/fmibNOqMBEPRjQdmv6v/F
i8NZUSJBZHmG5+gIRayIALgMeZ2gwbmi8Xrdkj3fNB8rZiTRGASugpttGKVhV6G/Vcbuukqs1ww0
Gj4GAHGtiGzC0bo6ZX5mZY1bT+8WJe8zHTeqWo0Hs3H8l0t9weXhHQpaRkvjg6Waks5tvJ/eWN+7
jXhxPWNgxMGtsRRCA+1T5fQWjoQS2ow3MKVDWofZkYk5XJiNt7OmXolaukhLTonWWAjPlUlloczQ
keQjbtO1hOHmt4sut9GiO1+o+jyPWR8EuTlVr1+po05u7Gz4OFhpHAauFp+ZfJBCQdBYOQ1b/eXi
54m7ZL+mbO1UMhF9GSH3NtYGQDc6hYE6pDdarcp4ir3mv3qwWWQ4MTqH590RCVzO4757Ox9hdb4u
FZxC5sGWG3+Am6+KKW9OuRN1i9eDY6Wnf38VzvJf9EHgXfwd+4DJxn5rwsyYFoduZ7tIksfFYiiN
G5+FDevZqhemV1st/RLgvVR3IExgJ/Vv9ARBSm2LaQqrZ5ayXGvA8ZWqBmPRkyxltV4ZMFLUCoTa
rlMpVFxmYzWqEpos6uCUhUR3CYQjaYLov/yaeR4jMabXHpEg8u3PqBqpc5m8n3xysl0SOo/oou7J
jroNaMb611Q28XbmbOy539eTZ4VkFfL9oQ7EliPjPnySD1v9xL1b3c8Qc4mlp3eBxSFCTni3Olvx
+t7eBVvFn8nGiycbtmkCy8jPjQx+tTLr3Hb3JnltY8vIWJ5fO73PvyNmi9ByL6tR3pRPksqBYt9o
xrtLCJy7pRCBXPxFYynOhvTzBuVUBTiTr4WTClYjMlbIlrDCvVnRG/SE9dhL7djg6HpKXSPEvSsT
xD0/nE+k5UnKVq4OCrNkErNfrc2vvxz6vsBj7r/7rh4JPsVEEWWWXJT3uydnNEysL0oOzhibQKc3
9sqgw/aUWokDyUkbnAkOtUYafmlSO5z8RGGSYeyK1CJarmhwEEsqRhnBCo6pL5/+eAl+1B8hfvp1
1LMY1XFuM9UrW31iFlRjnonGy13nBr4h7mJRJbxD3bvgKbOMfdvTp4DaiY0H82h3sBa8MznHRSiX
12xiPTNCvZIMfQXMSjDJ5zpnFJESEOMGsjHXzBTuC0+eUQYrIrHLBFUL8AU03vi16HfhtKqGA9sZ
FzXx7wBImVi51m+aPvkyi7eqm1soBGUAsa1cIoQWeygRko7RhQmiDgYQAW9/448t+6mg+fYhcLCA
Pzr8GKtcp6WPLnjY468qRB2uzGcf3WiheIWsyFyMIQe4+Bbm/XpPTVIlae/Tx72M43R+mB3WQb3I
PpBqsjE2MCKi8rQ3WfVptoXuhpT6YDhlLX8EKb+6uK8DABb2g8IQDsWFC0JdEHuTsk/pw7zVQWbe
22QmRKAfRnpUJ0Qk5SGLjZyBw8geR0zyTOvTpBB6Ua57W7EYW3EFwAf2Q5nJVRrU7aYVmQ0Pacgz
ruFTF+n+/zQzEXIWKn6VGtUikf9JPmGifsUKvTUidDbZyREW2d6OZl4urlH40FdqtOrhEZWLR2nX
aJoHX4Cu4enAA+aGt4cQi5TrPUPld1FkWfFQpieA/L6/dh5bCa5q2S5R7UdI4eo9+c3XiXsTVEHl
60HsHOKG1EFroW2yqIrRqV1vXVLUEMRoB8ZwfrDx0hciLo/o/xmW79dFhsar1LfY0/vBw6gmW6pV
JNeFDZCNzFWqgqJGG9HEJ3N/rBMdLxm9anzBlnV/pNVv+HE/zRoB9PSyOc6W4/HnHc6e8eJuIvVD
V39p72l0d1FqT4S7q/c86KCrY8doH+DoZVt7J0Xv9ipnmvBUI6eHia7a6q68LHPP0+A3i8aobdEf
bcviwqSAA5Tnqg5i/Vf6+0GQw0OeV3BjO4JrnfBF//Gxxnhp3zB48R2yJEQjh546wGYKpih6A4fM
lyakOmqX3U9fb/SXdAeS82BT6l9x1/O24b08SixK9Std4MsD8JnK3aHprtq4+0STZYBuZmmeRYHS
Wy1+Lix84snTeNrJKUESiJmTBuRwRjHAdCQPo/MfDMB8WEJMudERll2By867yx5qXkwQwvFKZxkQ
VsvObOK1DLGCHj9tWOM13gpvcKo9pURJg5np6CJ9SZ7wOfhKRigllMi+LMmBmt7Yh/wSyCOAVnoc
oPp/X/vqhJkyqVaD17VCo3rH0NHB5at5ZioFIWFG54RBw/C+2oag+X7FLQ4CKCMP7qp9oNe+QW5H
wIqEUBqDeVh9iD3FUM+X04rB3Nd6AtZr67MOsgk2Ke+0tN3GC5U7C43kOSmSvrXNblq5rKX6eKJL
NgqrJXD8a8gHoA9aIrn93IQcYDIFqLaVsKIde3mYDDTcC9ohr7znZEL2LfcnLTE3k5X20Dujz29c
fzX2GIM3WFMI4U9iSwobqnwA30sNWJ3KZc0+fXKvxHEkUW+ebus+h2Jq5VUgUwtrfWnI0EFkHIAA
BXz3S9Bd4swultx/Fpj/ACCvxPgYap1UEY04RzAggD1QEAnq2xKXDs+8DNdDnnEOrvWslnsf0g0/
PeHeDrqMCsQ18EMEMQjPpDLQSk6ALLpke1oLG+Rr+tw6gKg4kL4Rg7G6WE8L3DYKYK7azKmMXaNu
RsVn4gnDvEKh62gEerNZMgScs1N2xQ4WvRlwYSZWYg5LoPZkwXaWVrBW4m25IROrb/QDrKfMilD/
8kdV6DdGAdjXrM++oeZXHnNRx0Gh75UcIu/f/0iyCnzLCkuNmbpqcY4O0go8OzBhd+cRjrSYc5L3
LW/Ls2eqFu1v8XznFfBB7uZQav+0w//IR4H0g3XyEDTuo25rZeK2FP50+pYBRfaOvSo0PGFK3ucZ
TLiHyHPtOvzpqauwVOfs6sMEOLUH7Op3pd5fJ+PM6S97zcQslX9xxtCRwLI8HxlP9UTXFSp+0irS
or4MTFWho64GbJnZCL9kIZaAwnnqgFEFuiAj7bqw6p9n8rK6d/szpoM64/HAAevsoEza8OjzTig1
mGmsKBzyHbmnJ+FOau9tkpOw6Ke72T4jq3G2I9b9ponivjLnU0zfsiR38R58vorxEfaN7Bg78d5z
lReQNxDj+nAiGHYDQgEfofWKIf1CDaQsyk6RuqjLFYay9vvzIzzaSHwG4sAZSBBhZh9MKsxUqV0G
lje2lU7u4Socn7cNEz/zcCm4sDpnMljAZ8rVmJJjdBTR9g33pZoY4J8nWOWWrKmLUAh5V/IGYk5t
h/LK+BFACgPUUxAWS+KvRpF4cj7fjY2HYhFNu0SAmlCCvpuY2V6ir3w8fmq/Z6uB8MVJ71vaJjHM
1QFcIm6GuVh4sd25nqM2uf84iV1/myLSoWT4i/ghTvzGO22leDDFOyEf17XSlwveOjwf4vOikQIE
eSqXEEmjrmVRyAuBUhbd2DltMc8mnWJscYA3NGaJRBUSHqOXc2sHKScsZd2E+zs8yTc8yTJ3mZ+s
il0A+oBV6U904Ndm2UP3PeHy0iVDbJbjmQGvPAkR57SpdPw8CvMKL/l02VUq6u0jWTzGLUgg4/Hh
S4gLFVBstnFGkd6k9yQdhRX2zUc5ZvS/sFcU4dpNQ7RPyywg1/vrU3Jwi5JUUAr5uUim6G3Ls9WH
22Is3MlbD/4EUHAxRLBpAIaX7hG3qRHPBU1W4v6y5YSglMZTvaDk9UZJJYod4MEL9SGJVI0Of9GR
zYuRZrOQ1fxrKor7ZhNGTmKNNkn9Q2gAi5KFYI7wsnaXDOOfTu3O+YCSb6ZwAGieV7GJ5rRqyedG
mPBmWA4WcnyG+5PZY36zKT1CZLZZIcoPA8ywKETX2F9gEtb9VABRWMtY69MrJhd14uYLHI+/ES3T
L76v/rR+BOWxdK5FTz4UZ33jYOEut3hJ203yYn+gTdVbHbP0wb5Nxs/dCGVcFUJGiA8Y4mNrlRKc
fJrZnRwnv05KLbgDda3AC0KwnOX6/vXXmXhsM+b1QXvdmO11I+2wUhRH0yODiPRn2XnUFDY94L9K
84+zZ+imA+erlIx5e2Dd1zNEI71AYjAmfNXpXA2XenCoeY2BxqrDLmFPiLrohbpYc6gM70XmMrPX
BpqUc+v76+sS4u10jjnhhWr1w2RnxUkQvpSzs8MFrFmwDGWrzPzY7fdp2qtfTOZqzJ4USOwmhyWM
tno7Hqjku5c1Lj61dOmgNQ5/To0+4nGe5zQSdIp8hFJhLQ9Wgg4zbeC6NF/CnSrWb0UVsFussHGw
5EwefwR7jPtK7RWJncgCSieDJq1NZ5JZxc/4xP4gTvGmcAWwAL6uuxgSwNLFVohQE2y+wo/jimWD
QRwyu5gQCCDSU2fDos7tzQxAobYfpqR9WXwgpu4TReFKyaV0PwaVkXAn+nusR+fF7wRqqmcWJ7t5
9SI4spuPy0x8wgB6N4P4U/dLn4UGma8Y9tqoFvG9/Op8/sq6YJJv+B/tdnjPdzEY3Ns9O0OdvhrV
NgrB8WZSyX8g/442ocmwzl286glf3MgrKaRxs6BQlwRScXL+VREeZhZC251ZZhg/vq0EV0IJXeFf
8wsI1TkH64qg9ohNSk77fFu70xp2kHcZOj7slHGzDWa0lddLIdcJSj2uLJIf2K5Cnilz1/l540kT
rQAyltpwA4cr6CBV7wSDfKaKkoCOHzofBmx/y4Y9uN3+holk8txHR2ntPeNPKHsTLxif7fQIdNNz
W6ibh3BqpeWprPQZ1LXUzRpoLIssknoqVgKUt9+xKhzTRWl+uXafJtpYsuzPGQLyrrFdTmSNenJM
k5TVFeK9su5LOJt305WJ477s274o+/FcaAGAc1OK7mz6cuYRcbbcY79DxIYU5XsU2HBNjSDutkYY
y8zFJLJ4R+PBIRLEWVwl5oGjcRoOCl3Cy8iW9xqd3p09e91CP3bzMbm4mR1kn5lc9yCXL3g/fo4b
IdT4VJLcKlBYkWb49EgvLqzf5m/AV+DgtJtqbZm/WjylCBpElyIczmSotpYbtxAQcXLNcd0ovbhi
mfin5pmOKj2l9Au8WlVetd0aZsCjf/L822sHsEFOUBLUq20HWKgusy9xf8a0ijYf7uUN+pM9xlCz
XXYOsnD0on7X+SheYLS7siXh2rnUVxmIGh/L9qLeVEZNqqEI9UyIZEqKEDTGFhAik7amEIujNM4b
jzLAYTErmF3C9XiweK4mvKSUzdBDNxIciJXoJNfYQQdZ9HnyE5hYzgiqI7ULRMqknizdZv+3qdTO
+QtHfQuPJxTBKlOYI7J9BlgOHtllsAqhMg+MeIuFpS/hn39E/J8m5YRI7og1pGsZX6eMD560Jbg6
Gc1eRg9qGwVFwz/3RwRdjIQzdOqBsQmVPt1cmC12WlV4JFwMFe9cq4Vr7jOCGsfKNEidhlmLlZqJ
LLpPGHi7ttDL0W56TKkCUgUdLIwuRG1qUHKKkZOy6wMRCUJ59P57afP7j7SQQC+g+2qjz1DnWeEr
FiGH9u+gmOxVytWQlIQFEy6bBoiOZp8S5yLhxwVo8vjhRuS3SymXNTXeXeQxh84W6w60G9liR61f
iqC62KRBaGmcO1+AwnWaAqKQ75drs8Y41dfPHlAwKsFr8mt/jKEy/dutxXnyDQAjkGPcvAk5Awys
kCkVGhkLEGcty3t2/mxOd7CmVZgz/D7KP4EjwtmL35QSga9Yjg4NXR1kU2Ye+Ju8vYoEX0vf7Yg2
xfOGXQshOUKANul9E59qEyqgbCdnt2VPV9GvutSadcQ9XGt4uzYBfUE1SFoGJpfPKSG4/zrDqyAu
+ICpLViL7Pcjo+p3N5lxHvIsAEqRNllQv557P2Jrb0LRVw9WTyLcJqURw0YQx2vhZYMZy0UNFu7u
sD8s544zbuz2YUiz1VWzCN3jmvimtHOvd5GdVDEk0x1a61kvL4JrbkQBQV9rx0fsarMPPyXyUfNw
TamHqxcckYCLTEBJFwRsASp2hKDKxOYzjPsBpXg6JYr63sf8fECxZDnKvMrNfD/VJMRknhrr0r1V
Letq9hJ+PL/IFLee8xECS94nKGFmp5RKS2fCKSe7fnZf6ZF7U/ryNYof1U34RGzY3nC15OkLZXbh
GEKlc+GeMH4KIuNpU3XJ0rU+1/znk89L9GqwkwTDQD1T8CbW/ZT7f9h0RU2Lc+RnqscnRpUj5R78
80B3ROPp8ugkzbAqH5jgsIuHpOexLr8bqtCdtWafoE+ZA2DtNP3RvVLoaav2mO4cg77qT8DwM1uM
c1zN1F/Fden0NXv3ndOGdc3BXS1GzIsB3K2xQaUN5gLvJUZkflgVXtkV5Aa5IxIZX+xlVi26B0nX
ATcHxdyrPRqsXek/NYRePHq5MFrRkBkXN+sCzbA5K3JFFqiBxK59vapusOduBFCW+xY06JhLi8S0
cLbLGeUbnZVr72TPUq+LaZ0qAQRkV0zUUl7VuUNTmHo2XXuV+LQu4mjiK6xtVhIko4MMFpEGq5hY
Jdsxqkhas0dxQWQArlx9KaijEbJVSFK7F5q2CRFC9+CM/y5YJaP9pSQi/+BoJZcgFR+8gwH4wvEW
8CGHykom6lgmFC04eHXZ6ARRR84mbbe8PJobBhH5Du3E3awxcr7L1eHeoXWSWSDXU+fmmZy+D4gD
IMn7xCbImTwKYSuQMdMAKYMz0s+CIKq0dF2KgBHovYO6tqlzeSsXn7mbA645xVM+NbL1IBzWysvd
e3n8us6A/F8mRXFHdARs0kK3A6Owg137y45mBAso8L4JTc5EZf0bNLpBHmTDSJtfMFWkYIC/JtU6
gGvo125BpUqF7YFi+qU9VgjOxyqr9wyGgVwXxNJ/BEuJRbGQ+XDbRzQTzjVPVDMwYthN3NXcPhl3
j0Bv4oFttrBWDPrQaantMSQ7SC3f0TPOOlwqbt9Ta9836n47a71P9Y5d0murqHPO0KtbhDB9cZim
+gUgspHRUYyAD0uvnTiAuLDf6PLuOOg02fdQf/9g70eNiDrWp49HBBWJWcgUX39+fQ3yALPVBASz
DkNjv50ieqRixYbrZRaYi63pPSWP25fFSOxxiceDKRyJymdL7UkI5WHaKxNeMfXmlInnQZg0bKPa
BvkOtBSjwrG1W/iG63CAuiSlw8bf7ndWy8DWhbP85OB6RQseNNqQkUM9UPhV2SCdwpZ3qnedh7gQ
+MLQ24X+IaTNfy+TVA5UAORLYtkSr0fBvksiItQJKmTXayLIFISCAjCqVlz9IExe4epymznhl+pU
3ZP3YlY28WIKQ2wOh40iv92d/Y5mYM1p95OyD58RvuYub/KcCb+Zil6obcKaq5oiStLInXiC6OKv
TJcvqF0Pz6bmZjs5ZgyxfJWsNv+LnYG2EKN6NgWoQmyoqUw1hzkbS38y+/E+tnEYM/BPaYU4Rk7f
LN9iRbylTEbcFKA4dmaCOmreJASziVw7f4G0iHJaGiYlOak/z8cUyxLEycHz9t8WyCM0gu+vH9L2
z1Cx55pOSCEjom+v9rVNN/opmd7WVMUESbjm1aVsLZCDlyy+2x/oLUxoIZhPa4I1wXvC4KnuxfXW
1j+gP4bRk72UpxK/iY/Vzcg2xl9XEWY3HDGd1kZBN7OTPa1ignxWxiHz3JyJTkUYYOJ+5tBvjj+0
4lwhTlEL8/RoWyzJUdbWUPyyJpeGitQaSF1ElG0cei1lHVVGCgZpJcwEyIl2EwT23D8mpfjSDMQD
KP4BTox4F0Z3fgWyklhvd6mc6dE4OaAdWHSqgkEn2c+Vcxn/9yp884i7mmVot1O4f5nHPAOGS8X/
4l8A8iUEsatoweSNy+UIZhDH+wDMgkH7VAk1xi4mZLG3bM2lE1fVsWjbWVky89bFF7De9THOuvxW
2WcBnP3Y5NdVtcmOU2ruhN7mcafQNG9IUfErGUq65JEaSG7YM3aXeSK4RoPB8930sN59mgce9TXW
hnbTpMtl4r+Mu2wQAr6VIsokddgRrz+fhLNUNzzb5TgwPfMWHdx7el37ZBjggR1Ar/FYOmkbZ6U2
F1QJ+x+ApqOfmoKAdRxCUi9YmQGbnvgppKSQovujvjTdkQP69ngzmhggie1/tC2zgt9DeVXraH+i
UvKwz7weyH+mATcp1pOUzue3r0gU/ckRgPSmCDaDfvQNWueYVEOeopcSB+8QYczKWzoD+nhrGQMM
lqzb713GxnCmmfuGmhVrgAHll2hpHuZGIP3IemGwwPeA7dz/576cqj+wh0F/gBHgVL9VxaBbEDx/
dn8H+qca2GRziKoixutg0els7jW6H2NiVRG+shOyL6ER8aLzuctz4ybwobez07s1YDOGAVofXrrj
bcgfHopschEeCPIn9uzFPvq1AI2sGQLu1yjsOR+ExNatSk5H6jQVLBlkTHPTE3eCRRP/Sz9OhvuQ
RVP+B+45ZamnhqO8/7z6zPvYW32F3bMXPr1HCtf8n+V42UuDG49GAruzrHitDyBdJG7zUrQQcCQr
3OO+VLQqBW9AG/12NYeFKDGPG1ClZuHlXdbtMBACikdfn0Sqzozga52cr7BE/XP/8IU/+qVxOY9Q
QC1kJomxRKwqN8tHaF7UnFIDJx5CMW0FeIFKvfyxFWsyekRgFBHsH3gBN5+I1vrXsUunelAlnFrt
Ur+BFcw+Xbna7B+Ysm3HZF4yDBSXjFkVogBTh6LOCiJDFib8Yl5ysmH5IVT/li+AqA+QJO+IWFxH
B7mJ3y9HElkcYS01gtizF1CH34+iIs7R9+XYwkGIoG8DfcPoKxTY/yJx2OB/kV2h1cjm/seErG87
+NsW6KIb6ReG3MvJAWjUeWxnU4GmNHF9Z+h3uHTCrD/SuurBRkrj+TJOBKPC5yFfJdZ0cS/vUCET
BSXzgjxNGEZJQbjWE5aUpQTCrmlL7OsDi1ekFmhBS6KvhF/7YJZkU88xEiq4DcUHfXKt51KBRXIw
7xbuYCHp8LJjp7UChlNRozyU0861eF31pHtJHz0DaZS3JfO4nX9Q5igxMgiPE6hEdZhFka+QWMkD
j85kF9D/KTksYQA0TW1eF+ftoHrWWmrxhu/6wzi+5ZOfpUkV6xMBp/BgGD3WV2NtOCT4A8audq9/
ijt5M5qyeyT0Wu3o6jRZWOilfHMxOhpQUAR3pOXOBMSqjUKso62dT9jMR/DkLteSHdvk6fgRz05O
WG+cAAoFN6xnFvaG3CgscxAQ7xpxUoBxU4DLldbxyNnf5jgyoAdMVTMwikBf1kArAlb0HNagkWuF
e1mN/locE1vheiXI4/ByJAjocuXa5oEl/FbuqoVZ00UXzoazZ50nb/jQlCh8l4kO+n+AONCPVHI1
9RjfCKPPeR8evFYY4lQDfuhQnb6yfa+xmaIZ/3BV0pJypPwMqzo2lk0a9F7P3eodjGXMzCEl+CuG
mC+/OCY+OWxbI6WtxlrFATKg7514BNySKwM0d5psNZC/8ESboBnrFRayOHRYTyrjatq62rvybll7
5RHCCZu1WdlR3MDv0Yoh5cU3xPbpJdRg6pRxD+qGC97f8pdFcK3Bkxzh4dgmICpUECxlVdPp+7XN
z9TCK4DoDLTEbh39Qhc2nQfGMHVSoJA0BcT6NMr+jjdODcJQ6yTWf0xazxjhDNUuKSCDm48/Coib
0EgAcuRFaRWaXoOYT5B9m9yKqCxe78qGe07pbpJ3yyNCFN6z0dgsJuNwdZjl8CHfvwM9IygGQafI
64nnT9xlRSN+4aMZq74zHvBFgAWQHnstZ9mivJehiwj5bNUGwZYmFJEg5byU1VYMmlp3SS/0xCdo
vVSQO5t/75hBNx3YMSH4xA2yPgbsc/XYlYji4dutv0BlE9EXsstTS6hFNQaYuD70lidGB/nty/Yy
CnfnBf6e6qpXSAKHG/z3rzpJZJmypy7TxkQ/gCJ8QN6k7UYdGsyscGuOi6vBQXdi5HdV3w82czou
60XeFsS1bQXCtxJuS/GZQCX1aISheD6TVeYw+OY3++o5r4Td4aJdnL1KFyw9ArvyqhzsmbO7YH8B
hB+OPRyjAEDlJNQhXr7V5+JYXWoAFvT+6h9cBfMtgRoJdcRmbSxyWdIYJIsY0fXDpapRkJzJKoxl
ngV2BeGVz32EQaTwLCaKOkqXznJ0cZk2nXcbkJakfPf2QzLOh+/dNSciHbnAcTj0R0QCoZn/GQ6e
KOOEpMlJc9p6I6Vd/eqI/Mc0ro/zsfFyHsZ5abgCjlnTa2obvBlG9wrQOSbtAUhVh2xLeqcDN0lx
FTihmRfHki3fyxdcy6lQ3m7IpkZPArk/hjvXqCT45k7JiyF1/DSyHdrAtYffcP6pcA+WbHKFCw7/
ljQ1u6n4KqwIqCHn08vMDJFrGmNJuLH7+AOdFqPOGIXp8nHPr5Mw6X4dWL4e34sWNoX5YkxGbjEc
4G1HyIkFFFxCdq406lqvoJPWIRsYYwj3zrYvNZVx0aYrDXaI6tj39Tre7Jgi+xXy+U2BOuFb4/NG
/nn0CmiSftdV1yyLRK9xM7brwBbusBn1HbGtmoqqhDriEKq51I6AtF3GttTMup2oIQ6mdregqVKF
BTlGhskhYGh+4oW3IVs/5rEVShbVSzRrzHPNtW5+JAChVbtm2+Rdc7TlY2BK+GwBJzFWVxu7oJX0
65sfVGWpQPYWWDMwMSuw5bo3+sRGblynUxZYVCSBfypacAjKHjou7QSH51i+VwlH1e5isSdCuuEH
974lr4Q0ikpNdPxoKsiyFEGQ0zT5a4LzIwez+96S5HOSgqlGlWUo1cW8S4O/IH+7WkqcUFnfGzas
vh6INXNYGIqHCw3ZqAtYytrtKAlo9Uigw9fygnnkI1FRxHLBu4YJ4xAJLC9COSmbhksfoC+d8mQ2
dRb+gQ9wZb3nbfz++vMayTaXjy+IKAFFPeG4SnsIdlaCAY4EfoETStqHlW7Ix3ZQXUJOMVNeE906
faHkeDoR8lV+MAvDCG2n/0uAiylsHjPfqSG4LbvHKXVQ1U/Jfjo8ha4E4Gg8PBNlHgM/tEzsnI1r
pQ4xcaWl2EdJL9iC4C2Bon2iuwCWYvMGNS33a7xnn+QNzYdjnw7MhLWQAkQo2tzi8y5QQTnysK/B
UIA9qBrGVg+G/vSZrpoClolKXKm4xgql+Fgc96csUgdOTIYJv499d4TlcvxIkLQKE/FhHWXxF4tx
qZwLbJP/xYgepS3EARxMyMelbZT5WwN/UGGTb3M2eeKtJuJAJKabqR1atlmzirYLsfeiw8Zx9Y6I
DqsyeCWrr+/af4WLGaQvpKqIT2mutdSn3DjYsV0lG5/ZiHD9mtUOrfhEM5ywx9NXihnInfAa8axw
rGBdtX2Qdhufju2V16MFDOTJcbrp1rWIBNYhQbXbSjhkfBFb2wX1tueC2WqosYNLWJrUVgDIn/qu
ywSpJGhY4ShSKRVZz4LjMSnBiGQOTZEoD4eXGk+aZlp+K7Dvi2g/FvkSJ7UhhYO7ufE3Vq4n4b74
qZvT23p454asQkdGl6r2NelupP1gMbpe5xgjEGxUu/nj/5w3BhgeFfpBP94ayjh6x/5oAKyCqAGH
62/QiYvvGp1SrVeWWR6Tsqgu+lmXSKLbfGghJsXuwSnVSka5adq42qvRHr3mRJ21lQUHFjFIf4aM
3w8c1li5oM37v2GRDmQtkdVWYY5wUOOXkGkM09cIQIIH9rBRrXI0pFdpYC88cGTMJ0R9F/havEL7
H0IOwndI3KLelJcuBdPTgwjB5Q6W2F6woy9Rd7w0rE9NUO+Q5cgKvTto2wDQnYbi7WMmt0Bbpvko
t0yfxWEuviGKlXSKVOCqbx+kUERhCyqCjSZhyEsLD/yDvRs/ozlh5tQBq/eMxZLYRwST/vR9zJy4
u/8IzbkX6mHJXgdU5SwDPxVM8OfQtKisU2paNFtD+77FXg2wdZHpCqGXui2mrylAK4w9neZH6kKI
TwuqL6IsmYKGQGygMViiwHjy6OC/1jAwgTlQ+mZCrcWMMQeLQRl7MwChpGGOh/qaUfusQb0MwM6v
0eI6MEIy9FAJWGHerFJV1ItYsfisU4lGhEQuRbWOGF0AM/kKK3/afjsThI5Xvr6ePqIwbFDCy1tP
iQm8csyfoS9f4MvQusE8gT7mksnrA9ZoRRXxNPaXIP2VCJWoV6b3WdHdZCfPh5hJ96nN1xtY/laS
qSZU5vBwNLk9R3c00FF1/twbKB5DbDhOjHsUux/J2SjB5kjrSzANNerflv7S8ZXE5lGaaUvDWyEC
5F7EwOSKmJVJJ+ewzMzCYZ8cay7TgJ/dWaeoPtdC+jEIw+AvtbrlkjyKEPnyVnq2n/qCbXpQxZM8
dsIxlfg4mSrX9yZQKXCsI0au+QhBzh2RbQE3ImwkNup0wuiHLfbtXJz+AWsWG4FwcYKsXIEH+8ww
aMqoZe82XyERKeO8tGdIQXYxyt0wFv+pFMTJn1V6is6vVMOHhAVGIrGUcRinf3/0VrXbSRSSd01Y
p21wwvoMNqoPTPt6tQN2XWK8Lt1Dg6l+z69HYLw4kd/ZQGaGzvtpzRktRVqxO4wUnbh6Gg6joZxW
DmjDsThSMh2C9mLga50NF+KipxBicUr0nWQ+wVZaromIlNaImp3U5NW2PQMcc4/hJN5oGAf9jk5G
Ho7KWnv6fnQ+eKRBzmqZ591CGuL+0vfCwm2p7X+5ege8cAKeeAFbzjpwCM0hJuOekzfNQR2zC9bF
bYdjHhJQHev7+FxL4d9oFfTCfCR/sstmzu4KG/JbNjZIXIGaa5nj2WUxfWc/CUopMpNgoYwoNCkm
ssaBdDfxHUpdIv1DZQBBMYmv5vDfgJ46JCrTDoRjvlSK/0tMtCYkuZgZ5+sVgJgleUONDq7ydjmb
yqpuq1JTtu0Og0zMMWOhX2D6krcMkkqdi6pXhXIomsSPRpw7wTn5aHP90hGIDS7IMdzNVeEdZzJS
FQVIFLL/jtrn9/059Zyj1ZLKv+G66/YiaK21YkaS+dasGIFhQKxlr2FP31svuF5xOtDXcEiedsO7
sgBnRV71+X14UDdJumo5oWVD0cKDYUlgd9IVu+bz1+naNgbUIrj09ZOLWOVr9fXTpEBwUzvTyIhi
mCBFm9EK391p4X1equrNpm4AudSN76q/Irr78xp1rDSlnuunVh5JNm9VXHZKeyCwr73tx2jdrXsy
IAULwZXy5bRO7TnhMlbPe+dkLZJ9FU3Xd6BDThmEMZ35j+OFNAytGyqxcGVMbRqAMw9TBYLKaQp4
G7afKZgQ28G+fcG+RZO4IwtzIq3cYi5ZcypJWKRe2mAU0bG0SONRiq4b3Cx3AQb6k08wFdHqjW2/
WIIzworh8g8/Z2N+0gT9B5ZXTu3+EVCLDFhACeClyfFLHZ+Kqdmcea87IPInBpxC+21sJses3bE0
q/jV7TGKKv8vG+HeKsusVQfY32jdSQSamZZXB9UlqGf/DtyC+Wv3+iblfgJReTdQloJi2GiyLbVn
/aP9xLdkqerCrlmVAZnCUmydBoIv29Q66paJ1VC/uocSgrMop6/gDiDKuIUP300NR7OmgRnhg8Dm
w3ao42grNlg/RrlGpyUE0GKnH7XSIb7+dexsGqzgnZ53zUDJaNmV5wSScYAPOEH1FH98UhQ6AOoI
Za0GCdekxl7JNz7RqtAXPndthZFPzoJi5jgPE9kIna/d3sRfSnPMHgQaBD5buMNdZQfVOj2YzUd/
6Fh1vbH0N6lXpELX53cOZXE8nfywDep0wik/XWms/Y1qLfOKksVxLYafK+JjpFRdGtfvEnMcvEmc
YccGj0F6Uopw7hOk612G03WZirxbOfr91ts0boRuvMxJZHcs9BoeQIrlOw8TB0w09P4wvkBx2UCj
u3F8ilOwq7D7hRuPqYwWJ9EBkYhek0NFvYQO/k3QYRio7vK29wFPFknTiaXDX8U9+qQxz+FYF2sM
MasEED5v2+4PrdmPQCNjNYqwhJRbdJu9NpkBud7EF4OoSUUOBlIN09q8i4/XO2uPPSIjEcMKA11S
svhTeq+aIxebKBGCvy0ebGzb07x3tZDPN0PYkkSDZYHCpIHXzo3m1HnEywni+4jK6FBc0/zscAmu
6rwAdwmi5Rei+STy3OVG7H/dMTlbBYmspK1PV+TMzmNAZr80ijsVbFgWzpYXo6SkQC31FivLx8QY
mOLc57F2UCKXmX/JZruI0XoWcmvfVchQfhXwHVfjUcnfq6iwDWNHFz5oWOrH40FUV0oF7SdtlHGW
sz1oC+c+2WTuPuYoiFGhbLqh2jISYABsMBiBJgzaXz6RC73x/dyyQwtl4n8VdQeSOwht0RXMtiHQ
niGEjGZdM3fzP51pyvLOnW9MH/3qdE4Ki0cBcx3XRrMUSOHOxqesRs7ebOwsplfBGG2GYAVAR/ff
JCs7wwc1kLSKI8dRXykymdPxVSUtYTkB3n90MhEuyKyyRq5TIR1TzA+UkYBm+Kjc4rC3s8AkMt1a
/KmXJeKG0hUhC8PggwNR+/HLUFbYLf0M36jVcGkPNIBNwoDNfbzuNDNIJGb9lQrQt5sD/A/uF3NS
C3VzosjDEYqFHsV5R1PWccx8n19T+1TOXUd3SZikQ0i7Acpq0lkgBlSxg15MJB3/NgLZALoJJDv2
XUc1mZUOtVXJ33odBwgxnzjtTk/iU5YKs4PCm0pDY3JeMiA8mVA0X57mfUBfEywFCLvvtKXip4ZJ
PIe91PDmCFHt3zi7o5RdsMo3edtUloDigMxmvAVnBOEMgaCeBReRQw42O/blpS/Jw3gDXuDP9Utq
chK8Q6Pg5MkOIsGK1Z/qPXbofU2IwRg8R5fnjgFi/CVakE+5PRaZwZnFdo43FyF/7FdmuoBDDmEF
GInMff52H7sNuMmfb+Bxgvb66/e9f1C/fUBxVl9lw0OEi6trBPEvnKbxfZKAP5pIiHloTCqAbc7w
oqWnE0M1Vr2Pb/li/j3VOFRNXq48lP9vCa2uTpMRxu0hJaTPTExSRPt9K1ILZAQJwxA3jbRV3JyO
h7Bmqu4Bz2nEn6PABYRI43Tg2NpAXf/xFrCjRxUAQrDQns27gZ/bs2d0iw8BlnJmOkgvq9BgMrq6
vxO++H3bk8miW1znJR98KIjLU9604Bn87SXedbhsGmPVB8sZMvOeC01X3+z61hdRfcYKxgbKLcIX
Os7fvVElx3EgpkBX8fbsuG6KTogyMChxittqIP/6bPo+MwxjdNhk/SBeRKLNR3KJyvzlemhlxMmf
8tvfnZ1jFhn9m8lbmaUvDTmfPOOzZ7F8WXxPAZ1kXrpX1xpSrcPEw3bq5aX25Qv2pdMDr7WylXM8
b2r+JeTAggk0MCpa0R5I4L3LGFhr9u3bC+zFt3ch9luAdoBTrdbZD8doJPyz7HaApLsbvzmzYZze
wawRU02YCgcUvHWENePeH9rdifZb7Kbzhh6u9050IUfWgFDMlnhPWzxgbxZbKr2s56zf0CwLLUGc
nzq9ZI3Jm3irxp3Le0h/d/Wd/HaTT8KjH+WK1I8ivVvY7DluZlwAqW5UfFaGdWXj00kg7WQyJT+j
uXR9NpRQU2TIRqjy7yO8ahVA18mlfM1/aYoUMobLQwL0QWn9AJ97PzfYpBxo8uyWw6MGQIjYrQwk
5M4f2g3kKP48eB05eR0ohaLznaLTw4e7L9Ll0ScPPZK7bfmiUU7zVN3Z1hyLt4GkhhLFHofAOMMS
JFVso9rqRrQ8bJzDJ+kGNy2N/jg7GscVi63IhxVGA2MNvuhOGhzPHoPufWAKR5Wh31EHHRc8ZiYT
XVfdmdXxt2b0G+Iqvchkkzef30J0mfJmpsPs+zEEH1+GhMVm5mvYJOW3+V68rthSbZi0mbQgVMLQ
VtuLODmnA+V1A/BZ93hY5k+fbKE0PvzVM/3RfKxEUaVe9XP1IpvtMgBieP983W7pHncYLFk/A3Cn
0mD0L6rPEtnLRVxbnyiJJlmdnBy7UeeU3nGrS866EDLFswI1INr6RdLWdCyrJa4Zmaeq0yGI4SdB
qFn816elSysphwF8idptj0ivYTKgNwewcA9CAsRIZY/C6UE7gEV2hIqqpueUxMMBdPu9SEvDgsHS
4W4I9YGdgc8OXkfW6J1vr7074IZTNDqmplL203Y5AEVr3H1D21uX+kLMGpfXjqzCIl2xw1sdIkw9
+5+5B4KrVrZdXoNkyRF7bFru2wrDlKEbhXyduM1Qhk2RiQ2FdJeeZIMJpcDyEvDcvj2GkEq7zHw0
DaoAkeyFVmaRAKkiiuB/po9uzhccemHvDP4MRt3p4HF3TDX9P05GrrQexi/c1YI12GNU7AXAaf6I
bh2zvh2o1k4ESW6lMkSkP0Tv22b3fnbPQP+V+xxn/agUklONFegelkCO3LireuDuAf7Xxd4GgecU
mV1fLPltWUpxikx1pjae/9Y3qiULy+BZYZy4PSpE9Rz21adrcqc3AlNBb9AJTw1cuEprMe+rv0A3
fOe97iJXFXZ6Pcy2CWRMXmuBt1SGEp0sHLDis/KrpH5yLzIyBcAUlVsgW0cbRplE298H+gnr2HlG
q3ldJPGM1HWvBLCCIoX8VMtji+jiEZ9SeYW+a56wdA0EBSG07cckS+W+lBTPWu8WtkDi0fJ4qQuY
zMGURy5MJqLu4OC5/eC1HGGSbSB3oouOxZg54eLF9tggWanK5OuLI6YwAVy/oaRsbzP09mnO2OXy
0Z2Imj/UTexcQe4UtqQPe+HdyFRTFmgsDWxQNIVMFBg9WRWTCqyR74SAaBJmTM7W+RM65yriDiIr
YkYKLM5aCiuqQDk0mJyPt8enQF44+e4hYlq01NrlJdnKDFilqE+swyLQ++AduKTM7jItxQ5xKsiR
ORaaPgilZeXvZiCmYWrI/sE+ztzZl490kqH00Jm31Xil8fze81S+hu955hzQ5kLKzMIGqN3B+NSy
q1tlNvkuXr81WWJhWJ9OYTCBJUmcBVlEbJYYtV6GKX2SdceYDjmeRs/hDFuwJ8M+5d/XgP2gBMD1
N+Qieep6pFgnhqGbG7/QtJKC0tB9AlyMsynen6OCMoXE70xGx7QB7UdzyV7T6ADAkJfI6NVOBcZr
m5BPk15l/zQfWptRn4cbj0nv94XAJUIcvhGEIwjBHVHwXCL0jgxPG2POr2titM440uMpEH7tG81H
P6b/752PLfaAQsGIQ4ehkHq5vBvOQzCeCnh7J3rWO+qL5oKZQdoLtLH6NZDvuOJnSQ/ugJZHXzzF
sy4TXDqzRfjQwnVBwWYVdK5dlkVqWB+PBLeghoyYLeMSWs5vJnxUks8HdaX5FQFSGQimv6gSISuV
TamwcAdAjtinTfPgNr8Trjb8rlzcnZ0aNqJJW1YcAPXnAnuiISH9iJlhjPGrQAO4jcWSWgbK+D8I
BRhwg4/VO/cG+l41piDnQOTCLd5Wq+1WXukPb87zvg4+0aohZdGRjCiKNFuWDsFeQCUhghNHQhzc
e/PfzqSppVmye2NhSRNbANFNlr2wMFvFMdPaYIGosjXgmMTlfeznOfokUYT8xTOpA0AttDTzjk/q
YFA62ndXVLK02KelVWQR1f1CQO35k4OXRHxJjJVPPOWnzICKaHFzOTQPXTfUA8lM1W54zzHLjrW+
EJCCJEikbP98tQL5NLlK8WIy+pjjeRy7gsWXR3ixVWqf7xfIl5+4WKxT1R0LEaPR5ThwNXIYYK15
REzJHMJeL4iajVA47zDqSK/3MPLpR8ZXse+Tdz9z+lWI+8kAzDmE2Yn0u73DxpT2HHiy/JTE41lx
9fiWb3qBlmJJQwXEKM17r6tkjPxLHyHTrwzAURHcyCm5myP4/SohGV4J4mKML+kaEZl4QKB8P43Y
8fnV3Ul9Dy4aLpZR0+bHh6ns/8TYOs0/zeuTmn88txGMJV1luvXC1sD3SdTGXd/OJuHzqTbgu2ld
njukdJYKmo8oeP/mgpsklth9RKYXox1vnO2efXHcqBzXy+FL7MDu2IUyMR4lPYEihbaNzzn8CRXw
w/vAdBG6rdYXAynS+gCb9J8XGMn0TpmyHg0Y77H3mAmFf7/A4hhV0Rr2W7x6rbILdcQJ9cnAwLkp
7Jlr6ZepQI2MkdBgNn/EW4XakcQor8mUlh6vZJglhB/rW+ysuQbpjA6u0bEyrLLm/GJQrR70Asle
A/+4KGML+frt3QJjOA7+RvYvsF38mjljaLJPMdjV8ByFBQvEtRC7OyFNKfSryZKOh8pnMIZttozW
WZMZo+8B8gnXtCfqKSSqvhCbiTgDh9wQO0TWCYU8PGagcfO/23sV5tfZVrioHD0+o7QYNoYd+MPg
7fOC8acCrEqxxpB6kQaiMRNgVMRwa9NhJgvNHtFf26CnOr+FpFMpxhvBO1+hOqza5cNdna1fFQf3
9HLVSjWsdR2tBCi3l5Q7eTkuzvPJKh+RS2futjofPqs4pup/N1Qp1+NfIgAA7lv4m7qlLQ74H3NB
l+w5sEnajsPwR8G7xDhf9ygfd+g0cmdWrMkEmkpC22HfoRTfdC6VyUyIm9L4x4uM5PGqCfJ/p5HI
hZbAdcKps1kLzwGyO42DvzEqemwYh5SMGKuoYacNrnWak5+wEC7qS2KpwmzLdIvGlLZ66BC0Abgl
XEdiZF1Yx8hwm8WQ2sh6S9sb4t9RXHGGyrfG1JLcKtLX2RgMox+27t5yuBBcBzm0djlFRCdxw4BC
ODa6iLPiL7VuwlKKXMows831mrN/J8qbZj0R0gJBzLCbgYm9bH6udULV6ncc5nAu/GVUtxcpEJ8s
tFgFKhbAl3SuMMuZKu3+Gi27fW8Wcl8+QiWuK//XrCRPYm58rRR+D9hWKRI/+z2XFzZ1U8ibhyAE
bYmn90y0SyZyRxkjwogcf672eT+LOS24jaAeFU3b5HLBRIiIkh6HNfGny2AZx/v0M1BkU0DO25zv
rCvsq6E/4nHRBmupBHesZnvOSZIa2vnMNvpDMHOQW9t2DQkMgVnL57VQ4iaU3p8lOE+CnHt28NXy
q1Q0NzeFADCLmFp6QE1OoMvvT8spBCXmyQs0EuAp37f6WcHOerMesDNfc+MXXBanJUxdtCXXktA/
N48j1b+d+wK5YPY6krAJkxsiEvWPygRmloMmw3fDb1WOJg+BKj2F/NNRISoSiCMmUjc/JKBv8Si3
uad7xXxc/hdFFt284R73BAQeCrSIvXXYSArDnzjs22VXxoWSwOiC7BvbtLyqLcJilPD1pMQxmk4F
lZWAKSYNzzO2YXD7B8PhuCwJx5ybacvjqUNCIDUxcXVQ+emW7pB14eE+2kPceUWin1eVf82kvCC5
BINHYbX9B3kTWBgx5+Hy83/YtdIbFNl+EdpvCHWMyspj+8MyIJLgmgDGtDPeLYCa/Ef5j1o6GSxD
ICdTZxKl6aaU5xo4q/rFuNoN5RVglOe+Q3wqpRbFfu1vz/TqZ/NVEWFOT1AeYiZy8a5EUeCGN0Bb
y064OURpHgds8C8/7S4TrnDLCFl48ivOoq4Hp+RV7c/jpLHO97HR/AlrxCwFjjE/VgZA52meA4vA
RQ01yRD6gvZ2O77Iw8Fz1rdmuhTrpYhkGYlM3lpXhjgxuj/ITkDrkRWK6T/UyVb4djaRHu/Q8ooK
420MlmreVhLzVrUbqjM7Bf0Q6ESkQHg+nkN+dTO/Rn8vr50U8nbGAFGkzlmQ31LWRIGwhQdmKFPJ
Chv5ngJASaX6FqLIrt2yrJZrCJmYRFZ8/l7XJmNc8QQxDe/25ILcc/5rDCPcdnQqjtiVYVdcUNIi
uLkYIrhdWGgkJMRvBNe3umOGfUHvOA48dXTR4OWcATVFsAEoX3LIA1clABFWorK0OFuKIx4IuCXE
lDAp3s0VoFy0fe8UREVTSu6YQb8vxmdCDx4WSSYOwFHSdVW+A80LoGQxuG8ZqhuLGoa7wWs03cZt
mpgKFDoxXlrpEpzNJ9uj31j1RMomgNP5G2jNd+Yk+kz1zQXpv1v+62vCPNUOuMlhNLYmKlszzNFf
r3mkz+P4qquxND58l4RtLUCWjWHsHNe4llwiUTuR9yKR+hfNzKPsU5O9J0ZAODiRNyE8q47xJfTD
3JK4yIZDffyv1Txxp7K9LmSjX7WgO02j0aNt7W4T57p+EfH/R7oEIIKeTqFyErdLiAtuqvNVXwq9
U5bBpF066V9I634cURV0UFRg0b7sjoJ0zCAGh+7V1r/1SLKaLcloeaTgRGqm2FnEvpIYvaQsINek
PNyr43WS3ZQHo90tdJjOIyryYXNOppcVC7AxrY+vkx372Ewm3qcFuTMyWsYH3Wgp6aQb9XHFCMi5
VUiQltKguZvXZ8VaN+BwaDDFqLFvfSFMuMb1Oj9O8IpkZ4MICmo1XAVzEPLCPdoPgdUKFVLwT4SA
mtYMplVxsCruZe6VFMWnltWf0y/FGwr5msjz2aUEYPBem9p4wdZJiPOwTVcVbPLAdEojL0t94ABG
syvK3ZWfQgVOK2cK3NohJ8XAaSPiWNAxSjg7cET+NEuBv8rqraU9ig8Tm8s2paJ4dsi4CgJlgOMb
tzxedad+7lNhmLiiO1mD5oIWiYR/7Rdw1qeoJTfeAupFK80Sei+diA7J/uuJm+uohrZpchHMl0xy
SwpNAy2TrAE18gxp4fYm0tLXBDp09BVDQBgcdzKEzW/IDLcnileFN8/+UjeNTsg6ycoh8LQ/WuIB
dxxnZBrilLbqURoNuHjOBZHMNoZCVh+ihkdw1y70HctZy9wOGI+2WTkHM7djkRtrWHVkRTrP1aZE
NfJ8LW2Iw+KkZstzDm+6n5P7YsmMLtQP7ofepSEZ6YK7ai5VnfTFaENrmYHyu32tAV0bbNwcHhfq
a3dnkfCBZ3uswz6px3ztFsbslEAtvH7KJAZ0Jscn0kK6GKQIdhXhYJ67+HKPKHyBK+g9AOEiPZm/
BHZISsMNMcgueU9qi+aDsCv9daXfk+reDEKsihtagnHcwsKXB+C1ykaWl/F2jFpHF5xWw72xOjCW
e6AFZcswW410Hhv101AWXg2NU3PIJ8BBcPx+kjZwmgOw66PJLslmRPZAAJj9mVBcSZLL+iKIu/Pm
9xP49nfJzj30Yil4EvfQTWQT7Kn4uaaHQ0uc0Nte1Y1TYsGrs59jbM+vsyn4abHhmG8+t9A+IQcK
wEK86bmaqYo35XdA5IDof1S2+ULvxyKg5QN+CM/IxD9H64CjSvqWeZRhDYmeqZ3fW51xCvVOwHYW
Crd+geB/TMWHGN4tA9N4eN3quzzNEZR3lNl8Uyqk04BMqPKdwR5yMH2L1vjXqrvKiyXBKxGOXizz
LGJ/e/ZXYOP2G6RVStIK7EXuEAz57K6BvxgY5gL7HhUC6ci+TaWq6y6U2npkcd//4PynPQygj4V6
aReo9vJmNLS1siUJdAHJuqSR75ZcOMR3oSdp5ESTsaA6cdp0LkGUngBytnGmxYJicpzkDMsezW/A
89hRuCRMZ/URSel+w5IS8cu/BpNJ1tQxRvUU0r3LszjAR+sIjBRBF/4X1Z38glq98HhCzHyGW+lS
6q4V5coO7Jbdd8us5VCc6eOeFYKkyB41i4BNLr9hUCw8DXI/HLa8aHSIHlgY+yFNjCEY8nqjvQqT
QxCcBBdSPubhYDFPnPQnbFJfuxIdeqArXMET75b3ahAWZkudxEeWC+NMBcXePe/nGCbrF5y3ZyUD
4RDNJXuvBr9+TGdGtoTlbAR9XBmT4hNOTqLk92rnoB/PtvRb5gnFstvTeaIeF+s97I2VuUgLk7at
4GlqVHr2P+xnP3iqZ9Flz61Um0s04g27WQZtXdcuY3IZmEvCOoC9ZbZv3QFiI9gOuXY4Ir3xy2TF
NraDz1a4AbzzZDX9OXnkrBdA9wChlQJRhhZTixr/boWlnxbFkLtrhXkD76f275qs8kWg4DKULG2A
+V+m/fKX00c6XMXoqX8lN/R8q01JTjPilY6pFElfDIHEA2A2Y/NWCpjtL50XYCOZDp/n+HPU4jJg
r6GYVLEeduSBuMgq1N7sXOwQWgEyPvQOk+M40RjFKjXS3rSLonfg535VEWgjSITEQ0eAbI2DkskJ
GYZoJEOm21GYXJDaW+CrnQQAZj35g9741xDR/WjFM7CThxp4SnhdTQClqTQIC7FYBVKLTAl93aVO
4lQEyDkjTtpsn/IF51fP8cdxS2EARY/MoG853zyS6AYyBTWSsDwxhxrMVy3SqkDbW2gwE74ZDZLx
MGVaknYlpMKsKqQoJXeqF+QqJBHnatxXnI1jYt3wxoG5qsJkdPFSNV0R51o0gsNaglGS7dFmZVOb
dFQ45GRU/kiwxyyzjlTwx41ES9mxxrPa4bHlaILtObwSN40BMe5Ux4kA51lF3alvWooXTuUnA65W
FR4RdBo0lT+nxRXVzO4z1xXc76LZaAwSKH9P7wdrujRsmdub3WpblKRsy0w+FjOlMBlDV9XwAZhW
Sqb78uJhZoGxZOvTZO6BBfZMWSWypSidGLQRDnKqPpPGiWmPR1AwpzKNBE4PCPPBH6p93kpmSDki
eBxeu53iTwcOd6KPcSQQTkjxy90vVyA3qLY+Ne7gCWgeoA7D5LwjVc8pGpoEz7J+3aFM5aLoAzh5
omhVl6agur1WxBCXagE0fBlRhT8STnBIKjjUdYKoJFsa1pKZnWtPmPKvnEpxH7WAGHzCppCvtLW1
0oJFyaznyOOrIGK5uVtb3OaApgjpkKi4FThK1k6Mg5eeOJ2oYsQqnWxwRyslcOCPHbfi/3OULNe3
HbnOnN9GOUTga/0Ek8QltyKeZMzz/9ImmIDDNb8RSY0JWK+pstCY2v8diipk4Z4KIhjsW+jgLZ23
I/vumboEqLjEE77UneQw+7Ugttkx9ksK5rav8eLEqJhmF7U4FXG+dsd1Cg3QtsNgEtMHq9BuZfyo
YsiYW4OiiSVQKA68o8m094J4zyL8XbFf3a7jCb9m3h7OlCx2nftylIrK15ced49tT6DZZOLE2gk1
zmIl56iayIg3u1xwTlGP86/nG7FRnAaByeryopG/ntk38lNN7Mmvs8a4WPL+43sXt5pEkBLR2i7K
HvcVFW820qcqJo2blIG43ifuGaxZ5pwejYoXciU9nEBSnp6FJIYT8tNS0DpVo4GUZL3WQ4BhIB7+
m3S0CIrqpkpahvV90t6/ztN+VyE0/dJnvWwYzM+WOJ8hduSJuu8VLXzmvwcB8E6SDfxjwDR5pNgy
9iDv7zEGw17xI0Xew/ezsBZYk1s8fV4KFi3TAxCIjvV85pSvnXTfhNjeb6u42KjVIKbCu6mgYX7i
oVnLrQBiS4qU8Jzs7s1gk5dlznhHAPNr9II4hDwuZ5OFv0mKVb9QIOo+B9l+YUuxLZDVphuhjwCm
uzKO8ajBRvcI4+vwbC3Hb08IbNKFKHWUzzQceFc42ZUEOEGcIomksGnFww3k9/wxuLLtbXX/k2cv
up8b0PHw6Y8L9R6+goU6LaTBPhwChSlWcGSlAKzsUdRbasDmJmzTI1hZvg7pLl+ndGl1C9W773yx
2ELpNEdviG+x+ywvxzfZXis/RqaFL/S0RLW1Z8zy3sQkZm80BrBYuP/wrO6AixIrdEsSaTetjKWI
V3T+jHckkdS2UwcD9IiFJ33ps7uarsao0ozkv2l3ZFMQYmhtgY/+faCYuESIUm3Q1Hd0gI/T+Teh
3F3co/m09JBwpLgZL7iH/RjDNCWRXmNFZEh3DyT68tBfx3TSfiXDVAVEgdfUxdUXOrkuMguH7IjJ
e2s2mljt3Hr7aqSUE4rTw0lTE1I+b8GzNyOS2BjMi5G9aXfnmXpRl+Xn/GCLljnpEWKjDx2pVx5p
nTsLe0CgS+ULNlTN7mI+GXto+UZR1bKKsjcUoA5enbzdYfsQ2ZBwWdQbYhrHEhjGgs47aZfeyZz3
jG6vcf08+6J65ZuXVNKpv1CfwBI9RtYOogDLlCi+T1/aj7i/fNQjLpD6s9GiQCTQrNJpyXYzBn5J
kywYxz4njczA2VJy27CMU5+n5iRPJdkIHKrT1nLztDBly0IqUDT5mMdJSmqnKEBpyjiip/+Rtowr
b/R/8s+MJngH3OlEpNvMEqcubY5lTrP3rGEzPU/ZxmLuev4k11wrbRX0lIWI2QEUyuE/Qk4HhSX6
qsXfG7Omqv0C0RuQZCpsp8hzJ8YVFqo29vnQ7AF0TAHo5zb7DkthOTLsX75m6fP0+KALHtP9W7Q/
MCccmft8M5Ipra36CiSXnYvZZyWTDB0i3vVXt0RgDLpjz2sTUf+VnrUz3Jb2btavi0E0+7gJ2xO6
nWsxLYcsCzwnxVodlreKC6ynIWR0OtQ77/HeBXjQLVri0XUEQrizBEvk36qIwt7nQ3d9g2N9Gh5e
jcNio8DLmEAsGcl53YLrQfnWX373JReKa87C/1sLQX6+Zn0n5cmF0s3vL3P3MNt58RWttb/y/VQ/
SFXz4qThu7cKDT+x8uSu8oH2xwZ2+CAu7+v6hy5r0bz3RTWSlScGDYwDdJT57p//vHI98fnodI5N
l7Hft7U8i6cHtXTD+pvFkl8TIkbAKkQOiamHLAedr3YyK3ZIE5y68HrFjlZo4Uw88VST+VAWTrrW
mPwd7ks+sjDlxgMkbk6Az9tGVqXcWHrPvB1wlj6Ni8mWVyDXdd/ZYKQoPr/tkSsn/j1U8muIzDZA
D1iDOhqs7pZcn/W6ojXYbdBID3DUsQqRm6Zso4zqLKtYTYb7LiSqbje/40PKl3CNMivf+NsLVkZP
byYV4DWfqtJsOgMErzEQcS4SOvbsO+crXTBou4myGS51g45z4ANixe9T9pJQwpAvS7ptIntAnyp9
7d1eCzeLjvp7HUqtDeooTfgOqLzhch+skjkV+dqv3F9Fa2XHXaGs9YXJT0/5kLm8DudiBuQEO8QK
55XG0N1fFuLDQP6z6sHnO8GsSpRMe/IW7359oEVeg3L9sVFFvpdM4kgPxOhc/bgONRu70PS05JDy
aQCANUsEjzTGebZcv1bdGq04Z7c+CAQzQOJalfB3WZuZ7sxG0/IRR73yB4UlbtBmCZCZTFxCG0TW
FrLTAEwCljdX6zgLX+bqOV5fs/8IGcoy69m7q3/dPbOJz7pCSPmqj0lnvMu/C9ft3US4r20R3lNu
3FXk0waKzEtYmLG+ts+9b0DajmF9dTICr9YsqFmufnfy7rgu5uIfKtLjnwDUGfiIon78NJSPaZP9
gfZdav5+5V8nCsIg5HjG53o6aYyuSzNCXYFkkel6T06MplSlkwRnosqDMQ3JkQ5+gjDWIUd6P+tK
g6uikhyvi9LPPnmqwgtNlpInZgWp+OQFgVwPjhgn+0k+KuobhcMP/8HzyUkkiyWfpX79xV/U+Jij
SShn6jlc6vanutnUQ85bWkxFB1cGCxQDPqD3yYtKwIv6vRRXK6qgKUUDVQgi0HlFsZ9PoH7VMVa1
zZxDPJfzfiSeq4LqlyP2DOt+MTlnb4Z3R4jmYAQyLTC40yhGHEJY8xpH84tkV+sBk5iA2vzXQESS
4T66N+hte5pbtwDMg8WmjJDSQ/T33Hyf5Y80d3Oq0qDtqKCa887fphEw3K1X+J+LNyztyYmkiTai
C2TnC6UwIUxKN2KJMjVKBg3f/jtCWYgqEsXrRXoMz+suRGbRJLqmidJmsVDDRMfypuUV8MetOfOD
QcQyp8H8ySObYNf1O7NVikMZwo1zfS0HGM4TvfuJvRqpAuT/D5mUNu4IzcjQeZEorfygUU8tZK9D
EH9d/PaQqTGFIbN6BbFXKKS81/KPBtGxJZj3lU0keOkE9XKQJJniQ0Dd/w5iVh53U+OCkRZ0LkVJ
kRXgt1qWWEJk3Ska1RqQNcL9paUDcraduCBhyB42jUHj6JQ7tpPYO0x0XlJhcWFgXyG4z4eXltMz
4lGHqEWFjfliy4/qyPMR+VgcsTyhr9nkIcqNLlsWC0guOGWTmfDQ67zuQ0HZttAWFhmy8GT/cCZS
kqCBGQA+MuFJQtEE8ALUxrNW0XPJXfFnBeKabNtzMsvTHw/hNEIDzyIz3e5l1Rh16e++e+pA7HT+
PA15hnXLe+NiNf/KVG5cGqMMnwkHJ238wDb8yESAprDOOXi82u0/M4GH5xIcOI0g1v6r4IYgFaSf
XP5/TLHYFCFj1C/gF+mpPO94yqqY47CzETiXk6+0nu35f/6u7BzNDVBQh44rsGrzCxVNhyqYAhg4
a1AWzGHGSNLPX/oT8ffQub1rnwHJVAjbuLyXxkz7wib36zl+Lo7kwHexP5dagiRzl8x6EtVJm8FY
aDPHCbt4qQlA42fXGawAYkeaKqE96H95T3AhrWh3jJtTO/6GHhDBQvRRNLPOkKKBT7p0de0bhBak
XqXKBAcO+vvJKkTl0NpjT1iAunNg7D6P5uCNqpZnsFyZjm7INEboNb4I0cqt3rIx385qF/vUn3Uo
bA6HDCfPzm0PVVpKo8UcIDW7kE9ZafvH5Sw5pDmV4SPyQjB5TcER8Km2FA9OsguooXEWuW2KNZny
k+d4A0CjHSrLzkJZXssQfZ7eHfo32o5zfrNaKGooq7crlis9QNO1CNR5OznQItWdnt8YyZASJEjU
dTzji+dV0CxlDrfs0kuuYuvptBK6uFmHip00Viak3xG2PLA3RNeCMTW67Xv5iTgnqn7c6wsyAq34
Y3jblFkpbHF+URei4PhN9NXF0DUc8GGCimuL/Ct/eyGFSJwB4babcRt+OjCRJBjukJtLFLy3+KGb
OMjC9HTuyTH4/dTh8rSI/eAMGAFFpcKv184kCjo8u81jjJfL8vyiHT/tguCUfi4vVGcM2DVnGOOL
l73zBvoTk904fsPlNNgtMxJNaxU73OLP96Gtzb7W0Kzwddpb78E6CkX5AbRBw/w9o12cfd25i9fn
eQQEgaIMux0td83lYoROatB12qstrOXziUfGpRTiIs1BkORDdgzwj7SIisv8LHC/sMcfK8ooU9Bi
AiXrVE1I1C4qLIv/C/6pWJWm8tlUzOABSkbue+VzRH92yqUONRdF8dqcEPXA9d7VHwG2M2QW+Kc6
B7iHkSyOcHfSGs8ZjsFj0OkeIU/Sl5CgE+VU7ALb8tbqUX7xj+zzelIwQmtZGHipjfeacmJuZ/lV
EzJW0UxW2MVjU4C+uRCSPVslLQxHi0Ed36Tada8IoQGVXqG8sdkbc4QfvVRrsBVRXjMpaIv1YrTl
IPQgYtr4oHB7UNKkBa+Twln4TbeAf0PBuFAWaKxURA3Bz92PuTyFkI37dxILZPpWANpP+AGa9AXa
KEG3BzeQM0T+Bz8i3wCwn2RUcFkjVxMYuUYimLnoP/4yZHat48QcuRUoeuhRY/JQAEeSazwvfeYn
gxfsEO5uxXJIXnBDvhkIxJ7HXqG/C7cFRQb48OrPpA3NkIxoD/4U+k/TWxv/nUxEAxMN3VLa1uyH
fA3l+19imrRM7khV7LaSud3pTl6kxxL8Glx0i7iZp8wzxURviydLQw4CX0qHu1bTn8zHL9D67D69
6+6hHonNTj447BTHjbqus5PQXPg3lt8hpEwgmeODg1eszAgvxPCt+TDhciY1GL456A3iAaeUaqit
HazTYOADlQRNrMdTf1g3vqIM+rHWY11v5a7m9J3hHKmwgOmxdNsfmXZlHnh4SMEk3YoW3+qjACbL
JLN0qv6dK9WV1xeyuDuZ0VyULXXqAoH/zUq4cXOKKtkdWd6Px43V71tU13mjNP5N4/C/LIRnnnh+
xnNzCuiyiWu8ltLCb47gM9IbthdrPZxM67Bh1Z9jUg5xf6OJCSqlgxgb02lNngqngo5QwEX6u4OL
ZgVfuvhpUuDG1PHyXbPa4NUkBqRr8n4kzo8h8u5wNO8wKUHdUELVLWShnf7EAmYgF/Kjtd+lilWj
8Ii5NObIBBHiSunRB2byiVRA6XM6+LvhR8Es6CzQey/nLYBciTnRbcxIkSWmspjfNIF228+UJoiU
Ai+D+TFf7mzmMLpViqx1EvRDkZ0Ka9l2JL2OFKQ7NoNCaaFgcJfbvLaVh8w5YiscCBpxspiSBMIb
87wNuhIPGV4JxKeZcUZVwILFVfruHU7paT4N6vktlXzTWin+ui1Hv8+WwhYgOfHRMsiZ5h7zrrbK
TgGZMPVHQ3RA5NWZbYBDlaCs6wC2KE5pTP+IZyQHvgEGel42ZE6b72HVg6EiZwOsa5uw4uyZ1+a0
898fctKMfdns5ffs6s3VZQ8JnDyJ1POK8pUJ8uNho7XrhJv+CaTK+xSrnZebKucVYYnIZ5DBl/7N
qMi68RM9yqea/mEQNeJbLCYJ8PSQtpL5AyLv7Iwq1hpao9jAutpeCwi0gn8rKfkPoEyKGPJrGkdQ
5Mq+Fwj0xiODsT0UlkZJCBDOTUpvYgg9vw6uYS1pIue5U2BdBw+oztfgagxJe46VUeo9+NWsZCim
HTIGjdI18Rr7Hz85yTRiPYRiCQakAxIbCFK+R3ZDZEMnnoV8TcyjnXkwMJgUNt3L9Ts+f/Mfeyf+
i1EKVTkOLx05q3iBL7kVsvcwoFwGa0VHG5mDQAJkqozF2InQE0eU5+fFillazwnIUR0bD+m+hlWj
CDnnrjeUYXc/tEJXiOZZOWQW9IlJZo8pA00yKEgNvsI+gOgu8oiUcGrjdsaB2fueqVOzQQ9EYgDw
UMOnhunR/h8iHpo8jhmDQ6XhkfuxW1WFHBxSup/H6NO5ODl9/b6FVeN+h+RtTEXJYiY4X3lckso7
2hdr/sCLKMHUdRnahM6JEAllC375oh3++e/MdpTMFilVUrrcUst90VQwtgDIhwUZj7jxWPjm50Gv
JM5NQySAxpPoNxp+CjrxnjIo2Z9bsjZiHUpxXYjYPCyXKg3As5hdp4qCfe495B3cKYcNHMXUGqXn
nC05kdGU3qkbF7P2JoSQIks5eDvX7+M6DDkXMYwt5DfwwvIgKevgdhq01AxtiaVqLSsDAQACC9Fp
4ygOUmldBHlX7OMd7D1cMki3Kd20ij5Gluiw8ONPVterE8tqegZJA7tAcnD8NiNBUaqbzHfODOiq
1lXEPbu7mj3eX1NPxL8JSY1If0fFUzODd2DiF6Q6QB6G5PK+6ZSjPveU5Q/eq8y0FRHqdgeoVLoi
O3SBSJD2dA/Ls/QESBezn4FJMN1fYJ+nxYH7YEzs7UvEycpGF+3Ts8ptVxBZEgjJFjjfQrC7vgBA
8KAJ7QOX3BtRwFlp3GVCptkO8y9Ke8UCtwQBcZLQd4g4/R8NYbWeglvBAfkQRrdcClM548eQOE/n
wZQkif8eOeABWwHgSzDCCYJtGkyPNo8Nfuy/+bYX5A6kOxfKIxGO5qALjtjaqK4w88n05A9xTutW
KTAkR9At6w7W/D8eWAgi8z1/YgK3ufRQVKoKmqKip5sovM69jQDR0ZJsgWJ3o2lLucFL9jvTx2Qh
V87xeYDFwXEVr1WEgHGKsPu1xeC9AxckHR7pp09B3fIQQqoyRs0Xluc3GVM8GjGH9wUUt10BIJVc
iEbsN2/a1In3M1ACeedTZ/w2iLILSuMY122+yAWyXz+y8NGcL2EhaIjxchbdH6FZE1dVSmXjUygw
gEv2ypu02zBgAbghvHvGrXP3frPxRrYekssCyZjH6v5z7nPpx4RKnxU+8XxucSjNrsU9C6VjNGz/
tS8c6TKW4ltyzXxP4FDhhWh7jyz/2azHkZgfbpYRJajzLt/Lduz2cMBrkFC38RSlgTDCWL7wCC41
ZWRVLYowuaiY5ZJ2o5kMz4lAij6aCwOnGa54l6i3jrIwnD4h16y24jjcV5OEjU0mAgper9AsqJw0
4yrtVERsFL+hp0rJndNrQp2vz1s1Lt51EPy/bhd4FrM0ks+ev1Ck7vu6beytHyDW0soe48Iqh2pL
x9u1hqaozm+1Vmf3Z4HyPcJGN4POm3YVh10ODk+K7W3uwj24VbVev/DkFq5rpME0CIlPobPg0vdY
QDiIkDMqKQQJtyTxwm34EoCNz3hBV6T6DzDwUfBn2w8Ch2VxJARsCCeoh/N6iMY6fR4g6M2LyUqT
w9HtWZyOtKP2mfIHy3Yc2u3MYQtLmRi4xorwj7v4Y9dLfvDFqVHKai9l1wD/gQBqgOzNpTOrKClE
mHbFLGWHrkvVLhgqsdHyJb15IbVzazjdxOTq+Tmiob9qR2oFfalOHF7RcNE6ifIZwPNnrdrUDLqE
c/0ui5iKCDbOXpLj5sPHlQzY28+pyo2OWfE4jwDVhA8mWadlhR01sWoqoKQ6YIz8qjJRLt3muxaO
rvP3m+G7vnX3MYHF6QE1kTkzDsr+Vf78NNQc6dtjojMk/BOnZapDdA5TpBLGU8Kplj1uy4/LxCdo
YdejN5Q24Vc/5XasqnrxKUsD3+p/8pnSHySHMesiEormJS/EFWOQ8h+/0TM+7Qw+s/5TPEdhe6ve
bU37XrDIMWFSlJogW0uwi+PLUtBBABDPPA84PfDhq1fyI471xOVcBaak104H3gAvGAgg4FudhhC9
ztZ0V0OMdmkcRkf6tY23B/86+aj17UdF3jbka3nf8IX92q3I1akX60UpJ+7FAq3A25mtnF73ObrE
7aXiAQzDlfySBirUsd5aS5hwBz8iPd/ad25EsCLikFSl+0pqZ11JRTC874LsN27GoWBVcwVB81mO
eqAL9TLMx/87RaNRyqJY8lat6Uv0t2ocBOkrioZsWA9GGxl3NKpjlVKELHQaR/BeEXuhNssTCwMC
TZqhUB4WO7nRHR24WGRPn3DG/tKxOuQLfsZWXGO1ixs75elILmaiuiAtGj/r6jDe1ATcVmbTM83K
v1d3P58o0y38k+/wwC2zVviib9BuNOiNNsXO9Tt/Ol5zdtBTmddn4xJLhR46rl/ty7kwdBcWNRUI
b0fRK5K5tqoeXEBohprx//FDzwscin2EJIpB2j5YPmOsKXA/3cHcwb3d+RIuItd5iDRvmFGAeVXO
7o3goFG/NWTplid/LQm1s8GEeyCsdT1gOjFsLliezVbB9sI4OoUNBFXWT8kv34iX2AtShtucmF8x
o0D2cJaUuS3BoQrWrF9XqForR8dTPcfWCNlnUIcmBB49te1kK6Qvd5uXYUL0DNJJvNPg8iz9OxoP
cGYiJkLTXvKnTiuOIVwootDhi1Wf9wJSYKQjp6UePPyKxkq9pv0eOChopctuGTr8vs35Le9qRGVQ
6+yMVwXcylbVng7xCArKQlYUTw1N/4/Oh55+02qnvZ0Vot5nB3vF+bs5WtPgVe4WL9jfmXeIUOgB
/pYd8HT7tPfSUQWYQUb4BgQGM/lMxi9InPwKv8srkpu052ufMaEMOdlp8rezTiOMbpnVr/52BP5r
DeR/etOCbCzwyg0e6jOXfv3iAC3bK6T6iYw4Yf3drXptqMvc+xD8xQ7DFx8STCqHInRgADZSO/HF
yQoy5Xc190p3M866JfYX5Xgg2wD7Zb/C3OFIpRRg0XQw9jVvS5IEfKuFF12GPpjp4rgN8aeULtAi
BZ4GkAweM+X6JdWx7sz7TTafg/HR3uO5EMAmh7DeE6+fXoz3EGLF/7BcxxrQaMlCBJCcW7xNFw6Z
xz3me0NOyaAoZUOFZezKeei77CPO8BVKpaVQwdpHKhKiFTn/55NIF4eaj1jSvow5skylcOEEyikb
6GnwyndEchj/Bomy8uPxKg/5jxV7vR5vjEWNGB115tB/b2V06qhtKHilynbLDYNwNP7ACeU3eBx2
nTkw2O+SAwLfns9bAHdpqo41H8ymoYGWDPA3wPAnEu3axaNySmqnvTa0jM345nSuP5BsoTvkLDdA
2op5p1CLWdfUThqxcdMnWMiI4LehqFQ3RG7lqLdzs32EXFpclAVaA3xHvXvojVKiBsR0dMSVPq1x
DGoJWKtN7uWNTYgcl7FujovvRsnVq0lvYoP+w7WVg0wUv2pvQ68qPP288TEZgPRU0VzTML3Bfx7o
LenycPtymYFafMCGKtB+zeLp/4JWY2pxEQ8pzVrSj9JVUPaLj187JM7LmOl41OAp2S22CsH3waaC
lY4opEDqtiIc3BokwTIwxx6mOLBIIVmH5XnC7aH17Pdtq1j3kFldmWc4p1ShXL/ZFDdRTKF+KypH
DOzddQ0WthZyi0i15xLDZAM/SCx4zs2oZxpPnOEAGkWChgZz+mKlQ1dPxcKnFhIN/eZ8a3nR2rfm
CATOrrICIclmCXk+1sY/6tv6P+22YUIGmnqT8lVn0T6a34uqa2hQXyApsrkw+ETl24CWulzkdP1z
IbrNcPXILeX8pD919gRFod0CeN8jh8NckSJIajW0RH58gwD6Y/zY+eRPklcNMw37iy1O69t3RwNO
9ZkHA6/8M/3gOIh/EZjnVTNMikL5kEXWkL5EUiAr48yQhUa2O7rIh1LNS6Ejwzvjzhy7wfHTrH27
Nr+aMFoXpvVSDmMPXRp+f9oBd9i3A9PHhu3gAHlSmBEUJQFDSrQP9KauqMcJ22Q4wUabbujcfyiJ
n4ao3MrTz57sVcYp75wit1yhpsh8+c6qRv+a5mrIFP6FD38ijLlw0rabImvEmxHqUyqd5joCMvad
UTbdpKEpitOFBtjzERrpXD+xZZYD13jmG2cEnskWrGvBRaMTprXz4E8PQ9dDRDT1oSfE4ghb98sv
FoRhyah3N3kXVbFG4JmEVlDS3ZGvFTbQe1edSIrMXMJ0pmopRBGEgFZovXiBcFaK0Fd50EyJe0sK
pi0h8xsrF3hmqrFAXZ7p2Np34ildqfw6RXUe9GhqWN130gPHib74o4md5sdjIigwJCNLQLWa7mmM
0AlTh0Nbxq4V+RWYysnJAbq+b+pDPMDFnt6GrPuuHs2nz+4nQ+Ojlx9xryBwJzkZz4yUFkH4Wc59
55ehs5NXloNOnEG/Wj4S0ujp39FJ+tsH1KQul8vXy4pyUmjc1a6SfvH2uYaD55G2vqj1n9pLquw/
bOJi8p7Awpxz6p3dE2u97Q16sq8j+sLdCCnN31cIMZoLLvPDUo4ke7jtnSLvLOf66UJ0OeAh2kVL
sva/vNdlgkW7tSL07k4iFBPwsv2z6y2qLn3L81ZleUfNIsXsTBBLYm9aCSuV20KBCdsjBdtaJnRN
RFr0JC4AFquJgTrIabKpOoTvww55lMPUUTBJbVYmzRLx1ZsUuPiqJur/amW+S/D8RB5hOqjbIeoh
1kX2996LGTa38MQbqP2NHz1x/pgS0gDQaVmHb8K7RxAZcOiKwnslnPY6azIVOVekyrGQ9OGbnjyb
saV0GCL8QkBZSttGPHBjBTbGylmnpyqD4DWWnqH/q18zOp7YdBS5Qq6mvmk3xNGAV60OXQ+/P2oX
X559ioJVBrsNukQZxxwPALf9oMQk/yO4ZWrbJeJIU1oMBFmee1luHL1jr2t1lo5fixS/kdAZLSHR
QV5fGCe44BvkRwjFjvoH3YUw/2hw+fw50TQ8XYaPLqT8LQL4pLZNGBTmKsVTS5bDebu0v26XHLZd
Fjn9fCVH8vI3fKhqPC2bo7wKDa1yOYoYdPWRPuP6h8IRvZE7/ryVfsWOxJuUb/5Sc+Xj+DZ6y8s7
mEO7UbenzqbCAeLJ2FYI2rjmp99xy1Qgux2/T7lRsLMI0jw3fKAkKRCD62IrNRxFyesZW1SZvgdn
9wQ0789BTfnmD9Lqf6apem6qlCE6+Fhg5O4NkjQlDZ1oEkHHggTiumgiCMAkS7RJMK+yeaiJfRNa
miA+bUYL+rDUT/BVh97mR5VwPFyedbYYF7ggeDe/8a9gVQ4PnbztQj+dt/rsqCo+mEJqYsm4zUIR
ld764f6xFHj/eYihxbUugKXH25HULiAVbsVouUCI4sstBMQuu8McIsge6hgQQ1no/ACmbwzRj5HS
JjaSIkV/EaWHz+4IVbfAABdHKJ5pHkqzDXmP1EwhyNM5y/sCob0bUEkvi5gMbyRNQnUTqzfSxhAt
Ypdlx3zXH5oyU+bV0DapPnq+9uEPFAz7RuT/kMErESJ5fvkhAENi9xOBm9Czt6SzYYol08fsoAcJ
XRye0CjNrulAh+lOBEqV6Nh3UUCUh8TCUg1CWLplK7tToTzXUsUDRPLyAk3z5M9FKTgpsmc8JUAG
P8wDc25sZggzrHmA18rJkXF84GFyZxe28AisHsIjgq9zHSeOQzkw8RO8WnnuRQkyjSZRDOd3h5uO
gHdgeck2xLf0ceYjEi+f6sbmJ815IUCTr3ncex2NHYDdcpmhd3/CKBc9ONYsQ6ORM2HaXIdNMuKo
zHi/3ojNVXe+Gmp78OGxy1O4uYawOBQ6Ngl7Ua4QpyGs6taK0R/FQuoYyR4ZZk0kfKXZOqyynk2y
VWOoaVYibWDNk8OJReVgL2n0mt8CKbD2Ulwv7W8mPJdoekvpIJ+4llaL/VWsSwyAYoDIpjPd3PAN
MiryWwYy/nT6/IH3TPgHAqf4i3GgfrgBDi/+dGzUbOS5/+xKcwJhGo0arMrDTsoHidMsNCpB1r9W
saus98ne7ARIreXqGHhHKcTW4aYybPDWEoCeL3P1GL7IPmvr7kpbwolkyb2vzQ+RQZJEj0bELLlv
h0knhrCWTIMW+2X3ddN+lma8iV3jscw/eb/UcQtCaNbdLT2VWiI/DUEe3YSpKmqZIKiCSk1+yurO
5kltlQrU3GyFjBlja5w7ZQYOQemJEiESdblVrSK681dllMjTLpISwkO3x7EY3tpcnURw9mpwQD+U
hRMsa3u2IMNuTcR5G6R90YMj/zetrNGQfrfeIQgjgw2Cg2QYvz3mkSl5qkYruhcBVdLBXkyvWLSM
gMCw35iu6/k6Kct6R7sgMOb7rhBOnaFCV/JfRN6f+Bki/crUgMMkSdt75EXNVkA/vY5ew7FdKK4S
1FMjFd+hCeBocduw3HP6qCCd3Q3Sxv2EWl/AjBExd45Hv4tb5cXCI2SSNTS6rtBSJoxyBcq+Rp8Q
JI2hvsgfB7MNaquQ3QM8pywrxXEer16YE1ykljJP3VQxWz7w3eVLWKxZe77gvDlq8musgmSehaIJ
MC8s+bbXiMWhHxiQxKfpaT0rW4jG7KgeUrdiVB3CmR6LehdKLtoGmm+p9HpTpCLKaPzhN8SJWS37
Wd/7EQ7C2depGiVrrpsdHCFzRBcr6Sb1cDrVov7iYvdJatKEzw3p7Va3n0fi2cgm6q1nCVMWhEWn
uuykGVYBeVP1HZzZa63Cs2j4ZWC37MyC5FU0yyWi/eMo01tWIxgU7FZmjOllf9EmKjVDTo1iTxQl
BwSmz64CKl0mMkOyAvWA5S3QBrI5o9c5xeIPUtgHCHdEZzHINjr7Ou1xB/rmgX6wSl4tl6g5ERLt
Ida/udd4xyIRw/+Q+kYH9OlKy3rmgC7JtsUuon44eRikQSJ0a4nuEr33q05SHmkWBveHF0hRNuH/
yMCI0a1BN+6YNgv5ZBFNxlrUcLPydmCjC2v00S8Q0Ppir/EdD8/+kA5BnDlFyRt4rhtSA2W5kieP
kH5TFtoqQRALwL9OSea6TPFG22vneReSimUy9BiPuFw8aw+CHnnUT+2CtClZWATQvVcXikHWxxKj
95nJKiiSr+FRkoN9gT6rHdeJcQc6HBfJDZ7MI9NEDEP5b72E7qdCaxYTkj//Ssdgv6gsa+cokkAq
koi7tDGQI/Hwy/I2D2pK4NEZEA8aSm/F+WNhGOCiZpACg1gNUID3+JKy2a1DsDLtrjTsqCiB6O6s
rDa8/xrxpWk2K5BUKSuO0/75nsOeq+9aBbW2riNDmFunc+ANzypTBbcjIiWT2weWysLd4KJLstnD
PaJMGSsiNt1rdr19mtg7bsdwUstBM32MZyPXhk7pikQoC3KDCNqDZgFDUuwmhF4i6GLIGoOTflFt
E2GIA+Pzipi0ycDlfO6SeQr7QgUz+L8ENbH+uLrCAkIsO87lc3PVpdvhU0vsZV3XvpUzRr7NVCGi
K57BTTQGW6OOh/mzqR2A7UsoTzYVEGTH4gJQNKGFJPwymGvtBQav7bWCr6sioc47WyzljiQQPskl
6d30SE1sstH9isGXlwDIGcQoO+TFFbv4sJ6JriuLieWBusZuS121yDvs5P72ESN66Hm8voNw7j1G
ndlHNJPJjIUtlvOfL1b8n2HoMNOsC2oGgjo86n8kjxm7QrJzYPXRvzwNDqb6vAGhVSYYtahp8pud
N+ol52VcVscPtcNK4LeKPMX9h/qlDwUkz9i5ILnX6cDt3oTtgojofbvfGGPZ1WjnMAnrXYo/NIG5
eZvdLIImYqlIcVYearERh0EjdXe1PjNv/ScIG5ZTaJZA2Tu+ETkJyETPw09RoIW2oJAVr/2RDZL+
Ku75sHo4P5mvntdMtiOe7q8giVx3kcsUBxKIOpChzuPxHYhk51BD9ceb3g2mvRU3xYZVyBQ9xEoZ
MTu0WfPJ9Vv4fQ+2ofB2MnKODtwb9wlgtyCAlx6Q7WYTKw+HqZigbULoidFStv7nH41yFzFPJRm1
MNjCUWs2xj6iXCNVRAzO+KDhoYmXNiPLxliMSmHAI0VhXmGW3SXGI1TcnpwpF9TyQgmVETw5F4Qd
RvIH9FzIg0y61sWlKfeEZbi3g0DFPDP44ELnkXlubEpVDQX1QH6mTML6QKH5913rF1+vXK+pTvv/
5XRUur6rhAxxXwzLMPE64GllU4cQ0m5HLNJCAmjLAZU50SaXUZcvrYPViap462y0EWgOp9c9o+dD
1nx3NvluHMoyFUwUgKq6JIFa+UDWwsIb5idRTv/gm12xLFUWqXDSzD/jM6OoBPLDPqi1DQ4aTE2H
uU41CvANgORQuWrV92p2gCQNBFfVv8ZiKqQjy3ygKMNYm7xfeBgir+9KB+Dcm1rK+nmyVS02f84g
uYtTvsLoNxygmapG9V13jhawjeQhyQiDoJeZXaoSFS1jkx3Fqd4yq3lylJU2Yb1S1ubqwvkMZWhG
uUeiozSsTgK4JJoIgzGUbuXegSg0hwc/DubIpEAonN3c1KRlgKeSWFF17eD3LXN0OR22vY1J2w7e
ve9SvksOZw5v9TvNjW1Zdq7uNBRCmNWTdtZdtuPBCP7zACH11xIPh+b7b8Cri4vubGJ44K1CikRy
xPJpzd6ycskfU67eFAwdQ8DJP7qZcRfyr2SYMwr97/7slrXmuhhiJAKxCj7nN1RWU7gi1lHbSaeW
AMhK/u2nGhVy98fwDmDtOTJxQoiCPSuFuzvRrf6qBcVLYhpLMsx+iUATOmBScpQoSYR50YT3k0uT
OLEARgkL+87as35tINeJ8+kL81Guprg7SrlhWjmUZxPKUIBhnuE3By6qhwTTwSDzZzwZQByt+xGZ
axmv1javcYtsieeV2g0+N0xjikqO+3X+z2qZ3UjFwK53ABQycUWV+KJix1OrWZeQWtr2d9AzY1ml
kWt280I0QDmm8MbngRMZuBIF44u2QX9j+YaYSFkehIh4OZ85G51G625i0TSKsbbkSnTahtyJpZpd
8erSU7zzTqTjYeku0urp39dZkfBjeKM3SKKKFjbs0TEIYT4DF40Sajl4/Rz0QWD8SpGkm6nz703Y
nrkT/VZvYwmb8Cgo+AoE+JEHuq3jtnKpMJP10LSwaEiopnm5wg3xr5teOnNzE9SmZ0A5WVHm9nb1
upX+dTQI5YbCW2zb9d5+6Jb1KFnpznhEwT0b3+/etBpztt6eqUZdlzG8kpaTljujz9DzHsC22qae
rjTDtRuMpYr0ac/egydosDkCEBjuP1m3vgnmE/ISMfTyySnMOhirrulYE5HNKS0TEmUawdS70hWS
QUwElQIk3BG0F1tKhMgzyI4rOVSPAgAmXgFbfFKtwgdLw5je/EFJQMgtp/PIoCmG4nxfwxRdrZcu
jYwjry6q6tqHYb+cs7Ad4AWNtqUueO7fZNwzB/pQ2nAvCKpMDyUJyPI7cj9kX2vapNKgBU7yerBL
Vpe6Gd97mDP5yhYgRxA5/bofuixV5IEK0ko04aRe0ktPpZ8ZWwH2RXlKEpXJYN7Q7tqRaGO/QyJ4
Z9HOoUCk19LCgJ8IqjjF8V0y6Nn60ZkmVy30zUJIJ5knM5wKLkan3eyS0Go2FzLi7e4GFfbLJk0v
wPbb0H0XgPZVClmxs5drAy8MjSa5lB2I7m3z0W9VUahbMjaQbO6mu615ULOKm5MGoUXJmqCR0lC9
GRzqxHS9rs6P56FvkbksdP4sZHuGfyg1L5BJF3ccoELCHJYJki0DmR6NKPph6aYDGzQt5aaD4hwl
AGyQNqKqGNYRUPrHARKPf8auHJxoZVmjj4irm2IsZW4nUnwQogi+CE456X5KlleFFghJ8ogWlo9f
amLxUd0LCoXeelGm9ytJF2Vjs5s7Z4j6xxjPB7/ppRYpSUUVQWc9FN12sfKGgmcfLMFagYQh2ZG3
uDyFl5o8CugANEEYJcEAKqNngnE8wo8Yy2yu1kpuV2ieUsymXBRbK4hg6OF6xzpahF4SDuWqrDrE
CVdHnH5Wroagd6XvZULkIFwB3d7n6t19IsQ/oNEnvSXl0ykE6Wtnh1hA2kxkQiDc78p4QEAtHsdO
ekYRzYWy++Ac1vKIgYf8pU7o7/Bm3wFivA54qsAwznJlHd9zlO38HBMjqnyKO2b4qXkFoFkJUCF0
WUA+GxzI/MUu0eIg3rITmq3pcdkASNEiTTALGv72WdUvnOlznROqe6jOhY6D03RmUPFAj2T/Z1JS
VvrkNANjmUtVxdkFLFGshvdqaKN0/4sdckRiJe5JPXQn3Qx5jkQkIEhIHOuX07Qu2JsGlHVu2MVh
3vXYYhysOw1zUOQbjm0h9WqXoo6r76XDHQuD3J0cx6ZZ7a08TsbzCbkq+JppvABLju/kNypd5Phh
dpscH0Q2GPpvY4LN/J1InQ+FkXQDBdkgSmsvH/xBpy7h+si5Q72EUa7UWLn0qCzhHdD6GMP0u5QF
RF1ISw2YCvfX7tSCNcgBQijvANgiuLDaoXvENlrrTVEB25rnG+qBR6e7D5tkrIWyqbCKfI5TU1zf
GXwCsdGcwfEVZ7YudTO9n9gWcqdHu6mhg3AKvs9C1Zw6vWRfS0X2APWwUWQ2h2NjZ4yQXrQvLEv2
/DgUCrUhFbww95chka9BzjNO4aipm8UXBAo8rhveg4uN/5Z3bXLVHl8J8FkxbIL3hKolOzwE1saM
kFxNibcDJD8/J6Vp1Hye9x6RM3x6pUaCdwV+fnwNgjPolpmNthB2jNYhcqjR/n2Kf7P/+aUX0UmI
CbQne+HQ9m7IhEq+Gfz+cCQTerZ4pvBPwzezK1qPkQQE+6/HMZMljDl/+xZtCpiU8YuG5nyKraji
KqNChRARujDg+84Uc2z7JclJqIBy7ZQAo7OMCUMJreeEFfmsBClXvoPm4akFGaCzqFSpPkmoYwdh
DJ7Jc3sFjnS7bMXADv6+LNJlY2Gjtd7T5j6h2cX0ysNFkgf4YIDfRuk30wCkrg3KeWIvSKbGx5Xn
PPGKN4sMp9BjX58YOgcZqcub3eSZZgO+tUBWDnpTtdlvBEnOm90890+/OGUfT1HCgiunjb/HU13a
YvC0LSntTZvvaTxXtvB82VHoBhKiEJQgo1OWPa6YvzeF/uI5Q8Dg8y0WGOV3ZWE36dPw54r/G/+h
Nx0xs87xUZqLaOo4A2NfFzilmyfUei8rTbUVwabLiNHNL10cRndQ26ExL8HFoiD1GH2rbvP0HOHi
XGsbluvSuZp7WHQ9rVW85tcdxVMG2GeNyiq5KA8HH/Ep2Qqch9RxEvMzJkXnmmuv905P1gkZrRAj
a1y4A79ti/mfieocH0i+4+S/V5oluXRNUGVG8DwonFj8ldvRAhJAc7uWzIPn8ofaiTBe3ZQF09+a
D6/DGfuxEYQdCkzaxscL3elEwa7gTN3OvZcFdmKdtlgNeXCMSg1HtBPe4QKx+BbmxfSiEZDyIaA5
r1Rau/kbb7FxtKzk2o64tlytIIX+flXxz4dDOz3xFprAVitusHfINR4niHCE4Pw3lZACNRjYoJgM
Fsq753GOCgpJ8AIzPb654zcXRGQHQ32DxtfUvWWmdB6qbNr1ANtDfXPmtD99+SY4V6KyuBD5nSzS
QDDB+xL9FJbS4hz2G2LIs8itzVhaHjN5kIuMdmvDKt9rwEoA8FAr2lrlMsBIAEEv0thSiNPTISpJ
nWannKCByvfgnIUvgyHZlH8WB5f1Ag/Ltw+XdmfwgXbkUwzt5deV53nlE1ISBoYRuzPx86Vg1p2u
f9HEqBs4avyF9np6KyKtOQqedJ1I7SvX9vmBsQSXJp0EI/jiGXcN0pzCikO/ALCwpvNdVFtZAgSE
4hyDHk8O8GrF5eq2drMuFIXKodZz9hBUKs+rGa410fFmz0nL2k/ipQsz8WtRGeS4DxVoP6vFQPU8
88hOrD+qNY1aM4JuhVcbCAOIDNrmhJV8cWXocksXPYAxPwWUScKkaL+NRP0nUhlTeRh9tDa5TCTc
CdcdgT7ov0uUCEPhJtbNbp+8OYkvObGqWp+viimP7U0pQ0ZUVi43p+QEw+cxtRTPA5h6EjsYTdZa
lFsLPdro1qHYIErlLBArUsBDdXIgQFWILaOrbNVZXwy41giA3jcgm21fjWLAiPK3g7wFQ7cTrewg
sodt7iSsSxaRFk9oVQQjOi+RJAXbP7X4KDfID9KxXZJEYvbN9j0LAW/n4ILEdL4U+PFE0zpX+oSV
0wD3YGJ6CyGLMo3LjJTLSAfKF+kpYlSVuMsC8m0PNw1t7++UvKc2vC6yN8bqGVauP0R5LV1kwaZX
+gcq0aFiDCT3k8ATasUG+ZJXcGBUEF6ztys41JDPJXFcsb24ryCaAu+V7j+0H4mG9MaoxLEHGdPW
EUTjYOTEjWXx4obgotM3K1elv7w3HaGOKaubRFGtU7AzlDUwa+CNOlib9Z+nY3WcclVko5s6PBwZ
A1A1ucL2iOgYnk5sgmYCf8/Xdl1WfVYLvjst+UT6NTWfxwDZgy0AqDhu1e0ePReB+9rl346xkHA9
YOU164hsXucVOYyJzviRec1PzcopSvjVL9bHiXDi7tZxuhn0X8sd69bJh8sNIQ/bJwOeRX5iaRvq
TERD/BOtJ0bxrFxzFV97FrkqDJcYE5UlhpYmhZgQBdA5qv7OEeOThJ2z1Vem0VSKTdXhio12L4hf
zX8V02nnMaZ6bq7vhtiUJXQpbot7532GD9jct17/9IazAYTzA8e7T3ZYmL38plXlGtwfxoCvAdM6
8erwS3zz4JB2QsbOAweBSGBtNE2DlVKSf9lX5qloPeAXUiFrJcgVjPAlFENYolkGcxdFbA2otJIh
hLy8Usl2oNRGnkLuuL/TDcIGo22t7hFzRAapycQVbTvVbd5/GoQCGbV57wy3j59EmHYCPq3bnzG2
gzv/SN8SwNgS/hIm6C1lHzIchir+B21lP3F0bQo6XzaVCK2oBRefBs5Inndk2XnnkLkgAnzJ+SWU
L08VtOmof+RZx0W64IROG1hcQn6DTR2Ki4VW2mW+wGp6Wyu8TG30U+pcPRWqq/yFLuHWWZgZXj6n
ozfYQRMq3Sw1s2stlbSTs5j0robk0XrGKB/LcNILp1k6x08WoheNtye7JilAyAcRH499V/2nKAiZ
6VzZmPx7xFAB7UpWg/OtcKl8d04SuPNIoh8qXgXMvsfmmtB5UBuG9KdlgNqrTB9SuX/+fWoa+KQu
YiC5Xs1Hxw1L5pb4y6RXBfySiTkDpi4vEW0qrpKYeZM+jTaJ1xhtrFH7se1zbJXTlYBGI+GFEc//
NSL8YcOzW9I30zrxo6XyYPq9wbSguru1jZuqzwDh2rWHHQVJRjGGekhW1H5GZjjZ8exOvFJ1fiBO
jPvsgkVjeX6ts/dlGg2gbff3s8ICotQofETeTEh8uVsC55vazNPUWN1QHdaclxMsIWHkm7ddDB/p
BtPHLXq89ioj91YX1WjfjhZryugOvQMhKzS7I3gKJaha46+dkRki9850d285nqYUguoDU/bD55UG
9C8WwWZcjmGkhlQAxRTD4yiFzADAq9CY4WLMghlaANpzAV3+W3KutuU2P77tVEzAjOHKNOurZrfe
BdzySKej7m/hxOpG6IzeO+o3ZvDYYWTddAyqUe3ZlE/39cAihnTt8eyZjmpA72UJPCoMwhfLAe7K
58qdB1i0EA3nM0j8zJ/FLlt4W2HP1FjPw24OUK3OZz6q+bnJTHM+cNCIajDhIBXOV3oOUvKM7EN6
WS/2kW0O1kER5yl6OW2FtYmG+vYlqhTPKrN9V1P26ViMpqNJP4x1xE9XYy4EgwKPZkh2wdxkAqqv
ZRY6yoUM0ZehQVSgny2IQNgy6qUk5iLG/ALSh02yVFhryngGuJSZySZ+bDh1OnZCr0ocJxxYoafJ
jGlD6orWH7KoBgDzDp2WZ2TBQrZafc0JVlZJEJywYpfAKxfr82ndr6h3kQUnpCB+B0w1w9Lj9vin
GNQg0Py/lczuNPop0ar6AelnGPoahtjRv47l+4nOqWWqEfLt249GvXJuULFgpKxMJ1jPOCAj3786
8bhQDWifeBqJ9ZQMqf25rvOtyUpzvs9mi2hWYvCGYcFy3NGiyTCLQtaV/8uHjWBMFK08iGGNit06
BX3ZuH5/5GT2Dlxt3S/7erdkyolV/jcknpcaXHlJQPTkSMcmKzt70H3vs7UcCznUYPn7emfgS+zn
JIs2J+EM82VtJ6f0us9TRWoiG/4Y7iAUJZjT9LXAU2uj7OQccF4WTkwx+wUQgkR3kEJX1E80rBuM
LHw1eZJQy907Rg+cpEDcOOeyq3uKzeMmBP+RhBxl8KALI45BJsEM/GgH98Lpj8MrqBXm8JEoY6RX
D++bAMY2forULWKZQcoxd6tOpp9e/CKeuL6XiK/JpYS+ObBuGpY1+Krax3ntxfZkxy0j/cfh7AuD
ggqS40R7LEdgfPnBIOdz92g67Ch0AwwL2lT2rVRj4mVXWSML2HACNBy+C9t7ODG57uh/CrN8hr4Y
FYUjEtmBL+4b39uuNSyQ3V4GcnyHGxrVqU2+UTeOjbfFbUYM7G4SFqy5Z8nTfajtBRN3qBuwPbFl
02xdzqa6Lw5WX0XZjmvnWg5POU0yPQ+4upzh8fgPcQ30jgLOUx7Cq5A0AfeIIYRu0qJXZ5eEYdoL
LrYxrqDattY9DqWuVPuTgwB1ChOkGUf06RVXp/zwZMr0Lcy9l6xxI5t4I75WDgdBP2FT9cSwsc5f
fgryyl6Dmr1csrFK4btNDTy3tMx5gk/sC2G7sG3ZmhX+9xaDSZ/1hm7gpRQ2WHr5rLgS8TXw9KsS
qA8RM+bBEwfmNuiOeJ+bSwuVE1fIXrVf+gCAFQyG9IiTEM0GtNTZQqt1IF8oIrsenCAh1Qns2EzY
KPme4TXPvonz613f1BqMxLVCJVlPN6euT0Rl1YVCmJY0fu07kviESUIL751d9gbg1lqqvjGqXXe1
rUxfIkIn+lOtxQDuKr/6eN+5eYNVg61/ugu5cMVJXMSPySnIhyY1jPEbeGZlxvUJwVcisRjfc2ra
CDqCNFdUZrZmS/icVC6vvx9FlP8xGsfL77yFYY1cOOAiNoNkL+Rx2bnD2xs3SiBIMbY89u3/K/M+
oXzst9X02+CAalF58LLbqAVnHIwR0rcku/2MY+dQcsPjlNHf0fSL7tifUWX5Qm63dnROmWrjsNyT
7AlYZHwbo9oa5eJz+du2c71AaDB9Nkv24Pgl/BMNAb4gC3T7PbcaX5towI/29PJXw4R2U2b7xYFS
2ojFk9sKdWdCHV3L3+B3jZN5v2FFpurP+t4/o3w3Z0xla+etMwXtcy2TEoJh8ZlgVa1U2KmVMqwU
8UTt5Kjy3+dhkO3pi9vp/bjZwZqlKqHxbOfr25COZHLVab6HP4kKd8d/jGdwGubxIdfPy3SAhrML
BAe/Wyv2omxf4/3FPdTmmrskkeC6wkkj8X5snSgU3/HqfdCP3qqDifHYcER+FvFqjFU8gXT3o9rt
3CFmbHx/VZfdVAxZ9jjgAcN9tBW/tFuYZEzWbyI0nTy7ndMGU8w80rRhPjMhuZbyiEvaGEp2qAI6
/MVzKDw+1UeoZrRF1Ns1aG06Pm8bhyW1m5sPntUOgbpE35w1gesVlVtbbPnCW7KovpjwryCm6vBq
A8YCLBXwGzmyI3avQkLDlAFRQzqiJ7k+s1PAtE3IFjCPLgBkO+38jGN0nsReBQl0nvZx+OG10Jny
UKMdsCWq2lX2CXh3mgkOJRfrFKETWGK1Lk+dvEJvLD1tsAb7d5auzEznI2rP9m4TKSO5NGCRt3G2
dYADJySQzc/gDaDt5hhQjTyvYnEPQ6pb9g0IFZ8U2VLXZk26EigXweFnTlCXgbft2EOmIqNpr44I
MX5fhdWt/czBxnMycyZfvcuaOXNxRYSf9/qIHHDMa+it22R07i7yCjw7+WaZ4fMBzr5r0ATyv0e5
Ij8tOYoyuPEeM763CQ38SLexKQIVorWG8ib+DtAwHpWLApCEKpTJdX2EIVTxGvon5QC5h3SE50Nu
uftfl8fxKP/lj2/BIzl27ahXZDjjGVwOxqUOsTMVrIRIuJRxRP2QYpw58eUKpWIFFv0NA85QOxeh
WQNu5c1G79yIk7xh9EASWO6oOR4vn8guO2ZAzTIr9o4Gofbit1ccxP1AnSVBMEBUdOmcQQkmFqMv
l9dXnPKjb5UTYQDsrqyZTgPYurckcRx4aZvQu9xmurmfCH9u1jxhqfqVQdBEwEFyIAOuLteZeFrb
3/p7huT9BYZmNVsRS9hJ771hA5Lan+4JMko/FNRQ0+lMnVUrUPMgEVeRstGgJz6wahc46ww77saM
Ir2v0NpCMFhyUKWrf5hEJvJnBtNsknEBXnevS906qm76WinWkHnCCdv6TBAz0I/sG5rzK0LfK0z2
WewXJuxBTP6Xq/5OGWK1fXqF2FtYfsk+Mdoq9/RnMBatJ8AtdaajbGyAO6FNTnF7OjVqF2yUlOTi
HO/DocPnDSDl7chyo7dn2HWrAFNehQY2BD47pc6YP9eQnMREBLCdXvxU4BCKoQW9s3fWrtLu+tz1
HOSxkNJZTJsL6/Ziec9CnXdzwMKYXSdTIfo5D0LaZa5kIQhrkZQweLhJgia9U4numU4yUFx0OGI7
dEi8CCU+3kL4KZDo9+sZ3xncP5rj/A/Mbp23gcFSVhOvxM+C+9Tzy2qxLE6nnD4j7BiwcGT04eof
ADWZ1Qr2v0kfWKxoTlERHVXSZeW5eIOQjc3oPl6UV8Ok4Wns6Fv8DLBrpP0XX9fVvgQYe1jsv0UD
IOlY0sNsOrz9/EgEPutKK0Qhxls8ptdrLoUxerRuXjMM309yKywv/au7igKASZQjQcrNF1bV6eEM
Fa1YVzkjPNP9Z5NSGzEUVc3OqVP49jqqDhjSfGJUSAK6X5qSRmh7dNjiTeH13ckKNlWQ7sX4skHc
xK6PcHssoGOX4iKwXv7HRRQEbpZSqDYja6Y5CewG8pD/usnEFKiBznuBXntktVGyVuYapFhW+6bP
C9fZwdXq/b+HkOzRJjCo+Zlt5FhjrwMMpi3XDDoLKxN7+bupPsP25qz6TuauI/3Za7FINCQlGdZl
0p58X6b6pfzrRqmBABO7qci38PCCOGJWGKT5Yi8r5qSsPNQviTOjltTwlXJdjIEMaz44jK9CDeo6
DB2BbQjC67WfRnHaOeFVNE1gfQqxwQn6GeV+SYbLKykztY9QHUNGENPF1AOa8CWNGgcNbZRdqJDY
NROMSLbYlgM7zCioIOWqXkcAJX1i5jnA7ox7hZ7AZAw/lzEoBj9TGi2JlID1w33ER3mBQphz+FB9
Awy2hipI0EExcOqnGsrmNTKk6h4JttaTtByyNGFXs4IZ2FCeESC33S758Yc7Zosju+LnY2WjofLw
FN/gpvdyL9uikGw9364/j02WLp0ydxk5wbA1Z0wo5nQh3QEaZgyjykX746Nilt5vaIdu0K9B8r6b
p8sT7uy91swGSONnTauZNVWCEkmvqrjSnXvRtTQICme5SG44cGGpBgJVi01xWx8tJYPoJG7REsys
ibcxe0nugHfk0s/AxKN5k0cOUGC9PBAPDU2YiqcTiHuL3opDYyolB7wkMX7fk6WOleAyhxuQ1U9z
vTLXHQNrm5Ta+6jBjGuJB5YY3DgccFHZNJ+Rrdxwt3XmvIsRPAmMJ9PNtmO1hS41n5LtNiHXM4Cp
+yXyMyHXpvpUKw0Ul/okLJNP9tbQWjFmbW3I20F80q41dsfOo8P85mbd60dlxtKdfGHWBTviP/YF
D19h1hThU/v4q2reJUDsu6zfLkIpJUpHaefRxsThzqZnrPGkJe7M+gqoLlxM2XqUz2rq/ghTyJ/5
6yxOfJDGQyTgadSNQmKXxzM2Q8RABOdLhkncqSPITvpXmE0a3BkWNscVz+WZ8UU/7le+I71gyT7G
WhQ0wakV6KPJgnB8Mfkdw49mZrvW+7whNIUcnnAb5E1DhirZP6GCBjdQQXnGBb6lcifAZTscVV77
BBqWb0MjSqLpS7ay4F36/QQaxCdQZxpusmWQOPi7Kd3ENt7dOnQ3A4rfwQSbnONkEHRHsGYALjM/
o2Jr6BgSL8akb6VuVuJUxeW7JlekG6oBlomqDMobD6IQYFH7k1P5RwDENJez4FSj8XLUq7mokctI
5pcPj/XnVOE5LBmwjPbejGtNZJ4ushvgTs0bh7C0z1QYPLMlq+iQup1LxKRk4YIpeRMkGIxgv9xr
kddEYUxcB1GNKE9Aw7Il61yaZ2jt1kcYOLvy7hroy+zi86Fzd/ql3Sq5bEoQQJKKu7o9VpbNiDUl
j3bPUg/6IGC573t1VfI7KQawW27i000WC55+UavbdFO4hYMUzpnuOnAPDQ5fei8hXaq30fA7Eenp
qOFcFp+n7yQ1MMkeyvPMZECB0scbDLAfoaqb+O+Pt0ifdtrt/lCZzfw6VfGDg8/DWuMl2rBSE/g9
V/fK4uL9jktqhEqO97RuyzxkL/1DnGUWZtIM2RnXLuCu9kTHFjgf+dRYX+1a+kt1SoCqLXlGM4Jb
ROwYmqyjerZg+eePL5pXVaw5giOUJtCRQIr0NK7GjG56EZGuIarg2j7SCQbIH/21plMjVYaOdfe4
EaOMqAll3ZYymFoU6EcrpfFTQpVVPP+4V3F4GCJ/N3oFnwRXjGGLqWDEgwwS0yCSxgGRsPS/6wLX
iSj4+QwGbzO7QulprKv2ffl2fLSEAMgZgoPf2DWHj9IboAJLJ9M6Y9vn+ETFwfMt7e/ldPhLlqi+
OwMVQQV6/iUGiqCkSEQISgZqD4DYUxpjSNHHsVIkqHn9St2vriS6Z45eqIX1bIufs+7WJRmZtcqe
LYQoV5Zq+mwYETM14nc1WeC56i/9cQ4B34vhJidNmS6Kq8gIHIqEnaBsQLlw5bd4pG4Eq0hxCZss
X6zXbIZ/dhz93ST6Ng4UzRjfrCkW1lunBHNrG7n8qpa7+PrgYz+OJiLg7wZPx+LTDBzQ0HjUqx0y
tXgRlWCZF7yIabjOXfSu8DYgPQiwYrufnroA16O6EHNqUWMnGPnzmEdPNQjALbV1ps4GkYE2lTEe
kFL2tzR61Bbpty0hGk0/9OT8/OZge6Rg707XuZEMPeF8CuwV7+v7muCuK+xbBaELf89MnPmUzcuL
dat3HO0ADz5NtC8p52YSk56O115A5ip5jODIB2q6b5cJGzPlzw6UeUpkWUj4mJME+vzP9JzgJ1jm
XC9MR5Gf0QbD+/8tEe7hMx7KzucA+PW+rq0XrRDdQm32tbny9sK4Dkm+uY/+VJRrADC6Ns+HW9Nj
U7gabHvokNN6JsRf+ZP48jyyVTXa483h5IZ1lWzKN3jXcuXCm6ZODAfCmPiolHBLPARhCXIDMgPi
zuVsHY4K8Re9WlgYj4pNPxc/USliAs1wvqVIA5FxhkdS78VN0rt38q8RC36filCy2AIaoNo7klnM
pj8inDBIN/xsAOCi5xSqOL4Zko+Zxvt20UpaAf4ieN+7CzEOIiMpBTfFmS6SprWDkbkb0S6bXfUL
WveXoR6l9Vge4u488ts3rJM7IEUWg/5unoDIpmo8SZUwTP2jkMQf1M4CRyTSEMMZeRrSq9EH5GGG
GxicT2Syo5Won8XbRJB0FDW2CKizMZkbr14bSZOQDBkYDWWsQcZsmZcz6gijxsIibvf6h6VoApNC
5MS/jxhWdxJ+My0+TV/LyVceLexJvCixCrvAGll//rbl3cqV9foXC3eRGvgm9V28vcdqLZskxU1F
AfD70NSzPvqSLnIIwdXUEhNNUXeQzx72b2sWrUBZ2SufAkUmRW0aUk1BaFfewFiH5SXlukS02Czm
FZ0GJ3Qnu73Oc0H4dtddeRdttjx65WDO1JzjYPwRwFaItCCERIxe5UOlHc6h6w+B2Hwwm95AoZmx
8TBX9/YTKjfGKMfBloCJx/+k1Xo7RGYZgXolLVcazXHWaIjLAFcb/YXeecD39MFMPWHtH9KJs1am
75tANaZNQXIrHvIBIk7NCZ6PnNl2i1+bH7zlgxzKYDTfAXts8kXHoqAm7fnoJgoJWof+v4elZD9l
Fy347dIrg9RSO4YCuBKLtGzRl/ulZskLaDUARz3Xn3IyjvO7rAZuP/dgdXCbnWoDEcgn4ZBa51Ji
MCsA45nQjWKEiFvSqzwwokW2OJNtQCgvWz7eY8FnhgQjmkNlO5PhwfIAyryE6vn6L14GI51CGGOp
oJml7NEXyUJ+8cLvr+uodzCCiWNV1FhcP8s/JidOLpmuc7VRZ4f0HU8wJH2wrNCDdAhHLIN7wVL6
hjbZkVvt/CdvhmBPIlOCnDMkC4EjdrloPLPlsqjbBQlgr4Dotd2SmhHbtjnvX4HrDbhPhETIJO0I
hoqtYMv/MugFzOneJMUVHlUPXG3UArY/L2UtlADdpenz8op7yRVjLePOpeT1R/0oDgqEH9INeqqy
q2h4U6C6fV4f1mMyBwz6yzgE/YOv57fSsyOYWrinrU+4ZOB5knb7o8kltN1rtBSbEZHsCK1d3zQX
VjPtdFiABaPkNT2svAKOtdoMNTnrRmWxjEEVPKzfGp9F+9jEp1fpRT9CNLz1igaeEBiEZk1GyFNJ
c6ARplc84AwSPQAFABXeBeyoqc5fs32ONitI9wHxVP+MsBI24uI8EwGZS9d++pivzx09/egSF87k
GW+GLL5LAADQlk7tA5fFTdawvZnDOUp7S9hp14q/1V5NitehmEa12DHc0wBSZV7khlDOTGFo880l
eCsvBWcIy/pQPrnyaqeDtVmO/dkKqygbdhEBV4KNirNWhFLyfplwoMbtZ1bCXJUm6lp/xH8Htrfb
J0LQ4DVy0ZWXO1XE/C47LY5vHm/49/VO9nOnTFuF0CW9Rn6sWCrGY6wWZPAYSbwUwLOysC7Rb9ko
FUmsKF40J9bLJ3x5aPzoUltKTYydvNEXSYAyxod54hbKWBxmIfkbSIuek7PkVsr1aI0L08sja5Fp
WKrMKP3tA5XY4XuZYaMebEr7TKLdt57dTtyFAiIDlEtqnDWLFaSSUEeZJddoTQd/Njke8i5gM1zR
6mFbK+1jD3DgY4TrsuKms9Z6B1/9Si5c0FM9fG3m+5sLR2e4eObhDLmvEblqTtWSZ92C4eBsjwe9
Ln8wDeT7nkGPncZdGm9iiGGDbZY06Tb1JPWUD0VPpIoZDMaJTS8g9jJ6zyXKqd1VOMk/r0ZXax5t
IcjL4A898gH8j5PUVvD7DyKCb3hU/ww+yd0DlkWD/2YoJ5LNPy2Y/f9EyPeghVP/N71eblsRlHj1
Yy79uBXJ5q20dHmYzuyWJut8OHV3CbU13HjwnuXSmCQ5UkN0qHXAF3Pv7nRCI0+fJO1hsclW9CPq
aN2uWg1qTlZlgJUuhiqvASHCEurbXZYXc8rUlywkFFVs6rC+vWJG+L4YZulGbe+dIYZ83fnkptJs
LxFIM4RUJt6qdh1jXAw8PQhS5s1kmigrT2/fsFIdzX8Fd+kn1T8qokcD/S91zTH+aZwM/iCPI7cb
Aug7uVinCwmbikWD79AvymFMEzENuUiQ8ecMjl8p7vZvUfa6pGpv02NouJKL2IChmrJoP2ervPC5
UMKhwps1uLIUuSkJvS6aJkkR3tlGOKIY0BSb0RHyhnr8KVIgUdRUPKNWdtYKpXEYZ23QtJkgqoSS
VHrmNd9JH2qwk+sCDThqz77UmMSFfyeSt8DbUSBmVqmn9OSsr8DG9J0IMWW2IosxxqnsSxwlaieq
j4Du5f9tUh/16FYwqBAuI7ciP+SLb20avdiy7JYEC4TC3/xNLKOnh5AjHeKaHbSozHYifKJLoT4V
kAFc0ATzMrtlHEomGwKVm5+QHhxfrNexNmK90chwC1D+SAHeKCYqioooNT4VK1zFb+BkxitfS0qD
5d5FpGdpz/g2yXfuVQLw2z2lhDXG/pQOgNKx81Swx9QDCm3soMB0hk+s7BxJZCT1O7GgywhbHLIo
tV1tULo4gD2US+U1khlam1ulreXOrYCzvRG1NH1gPGy9eYAsC5b6Ib1cvTDkWU2IYqoyb+R6tatq
hkrBgNz+ZBImcalORS+W/g2uYZRcPP0pa+ewmb3drebiCENaYQUncpRbtb9FsDpPQ5KHKa/MeKP3
3MkdUl+2Bi1Hd8ENKjitcpyh6oziGDOoi/2+Dv4bYe6PPIhtpqZkVl8L+JSYKBZQw//+sqjX/S+w
MA/0ShHXRGO6ofk3YN61N74vbwPgV/chSpgP2sYXi9PVKecrTUcdQjkcTWr43t3LzXMV7+OY1EKZ
pgq5kr4By9itMQW8T6vvuFS0L/Bkdhp4eji6PNzvrjfCu2jdc5gz3t35+c0m9U3/1nAS6Cq4RrzF
+H2EKteMOC8z5ahKl7UPkCpXTBhV0AIu54WyI+lN3GzPvy9aCNFbA5dbWvTpk/Sb5hrosnNCv58B
D55XqAckY8m1ZedimjXoSpghavuAejMjfaLEtT7LG51fTKozFCwBYWbofkZfbB4Dlri5Y3qZLXzZ
aLF6VOCpElYWooGY2S7ZGAnfegeG61TBkzlG0BmcKPaHeRGTVSfDvMLU9fug7dG3m/W/AXHvvXGY
Jf6uAeQF3wu0EEkVsp9HbCy5ImAcX+/PUSIh1AJeOmO+YurYaACDBDWmIDz2Kqnx+Wojf+YSamwg
aXzRnrzJeJVR+BzUa4wykMU8BqXHmKGsptHhLnToDrn0vhNy/0nDXaAyge35Q+cM5K0rArmNtBGT
zqdMDWKlRnqvM+8WdInETyugKpoPupUvcgs+whrUz6wt0sY++LU7xYFeVXMcXhXg04RF7lmNcCwK
HNsqeeajrTLzX6KAtGqFW+BXww6m5vSJRm3V37JsuYfWa2kCI08uYN42NgzbCVXyHGre1sDbTx2x
2HhkM36jjAgGzsdTT5UKQKq4ZFAr7qH7SL/j0j6mu8tPu2Ko4pXQaXsPCfb0JnXag9O2nM4UqGs1
AiuXR6wSuUm3DfqJsT7078RygmeffeILum4iduMnBdYAdQjhOGyrTEl3pB95g31cp6ylb8n2ZV0I
WceknP7Dm7VjEq6wJXnQPWhMdg3CAcOpGE9wTz4trrMhmub/vhIk4gXFAIdqqKmkHE/ekO/V0mdB
w6TzUEXSItc7LFilHggshooG1k4ZA+W5CxNXA0EdPWHYRl7MpVTvkONdEeIthE8empEe4ug33Ot7
9nPgqaya3ujtalV5DlQfJlnLsGznkFKxtk8suZG9EXznF6G0E2xEeifamxiV3k2SORsRVudJoLnx
8CgzKRTIENM6bdpRtMgeFj2O/JeYWgXbitVhYhu9Ihc3tTw7iNomeg+CeFisb01+hafHT7O3xUoU
fSinM4oSxCDD8XcIY+cVo1/6qQjh8HtA4JgqPPz9OmGn1MfKkZrAioIFn+E3B3+cxO63WPHFgw5P
BtU2MQ455yN038Bm7Cfvq3uWGfBsR98TF7XvGpGUKeZ8reN3kEGTA6inegqcO39h99Y4rcekFAq2
rEgog3r7tFlpoAS+fjMjmQDusQ1o6S+vODIHklyqkXEEV82QN3EKNuixkJqtxNE6PZcEGTVY6elR
hc1LrkpDlmr7fV1OgRbv3s4VDtd98mZRy/jF9HVQTa9EIBtXXnj45A857N+1shTiw1P78Sp1Gq2r
A6uMFVkq56Ka8xRuym2chOuzHStwwufH0U2JysPqHueN+q9MXIFdB+0L6aR6PTvCsUjeeMF9fINS
M++5qdVXnbqVwTNRb3DBBOcRb6FAbtkGa/WD/WGRFz3//UWMmAZiHr3dcNI8O/1w6JpYye6nmGjj
8VYVJTX8to9p7CeLMrUElf9Dd48hZ8BjdZeWixRYPjqLYEVMTxhwRaES0M0kva+QKf+4FLybBwiG
TN7/Ac34VBhK0fcsHvQudRNpmLncNwqjIenO6EqK526uu3WmET3lhBHcX+yBmlKbGhkcTIpfumjm
sYKuinFu1qYRNzJkUg2EmFqsIEvWnBnZmOCV0ZQc+c/7EuEC6iy1J3zyQHUD/vNxu2zcbkdOYfnm
pQ1PyvZqXi90j3A2QlqbDNyuT+gOQpK4zrOzLZyz1MY7ckLMeeBBYZ4/z+h+K4wviUk6fn6W1RO9
rEp9mXq8VI+xtPlS22iANkotg/T5SNyLoetI4bRyZ+c/3CmeoehuSpW3+BMfIL/JZTrFQGsKznbJ
N/bi9rFMdePDJRijTpxDwWCXYaZsvXEfBtCKvqSf2Jt87r8SrQakECvhH+10Y+pckiX9qDwhUZkI
CjRD1PA7DoMDdoS5C7v396lzYMSRz6JLEnbOZtxynsSj/kP00rJmz4nx40W4hbpakQYwp+xgflfU
oLOKJqD9zGfjveHJrjC5s/zoJyFXi8nmHM0oRQm7+VuB3tgwRU0MjLVVrdyjardNKB94UnX+CrXh
X1ZO2u1cCAsgjj+ZdazaUIAW/Yf0E8kym/2fsK/6/c1H9FxBUk/AvV0YSTX6dCNW0dXKJuYGGvo2
G58Wpz5dzEM1xrcjsIbQBhqxuu7xYQKdMqCQnRWjYl1ZzTIzmGswYZx8hVu1crPXv7ZyIAvM/18b
STx3JsJgjzkJv+ywkoqOrL7E38lU83Dss1Ei/IbfXpQ+5i6gLjp7xcL7/M4O8X1MnDKjQBSTFbpF
AuT4GdRbcDUHFhGVYmCmjK/5FsTd82Lv384jrj8MxgR+abROT7ogVfHLa3MuI888u/h6dUkEuApD
HZOmv24ZS4nUlNK72B/BHiChrHkgPlUSd9kAe1bix5MJYbLrY90kmO4oUUlcM/QCWFx6F5L3l/nQ
rdo4zZwT3oasci9fLmU08hIDyXVaNt51MR2OKUWNQ9HI8dvlB+JerpjzRI1jQDjVhwkwxc0GU0R2
LfocRd/XqYoldgrhaNN/1dV5l6iRnXWy1eLNh/IHF2g/wIeBz0SBUvAVOMTp/zXUo/dwTrPl6DVL
ZZmkoQoz6mm+ZRPRGcyvV1XosGfXtoukDUq3VOcs/xKGrcSCdVuOPNZgImK+x05jhBfSnQJu4Vtt
U+sdwD7z6RxqP9IzFtBbSI5J3ZEoyY9kM7TBcBSbEovbI/oHweXV3ovg+Ry8g3DlagE34OtzhZz8
Fc7FmEYcm5XI/9hEkuJUncPILyTymf9K4yxagLITiBiz3aQkZZdjD9QcUzK/82qyXN5yv58xSuQy
saGNtjJTftGYoRpnzXUwetUxaiNZKBTCcDl7QQRau2+NP0fhNfMD+2H1U8s+HjULaEp1A5/S1z7Q
g6dNOWVSKE8n0NjlStfH/OAf7GH+i4BI1h46FtByLI5vSNj3OQ2NjCKa2ztCcQofYWlIa4MJr+gO
I5FcGevITGN1Am+AgCiGn50dIrCnKl+2OIOYc/hmGwtmvbtU+V+o+MEpgzopXuiyPDGuJ0V18a55
nTpHYR8kmv1edXllnen/07UkbJ291W0l7zAb4/7Pz5M9CHiNZDlmJqKiuMRYQLq4nin672ZBeQ+e
xTvveYA7orbHO7eweJPvcso2lQeIhioE4SkKb46v+Q5I4jkxYmXNn+Lpx65DUZ6cw4aFZssnjIFJ
oEbS+261ur4yrcT14PV1z85KWoVBQnpaAd9mn8YIfoyNCUpT6nPIpTf4T62NPqbuHNENnqtcyEl5
drUvJS5MBwfTLtuPT8bE1+355bG1kkpR8FfRDdWbe/XZT0dCjG6Pdc80dvmBCGhS5b9+RNmtGVuo
7IopJrUMG62ooa1mj6hmDP3xf7HSr+2qa8z1/Er9jqgS2guRpu+OZhKBK77mCG0u+rgSyF7mVbUE
xaiKp9T+atuFziIwXHxgQMiBxBPB/ApTpSAPSKW/xNVx94w6yIt5oyuxKGNEUZ2Z0Tp6w4s6KtH6
LGW8Zc3vZ4fZGg4/7iTkGmttDHe1OWjz+BzgZdYXZWeHdtU+hKEdq6t8O6MKpg5MmZ3h9gKrcBAe
7ZdLcse3W2lTy+Hf43O/FGITzXIQCjcCFCga05+SYycZp6Jlhej5/6DgHih0Wtk3OeS/YdeLqWfw
JwAMDw5hafNaJt8Mug/GDjGvyJeZuiJnqbYXNX0ps0Tn9sFxRH2YW3eirp92Y+bDQ94DlC/GJ0+M
xII1O4v8aX9/SVedp+aMs+4rdx4ZXlnE6OHjyU97LbDgylet23yPTgKWBqDS1//0V/kNi0Avvekd
TaCmlmTWBJ0F3+Dl1gLiVICJef76YsiflvfJXNRNUzkDVmM7L8mhPGAdbfiLWyCh5NWJAuo/smDs
atC7xN5/j8EyeM7GLvftR+uP2pD21OtAXG+yOgQdI/XkSRu3DFAl/lkNCC1LOTGadEZoF/qThLbT
FcD1pl2asd/8dq88b7EomWpHl9uWGFKDksONXbnjyVUFbbeEv+dqrOKdzYSsB2Wk2lcbatCAQidy
laf+JwCyXTRfwiysQH3d3AoEycANpfvv14Sf1KKKgmxNxtz7sj3ambKSkeRJctOUwKicl/M7YNB3
+EcgjYFJVPPvs6dTNOvdJU+m0ZHF5f5FZ4RtiHFROyAs0ZfBo/yBU/cU4sVyTM/vHrfaRbaHoPeD
M3jXwCA6EEKXWySVA5hOzkonmy/N3OHTqc09+10yyLY5eb2FQgLAaJgYTDIBoV/2n4WnmEuAosMv
5VlPER6gRv5ufNN8XE7Cfimdmaby37fVBxxpCyXeOiJPI6cuiSCPU5VTn+lVO7QCorEBwuP638CS
+adzCfbeICQlIj6u42aGRuw9VumBPO03/svMQRxb5QYz6zxQflhj7TC5sJozxIVPSfSK0I6u3cYS
rNgRo7ShFAx7g5+9Dxk3WCLJ9U8Mvmr7xSl0nj54RRfym8eh9Xt73vQ5QrodvTpaWuXFIXvaFKwl
6AAUrFclNdeIuJ5rQx/3Rmm7jNYbdiFUk0vUC1kK3SW3Ea4h4UbiElL+JaO65tp9IFQjR6fZvq25
FJ0JMhNuSH90IAyEqLR/OBy3GZbbpSvMVeTHEDhXN4glZEnGCEDExqhMkCb0SVXDOk2PtWkmVSIo
/q5qDaXV4qrw4lIsACzw0Ar2vDPTaL5ykzekvt2H6qOFVZkhXnoDrpX7Fl9aJc97nFl8mlaUOuDp
wvkoCtkCErlDMosqbbmhKZDVEhVrIRB5/1aRXCwJVmiok0QbxP2IJM9seBNVnMDTZxmtTpgwHZJg
4lIfs6AZNFGAWpk4iqsosGn7prkcnt3b3PdgXDLSNWQhXCDijc09i+ZNcproKHlbFiHVJJYtmPfR
BloOLt5Ts2jmwyqaI9+kr9n9KENwcBitPvPyQ4RCvP7MOBdfm4EPmgz6fp9NrRrtIBFrBq3xerbn
8qBxwqVXzl6ok5SHigDZkqVUP1lzqNrqg1uigJu5hM7hVV3nwy67ijRHs0crq9r4c6Ec6dZivCYw
1KQNQ8n7nTbRp5pKcmpxfz1PJzjS76HUn1nvzwoVRfFKDKHKK/g+tY2/zRx9L0C83J+DSGog73F+
kFpUxjLUx4eyCD4HMngccWOq4BkXwUj2lKQQYJusrAh39sC58BcbGD5/6o9U56gcuVkiDF/TR7e+
PekVdEnvJXYRPZDsE6NOb53T1Cnx3GY67CsP0edAIQVJGtQqvFfDo4xZGnLm9pclvq2WsMJqZYAY
gghNAVUOnhA7AGZvahu9ywu98ltsAgUoLDtVsYkDWlG1cEs49Vf/XTliN3h5GV6hhqhJZGxKgoO0
8pzmbUpiF3uK/ph7HPcXMhawseKboRNqzVE+DiKTorXKBZKOaNHU8/xKzdqYntQo9+3MRPD2c5xQ
oyQEMFtLg3TEq35YHuO2mvUUKSHWfrjb/RabXcGrFIJ2cwAvkeMs0aJqPSL9eJN8OzKg/BC1tXhL
lvqHok+ko4ZIUdO0KBSBzOmtiCmbvHFY8cUjKqiakacPoLbxLu3KWhnm82v7eLc4GCGy1o1lCvrd
kdE/3EBAWjhnZG166i8txVoldL0LRJzhSuh5FPmbikx8JysAJVKBqCjhHKnb0hUTeZC/aKjyq0hz
U9afMoXHgu1iEiE/kBxr8ERhWuCwAJGyisfMYdb8giBhHBRHyYQNJqvYz4/B/dnk0K/8RZSwyVke
WrbjyQDz8o1Z8TOJWv5PeYMVbybmoIBCseY/a8D96cbtYwRpUsVO3EPvo2C9n/G2WRHq7sWNwCGT
6cBKsBsxlDhjFri0Am8WwZ1FsNIJnlyo6I5bdisB8LNCW0rpSgj1pmPJvqfxaMpdtmxuMYP4Cnb+
j07+hRih5sv5bDesWXvvjFpGq2bjkFITWBW9FZLNOA36H88W6T4Y9psstcAoHbLTcU1iprkwUKGc
KTm2qYcghLxH5OTids2CQILU5nr1gUHuxRnvkU4QBVyMxrxzVgo3GJDIsG2zkcXuDKQFh9SX/KAW
Y0QPE1396Re0kLc0uRSLMLxshZd6dyow89LRIDdySa8V6heN+adPJMg4l4DWWN51Nu1Hy9E6W971
FR4mVPG610DPX90d/2hBmr8HqUJS4rXBz1hqTHO1Bc9DiLXnpdSTpcDf62yAzMwRpEp1rsP0oO3C
FInhp1RtlcdIV+Bk37f1KipxRQ2KzK0xC4CSiIlAio8xudYNT59/HCtXqOdahdNHcddXMBXFCmAF
h1nNkSpJnQVGgYp60kSnqut+3Czhk9kZOX1e1z/UV3oZ7rXmDbsxPyuhQJYJpAmuQ4W4hlb3dVfF
5xWur2+CovmL0LQaB7T/JczznoFwdpiPkEn/otfeo+xoRVZcWu8Z05av10gP9nNo+bnamLHHRKyv
mviYctbfx2T1xq6eKTFUiuoU5P2T8443UZ5Q03oXXZMzDE7Gucw5WzvZR5fBdK6kFhPU0GZldnWF
DXgIQ/hdeSo7658zKdHtuySz86uCt+9u0+3YW5o0QYBj/0XwwaXJfs4WICsbZTY5tQOb6yrhQ8ym
tVzZNWtf9rPz+6TLi/jGXwwqopaX33SN/aP3a2hwwjQn1rfSKkAdIXROb70VjvoZqBjYK7Fe7VTr
QWYFb/AJqdCCTNox5LbvIPvBUXCIHidP49YkfMwMlnVZHaJbpANxUtcMDMpJNQlecKfVyHkrbkps
8HB/kStwuTBZ1igxCKrcRvE43avSgD/dHzQqnwEuKbsjnT4/jsUlh8dW6gaaKmDxJS9Cn6/+x+xl
FzXEoISsgPio/HvbdffqsuUjT8TvmClZbEQUIzUilzrlkVymPChCxQ7gATDROz0V1ItyFfTwkrNq
rLCoV2XN2X9ZDLqxlVXKpBqDVQl5cepSe82PYHd//utyw31YP1bxByoTCHQz8Wcftd50x0B4tWJr
6QbcU1seiIMaK6kJMQWSOLqKS6s/i6kIS0WnDoJtE+nrlzGITqpbI4pk57UFQTgikh3DuwW61XwH
Ody2xL8o73gvehzaAk/pADd0270bfvT2zt8+pTmoO4qObAJxECDqees9wvf24VkuLIbPJixgEUMA
q3Kai6QLyXniLrGbx4qn19BrNXdHrZcX1fvp7j5W4u8W0E4Qq7uPptwDBs8mvgN/rFpFUMAA82Nm
K+aKWlrbm3/sUICgHif3de6aitYOiLJCTWXqjKlR4tZoUifBEgizVKJltd73E3A8eCNVR4IydrE4
41Le/oizny0PtR6KBgLzdGkhsW5pD3VHT9notQM4/nRLv8T4BcWBBD1VhAUsOVPid0sDIJBkoSB5
DWapPum7gVqgaWEOZgUefQPlSuIYExftHZTTc7IbvTLmNGkMjbUqzjkNPMfFlyTJNC5ZbMJUu2jp
pTXNQvYMp6+ZPAwovX8vk/Dou5C1iUutN/DrMYUvCDSt3MjDDMx9kaMs8KSNQVTzO4SUljLLVF2c
pNzH3CfvxvSn2cQTCKvyAXEIsnUW94Jzy5gfXPBXg4cWZJtlhUxnai2jsMsS3UD+viC+wXXBEY3x
kUdqenkrlC6MPZKN7u5oQTTVNv8ocK3yT0RpJ4PbuSh6yGYHDOWdItX7eKk5Ed75LI1tfka94xl/
MRyoXCNXcbzBpZgY03pZp/jl9y32kVOGyfM2ny9u014qSMHinAKmCNhzyJyNqtWEfnDjaxdYTtU1
AohTBBJwPdVfH5uQR/twFbsO+l8EHTrfPqWUexOKJsSS0tRXuB6wTn9GXe177fdXPMg++BzKe2Va
zgcig2zazHAHYkhy01cIncuX3B1Nr5nnga8Dd/uguVKOBDMzv+MD6VOFG7c7OFyu6c0rw0WctOWL
gz9XTJfrGzYdCPQyPOjVeBNH6Gt6Gd0TYbNDQTNjs+RNTFBxO9PrIod/ypNiI43VY3njjnaY3WVH
Z2oTgtqoZ6TP1FimuvxoBEsaTRCQ+/fQUlYeI5AuScmuqLVbC9KbCoP8dmlstZmD+OOIKscZAk9C
8k5ZMLY9Thvn0Hn8jEZliAJ/OdyZuzZPjSeJogUvQ/OreVqN0FzWHf7iwM0QANBfPjj72SSDFtrc
iA9PFka53kFdl1KHPe8P9qXByEAZuOo4KYysrgqJDvX7sBOIgw7Fky3ZYE5C6K6cqzKMulmAo+Ji
co5URaGO5pHLDdcZDQDLsIyL6P5WBYa1p8rJExcgdQKZF4bSsz8GTzTkFhFrjWYIh8EGl6lU0NpS
Z4Guwhi2Xm4ux+S1epg3Fa/qeRBN03rThXM+KNz2ZpfRi5sPOJ843IyRQL8/8QP3dvK9pqlKLsUR
tEekDTp4vWSY27XH1SJjNut3tjlPBPitX+pvLFKJ3PokRUuXWMloHx4YukakDGLYRjdnus/EGVTL
mSUCgJ8+4sWHS2L6BiI+/IckQ0OG+uyeYbTm4b9LMsJGkhNYgvJAB2rvbXpj6CD96azBXPB0nhlI
AsYxqfOqD3CTqLbuw/DL1yKk0QV3iV5zBWZTePP64ElRgO8bOSQO2CLjqdkhIJAEM7/lO3NIysL0
cAuZhqJcDMfavjIoMedIwFJYDj9+SByjh7AWEkRdpZsK4HeX4wlAlTVCnDuApOOjNi7g2vhNwo7k
DV5eP4+bI2nb7DxE1ON/63jawjKivAYHpHswki88mzYYs1CbjsUcOdNg+18dx2M3tzvZ/YAOORwz
Qta88+CQzC/znj3rSIiBnURaLoSAhq0xq2WZITuTu6exHN3aHR6h9BpuLXm373gws80M3zzpt6jh
+Fcujre7dmD5BLWIda4Picg2A76iHmnpfYB41MT+nyhT/3zjzu9KSO7BSAG3Ar5gUTm2DVi7wk1/
KlYYj8nEEcZVpMpY7pnPyBBSZQHRVcUyB3PUVrjXWfoICf3AdPEzYAgdnhNVKSSddAMSlYjZeaF1
iwsouufHtMGubnDYuBzSUSNx6Br1hX83XzyMPRay4FURs9DztOt4fvSsbYje17DKrFjHCffO/a+r
PEdZ970IKWBnZVREcHxYFVLjslrfkPZoUVddNcCoY/LvkxNfz5I1X67OZFoxZcGSFMjzZD1Mm0/a
6mZAJgJPRTJXzR8sHTEKHUM4qAVNvFiR6+irbVMpm3VETgERpurhHdpiMl2AlOSjG29xhhqTc/Fc
l+tYM/jMxN/hiaRovHI00ottQdgf+aeyw86QBW7AaTRTFTWDkpnmNgdL7TiPvZ00Y3tqFB/GZBEz
VylGA9dNdrPT+1bIxtLYwOSzA/ng8C9uQUx8qcLrqPk8H7MaeqPLiTuYyT1uOmpv7IDn9RU8kdsq
qt390cQtuysW9U+O514FrRxKzp939ygQeAFa7jjOOHsLRd/NRglf8vd++mb4d+M8AvMPGH3eeakx
V9NNE8aZ8ekzVCyKfYknTADLhkiRflQJgv93fCLYcrhF/5eMTxW0A/A3l5t+suu24QyVzv6Ws7m1
OxdSoZqmu+fA7QIp51ZhW1E/ulTM6xEjncvwHyV0Y1IVecRNliktGkbXKlYFdIvji1aT0VOc1y1+
HxUdDktxKyGQpITxAWXUZQCV31a5abXTfpd1HYI6rMkdyr5nldTnP2bVXG0/cosrtAQ9pfPAS7+Z
yzWpLeuoHQOkGRZlQ4M5bfrkWVS0tCunWeoQLyvcbsTfut0P9Un1rRhL6nB3vPIxqWtgRL5IRQ5d
3/aexsHAhv6EGMFn5ACJzS7l8q8czCisym0w/Ml6kVOsNA+I9PVqtNM1netSvTlz+EPVfRlrPQp8
Aat6U9patr42j5q38+3rftj2CHWnpHCfp4HCtc94yU3qVDOOIgi2+/NgwFT8JupYaEPtGsojqvKh
k4W4wxwoO15Lnl0k1kV08s1fLwQcdnyFKsyBkmBT1yPgWvOLpbBeYSl3IX4v+q+/jCbYXrK88cS0
b7kSsgz1tm+wV0fymUmeK5l4ToGRafewQy5bamXRzc9iDKIqCLmIeYKeGavTpb+5hjEfJJco+Udb
K5AHXWQQfvUu7Y771QIwTP5QS18EkKETt0TOmzo6m+CAN2EmYZId9ehIZI2Zsx323gU08cBP+Tie
r/D+Sc+5+XEjRMTWAxMohSF1wWbOAUwOVgxJAiSbEy1UKkgdWTUyZCyNVQJRQICVAwvstd/+HfcO
BlS4Xad+QDLzQoElCbKqFxl6MTPzYAOgRRZKTucUhtdJBGKPv4srWbyse6BiBZdQCX4pp5ysxdyH
PKkOIvs1sc6ZTsg3FZP8x+KdxVePDUL1yiUOvfG97BiDVYlDPP1RxJYnnKyjnCgxJ+lpEivAZXUL
BostNNdMbJ42hZ3jmIlWhVaqOVop5/VgjhY3BQGgLc+rwSsaVSxDuIQsy6+1AgPjv8KylPle/EOe
pS2Yxxtr6KRDDrJSqnNO2cULl1FKWVWmy83Yiy+qcTWLhiy5cnoLF/3Uu+/lJJYw9t3NbSEvqM66
3QOKSK/G+rqeghuRYeGnKbdhUf3CVx44oFVvH6RJ9smZtwYhfRRS2nX5aS+tyxCKrzNWWuNfRlcd
uUirgE67SPMe3oHkIed3QxVwoyzWBa0CmtGvnvxFtYFwaxK9D2FUfLS3+YiP7quwHRP+bayAbjYx
8NZqYgLp25o2ZD+OXN+BI8n0IeK/MiNtBN7T2H+DEKMjftA5a2Kg1ZbYGWE2TBuwplU/OrOxSb/O
0rivODBV0RVl+AnoprdUZ0rja8jIhioJ/vqYkpta8EvzkxRia5nZqfWc5YHIlzmTsKnT0k45tljm
N4ATxP3z+sEKPLcHF/iEriBvApq7Ixpe8i/XlIfOK8C/f3LEq3BuoDk6+9ABD5+m9emBQEI6hIgA
5Ka2gxx/lO6S4TG3eSRPR6Sob/Gylu10LyQ3riOgLCrFUod4MIYZEELlTXHMIQr2xmvCYRK4hTSY
oTjWCVK0DfvbUamGXTuRuBN7TbDidv7ZwIv1tBS3fll/3wM0/HwpL3yHzceINiIwfn0Ow0y2dSf/
fESDIcnh49XPgATn5bHzp9zoQyENdCDehxlf09vCyJiLvciCc1X71GkLDe1fm3nf+VSIoagsNFdR
R5c7GopIvM+o68Amv2VN5zxtzKplGqBmYe9/xQEz93Joz4/4tMnZsOMO4hxAGobdnNpw8p4avPhH
/LrbiWTkhOQIYZSdNZpSxxyEYYToTmH8ZdF9Ovx7wgQobeQyRJlg5nFul6gLrdlPmflpgoISteur
3wsnaMULw3schJCnbtHdRQH7clV4LioZ56zCrD7V14msRn6O55u75R6KJogugYNegidfQGPgNf2u
DUu1YWrISAPn4cff8aKlW/ibopO798xaR3AaJl4hmeHDepa1kd0o7VVtzPixNCSIfQscY/ZLFaVp
gFw7UY8KlRWCqko+SEPtsv4rzlp2dRFnWTgnHJsqFjVCX3bbhkFXcXmBCZWXCqoTv8Pv4Wv1J8GH
OM4rYL/Lywf+wVF6M4nYuv9WdXESV7F6Bu00iuKNtdk540/jVQz+hPkqwRYTSu5QYnzcQp7gRrks
xIFj2WhuY1Wwv7Pv6/oLzvdpYcvWNrALNi/jWD2iIsmmg0cgMwNxLGo2lJPw2pt2QD7zRAxa9yy2
J6ioGUhHyC2iuU6GDJ+3VccDGxzEvlhBMqSz+wKXoGUDrj2w7ICwzGb+W0UeR7j4QT3kgzwUOVzF
Ksm318n3/LoXw59dCRy4qYnpL0ZuGsBqCux+SgbidBi5WeJnStfNWun3E0J6RyGovj2FeojhgaVs
XSQjiupsdzqXUojP0fYrGi4Kan48C7Zmap1PfONePLTgoxYDJhiIpqPHLSQq7/pCdA2E/FjBtsFb
PyrlvJ6Y1376GfSOoWdFjPm//PRs/MAJ9UwCNNjjqzWcbRzJjFlFQpYD9/Kfn8dSuWjwor8Psxkh
zVxlnJz4EGyPgKLytw8nz8yZysDeukRu7JclFjwIPPoYxF6ctKiFjGdeazqhILZSzknXIXIzXJ5x
q9eHzumANrGI3Vr3WrUHx2gsV6xGy4JLBJLXQA9EYtK0hpVPAleGGq1dUdODnlaGHqb+vRrreHh/
kXc7pVc7DZ6QnZPfIfhx7jLEzWSPiL3L4zlCr2A5qTPqF4BUlGPb3j0w2Ojqbw1sFPTxrbDgH4f4
0burPfQk2bcyXX0P6qKNw8yWhH9AEggEpo0uAJug1YNT5S72mv/neDdUqC/NfsCGkk2rvc/KMTjB
7Dawx/D7uakwin1t0/eb1ptjpMT8WbFCdmxCVEvNZzAYWBgkRqeznpDrw30J6f9GDMM+pRSYpT6W
fc9ETxyiQAwRQ6t6ldcycqmLF1xlzxG8F94SaW8wAzVJCMO6S6CQe93jGe2dEZMj7jgmX7OELfwZ
htLID8ovHdJOxUu/PQ6b4iUq1QNSz/RQSmHzoIyxmfytvgd/4zwQrFlLXUrFR9/sEe1uU+tZQFni
NCSJgAGUTWqIq9hD/Pzfjao+AzMOpUA9ypafqYZw54e12zCUth8mApUtIQh2PbrZSj4VBKt26hfI
+EP+vPBvhC0fK6TO2Z70eYfhcKaZdvAvvKdEuJ97YBMJ7jmf0U8KI8n+KVHjcIZQmOeX9AiFzTeb
zC0vunm6JuoXqVweVVKWDNdpUM7X1bH6Rzd1m6cek3vYhJ3bDgi2SLrjYwNICG8F1Ii67kE86dLI
AaAFovp13WsqTDhKl6NoY78A8MalRtV2IFmKBWWz5sG4eVJGHHsp1RKmGRuTcTsJQwkoNWixmHy6
kdlG58642zMaX7opNrUWa7MKc1kH6nFL6a+Tu3oNrm3XCOolXxsf1R7qhsBECDDSITNs1EGMVnxf
Zcce5c5WDSC/oB9PHx+HePH9WPKuQV9uk72mM2la9+QPVvaTDzttkToFWz4P5srPto51Zp9JJ9x6
zxf1pHq53hASArhgQl17JBvAVa2bMGaAeUYYdfCvu2yjh9AC9Nt5GQjNq/VgbNcIN7KxJFZ+xZdU
fSubF6iJEDujwnqjVxa0ab1FPva1kThDrfqzmWWVjmkMV97cBrRzl1BV+Cms4cf8FWtZsNQiv9O2
S+l12vEl33fjDG1jVfgf57PrW+Okm+CAToRFhoy94RHQhn/A/lqp1ckyJIj5iNMxYgTaaUzqknmu
gKobEPFh+2Gw43sn3Ye3PtZgBx//L2FJKwA6WiFd+bZ43fcj/d8FQU5l9yQxt19IallfUHakpkuG
BiCC3TzkvnM01f8n0LtSW9nYOa5Ev7kvcjsEZ6Z1urZk0FYgSEdnI9nzhZuqQKcLjT3DEoPbD4RF
pf/UVJa8ZClVqDTu+lGGfu+dQR4Vv6YzSY9CGXSygKw7WHXGIIdEpc8Mlzltft+0FXrK3WynKSKR
kNR85PUDrzYpF5Rw3TlpBXG1qzOEDigmhwGj/bPW7A4/qSL+fQy1W3S4vkFKhan8ggm5IyYJ6pW1
FLIcMNdviqW1A8qvpTUYhZ5rIRRant2PF/s/UWcpoVl7X/3436spW+VS+AgbP3J06j+VCZMLWdeR
b78QApLbkQ4srJMgStQJjLdIF6qnORpM0Kzu8udFSgg77/bL9JgNdon7TJD33cD9uOVAtNuyqCot
AjRQVt68FYhD+kY7QDZmnJ6KJz7Ic2qtl+K+AL62eltT1HfoxD5lVdBR0oSJFvHFpakcXDlWQA7T
jSiH+aDud/VAJ/DcJFgeVadCljsYLxpc4JCUCgQScD7JdBicwLeRWJmspDMrVCac/NqJ+KcLEpzI
5LNCrMWfyj1GN7gNT3lWn07X8kSVnigmkJe7ZuYR4OYDaOAq4OyMpj+Txxf2Pmv5NL4J4cOlkHCh
OEZPeQElNnI1gn7vUf3bxjPGKHGoKhh/FvKCUYo5VP3eCYTGzo0HCtP0fqtTm1kDpiZfO/7KRXKj
DBp/CpCAZZWUxinXhQ/PBOkW+Mhe9kOT+kmFmoOjzK43Z6JVoVAWHhajnBHllY7Clf4ydg1gPPj2
lNp2q3yYTb8bemK5JUIElXfb5Rxhu51os8gAoBD3PhQfp0/cpTOZ28CTOFsYwVxCvC8inCprYdoZ
8aI2JkPFb7ZHypuAsSSv12zsYboTL2z3oTe0yFnDoOMEScpoN3CNo+r4szcvcNLM/v1qOgYACjpu
j14Zbv4zNl0EcERkmrqE5dUZ4567q6nSEFWMD0FdwphNz10upZo6dSDWPzeRzHTUD3DguNCvnwF3
fCJdUPHfQsp1c1RxA/wNZqfWU6o7QjbivWWzNHfWXmYgAzSKrCtQJ0yWf18BUB9ZdCo+XYfSoqAK
pveO2jvdECUAefXiVLI+x27qGnx4OkU8KQyOhQuqChR8XjAaWOkCUJWw3pkbPXtHsjXBTZ0DB/R5
8Z2oRW6j2SITdocwsHmdU7rN6N49x1vXw+eSKG+TNdq4foNVosIuHQOvo3Vah9uaOExnT0+W8BKn
6RnmpZbVQ/brfZUgT5uVEWeJMaNQW+v5RcJ9StIsoiYSoUI+zYBRdzu8YB2896VHcmnbrKFdIYIl
RD1CAjciB/nCTEmrYTPpMCi8arOmcV+FG3EwylAHoRAaNEleGVOT/DRCTc9Vz0GqZukXc9OAV7bf
AU17vRkx9xTzhPFdRz0BucK7O7CusAQ2OaB5+116BHj9jv8UBjNtA1U/7w2zPazIPF16OPChB54T
rNlCQY9ozGJ7SdI2Ek+cnF082UOl2Qq6LFTKY4Bzz6Ymi9kK5GlqbTOeXgGhJIENoS4V3cc0umiN
kxJtmDXhS4vXr8WLpyVeQU9XGbUmMnxPaMrd+Dojiz2qDIoAVoFO4yvD3LF0vuRiE0ZzcOHPAo29
H3wCAJXVqcCGcJ1w56Dbh8b3SIgZvIyg7uy4Mt6y6vWUJlciB1l/aG2+EDsdtmIAY2glFrq0DXNa
Lhd6Kd+6akgulU3w8O+QSaRFYYMiXRBx5z6Phl6iUqWNCPbMJj4eU0xOaZp35MOrZLHluDoyo/7v
LSKOFvnVpDwC98ISSfXmtMYe1JrHjXbrYcyI5ncxRO3d31J+iDjEewxPJ5UG9cm6i57F0f9vbJli
cXmrcLIWSHFu2AfH6nWNJNjkdLY1c6vacW/yHKQeObZkpaywXbiIY+7/SaEO6M7lywWqJF2AgNz7
oMccEcnt+CNkx2h/tL5Q2/30g37kwANzvFtfenNgL81T3+Cc7n0fk6PhKC9vLFFmgCt3yCABfizt
iaeKthFrOHvBYbwp7CRNR+yuuyXxZb/zTZGhw21CSGejtPG7yI58srnYGqyI6kThjcgWkhMu8U3w
DRbs5Gdq1UcdFaHXQQ/97MC0WhNaaLsKu4Iw3W1eJfPpVzQ9vnmDjLIAYKrKLMRB6E7jm5qdFXC6
47JSOSRujQd/jLab8hHUW23HX/LM4NwcFQapxegWsvun7/js22a/ybPa9tumnooNqUNjAdSyc8Qb
mjcEVYBRtM9Brsy7TkZFKjZF5puA+tf+b4v6GZ9zGzmMvpfqsWiw4RZasYUJvcl0vUaavz2lAcUv
+zfc1nXO/FWgXuc1q9pOTnyi2B9IA8/T8gr6rg5FxvfSBTtuerGRKajZuj9si7Kwc/+S/E4D99OU
oQBSiCULfjyX8926H+2ovFJU5XtzrrZeNdYHbyJp2wLR0co2q6RRDRx04wBciUGf0elRye9pAk6g
oCgQ++BhVYl/RtgdGqs+AznZZivajcoQC3jj1YCKd846ISIhcGZu0TrqFLloL/RtfQ3zpN8ZiTsr
Tq6Tsr4JsCN4vBBe46IiCCreLe8u1JF9LQrUnvcwLTSksi/49Rpf6Ro90nAdhaof46wwcQDM5JB1
rW4VG7/vruLiK2f7WdfEKwkTfkdRpmiSBQW8uspPfbMUKrpsf/gyB9vD3Yj6rvx+/P47J3UGzMXF
9bi3oID3NCVjoph4OkZkXCn0Qcx7HQ1HWcOqm10s02oyui4BA7NAgstUuI0eq/AaBDB6z0YHS2EI
Q/HqzbeTakf4lljoknb4yvLi2PtNRkZjQa13YrxEwm6lytUo99tJP/DdlWXbFo86ymvv74XuiGJg
yFqP7ZqcRIb0vaaYbjg0UKGkXbFOAgd6LYhgTkDYGFZG90QW2aGrpTvEFv1e0+vqQsqmrTi8KQKP
7J5g84KueMUI7/d02NleFRbDwN6jylweqSMAgsqS6+kXZV7YbDTAJNqIvWP3onIFtGOu2dPYMUnc
UElPg6Gr8xP0lXgCjlm9lnt8/F5/bD0y8ujzMKGI7z909Hz+FYZJd/FDoPDa0dQMEK3Y1tlUfrdt
F0gphPCr4N75f7cse5mG8UwrIlxtfQ5QorJoyt3KHlpjj/h/26mLhzJcxLJ16YqDzXIBFjBtGDLY
QAd57YhhBp7Rw3NxAs+vZNGUJXtdHgJTOZV1nvYFRuZaRRmQF9IkOeq9C/uwBQK60Hj6fEYNIUBY
MIdWz7eRAbxBLvmiKJkSTC3WAsYwPR+b1P7CBsekNwBX/YWC2nWl9xhybOZA7kkRqDnBL4Ed12An
MFyLl4oOTtzaeW8cI7zywqOONAApW0nRnjGhvP0xpK5Rv2S44RvSzWQPAiNWT1P0g0b7c1XoP8ae
ENOHoAoTd6Q+RbzMQikbAiqSYMFdTsZBttg0PBci0D4TdC4/nqY1X4PQdtQHCmlNX5wz1+vFpOKn
3RIxxlmjQMYRqizKvwy4JKDmccn0/9ajvdXB8ZKCeswcuIrbVREXmV/YkbYKo2cdUrxsJH8FeO9C
jARw08m5T9KzRwbcvcdDT1U7Xr0N6oJzMpf3tuBOJzhUZI9jG51Dj66dZb3Cu8WrVkVQbMsSkbJK
xohuTc5nmHTYSiu+CRBfhrFJe8rLt9bDexNnMxYzDuk69E3D8UeNx26v8yPVSYTdfgcYw9eoDkRK
6QFIuPzn3bwbX14ZgUwUgUAhNOcpnw9YpxPHniA7IHA6CN+DGIfGU62/mA3QW6k+ZQINwv54q0Wc
U4klstHNK6Zss88YMp9OYW8vCWauMdybG1umJ+eZUYEyRwjCw5viBfkEBrH2kwudngt3+9+QcGrj
z90wuDMSpRwjL7DjMjk0iexa7++nUCjCnrO747OvAwlglZNNB4qzRutpyBBoGm0FIem+P5cJYxVD
TWDzObZCLfH3vwFEJP7/xd20hZ8fshz6iz6r96J9qtrKl/glH3umJlUikjc3y5FC9hVuhrmGMptD
Dnq9yl1Btoj6suI0yDTwNwgJe6uecodYoWQFcOS4Yq4lPMJTz2hKtliH+0oA3HfECqb+RIubndDf
Ijwtaig31+FoveZKGK5Kpw/VQd26mtpu4IHbbyn+b7IXa0J+fo/Z+lFP1v52cuUFNXqXRn/6pmho
H0LgZB0zfUwxP5ca2YiALdSMQKCmanBqgz3FBrUztBK8W+pn+62XnnjYyZOaPF6qoTnAJPHh+moQ
LpMMz5nnNgsxZq97aXGcYzdN+CqZ+wrBCd7p+RkzRRGEzmsfqmMkCefYrkN3fW+ePLBpW5sciaqy
xdF0q08KuevDdZwlg9FSWHAzqAbbvg16Y1ChRCO7VAh+++DPLbZx+VHU/kQ67pveGQIyErD8WTQP
juZ8SfeUECqTTnSEUNN0lX7JlwGbTsvaqqyuQ3I3uyxKanNnDQJ1npmjKeBxJ+W/5BMw6ZAKIqSY
P5SJsnM1oRdyE4glSFkIVqmqN7SozN1Gvk/XQ/6H6Kmj6TiioVWdjnafW9yL/0+fNKUqlNc76Ix6
3K+IuIcC1o6U6MZYNyNWzKefme93WBOLTH8okAsUqi3c/AQAxitzDjUDwvGkaGOQcqpq5OpeuMSc
zNGvlCyVAXpDkvsqjviSSLmRp2ce7snXCFtOjGuNuYopxZb1I57WYUcVLlGbAhsZakzlBFptdEkz
RLkR2ah/vGg8gFJQa7h6mE/8GBVr85NRzjU4PUWox30lp37hrgw4Yz94rR0aE9KA6rVx+ut+QS2U
oS/fhtp42ofM9Ipucc82W4ljRmAzLegCRKUrgXRXFi53QXqInjsJWQEyRV6Zax8bCuJGkGSOE+kO
wMva2tf0dTWaI/rfD+5FoZ9LTZoSJcFpfE6lMzeslZv1ZIVvYJmElCUxdrtkwnzWxEAuywJ04Iqr
sGC4WkAaAej10YBAbFyejQ2cIJiMtXeY74aMO+Ihr4Y+nB2peqZNGc0XXQ/618QGfLFnD6bkRO33
L7ohDl3THvkO8c8s6jyLesqbQx2w4WqGSFCCkwwk7n5RuI0/ikH3m7W3LFELzR2vfBTW5bTJVjVv
FRsBl8c4+KX5KqGOACLPurRLj4gDoU2cg2NODtro3GqarB3aXm9s9px5BkxVzeXB5/WdU3ci7h6W
OetvnJSII5+yQDw+2VWaO7lrzm5L7LrkzJUnHRMRxQg/Fv0rHh5U61q92puBRY/ZfJreaGw78dy3
I8X7cAgEn8XloyPq86LgYBic2G99fSeLcQJzzwWid0/blI14oXZk6BYs24qQUSk9ViNrfAPsSAI1
MHI8W4mj+p4TC1t9m+1s4YGxbODRciYxK584KIzDa0/NyzkfuK0RbdNrqAVc3JZ65cr0qKXtjQHu
F4oHe1NxFI/6geEnbnVEf1+ryJU2sSco//lMxj/MpEUU5Ki6DDhzxLOYkkzHACQ5Djdl0TaGfkjK
xCXHfTY0mH3J+mQ0ajoyd7cxVL6Et19H524SzT1uoQzAyyVX36RFPR0FGguOO9LeEwpX/biIQxLU
zPOPx9dLIJ32wnn9PKUayfjBRMMMzAkLeWWN6W1Lz/xUtGbGCoD8wsOAbOXK40RK66yTAZ9LzGWa
OIuk0ER2glzSizHy87ITUd36KvMBvWp52Mf2Vr0NCvnf7E/n2qSTWDGWSAXOiiR/xLueg3XIIp1b
A4ab/TYtKd0gAFbR1qOK1IMByg7Wu/Yei3pdMzHZjx4Nz7Tc5fOpdYaScMYjct6WERe26QU7Yvuc
VePsmTO3dHh8dgIisfnUVgw6R0m798tJzZn7x4GGGYFiludwVhZ8K1YWOoJB4rUITDy5/z/tI1Ak
NJY8bNd4Ex9mM9XYOUpLgGN75xwAYxgw7u8hdyhsq8v3Lz4PWI4tPrTy/aNduQo+2UlnUtQI4ZCH
7xdijk+kqS0H+loLh8RebyklR6DpJCNKe8HRl/KLuC2naIJmKw1jYfULo24/2o0DimCTxnMqG6Wi
vdBLPbky5o2YxqGLXFSroxN9q1KGTHEtJHdJG7fZTsE73zZ4cdFzp4mVn8kK1Du07QPsgzM092bg
NOLGy3oU+obBdLOuMjj7i4UBW1a1KmpYIxdm9uxf9+00MiKo8FFO+5ttkV/71Dk3SPPPrZw7EDFN
d/4O3KstiN5cqawYxk1v/uxHsmQA024kcbf2tw7jt0PK5bx00Qm6u5kI3KkwWagze8l8m/qJAQM7
txwyL+iepfYk4bj299U1I2RttFDvqDseY3mLpnfLvaGSdTiOlS3dT7OJOZ9s26vfpXdOdoKOBLe1
QL1ubq43oX9PyQTyxxDulrowMSQj2NkZvWK+le7me+mmmMo4LgV0DwS7QoQdHp1mjnJMz8hKWL6u
4+mgZeKf4POAwtle6Ne1fP9dN2ULsChM0mD6jexI5PkOu6YtsSdajmHmr5qz9RkLJ2Fan+WKpkbS
mYj83TTXJ4mM5Z9Oph1A4s4TPYant8/pum461kxJPeA/Zj5I5e4uaY3/lVkTMhrtZrcQradvo+TT
wzdDkx4V0DRWPWkJEIA7VGQbG5NH8KeSmJz4e9+RcWZm+fS/8zwUzRzY0PTxK5TlQTjA79I2kgwo
z0B+5Bi9cRBe3JzQ9xyROd8JuEE0rnVnO00YBKzEJPtoUOnyQMcYROnca56gD3oDK3sgz0kUJ8p2
6/ZRnAFTFI0RRwHY2WRMzNEy5x+QnthRLjK+CU9fCLNg9CbkFp9u+vgXS5xO1428L1xZ2mpf4tFj
mDhfL70pqXEbK78ZYrD7ORVGGUYZAHU8RGN6ZNeXia18yrnW8tdj0/VjgDsT/gypYuCpiuCRafIm
TDiSlYZFUR/lMcDtdv1P14ZjLc688nyAXUi1Je0rZN5Gjmbi8swo9oncavxe6zQNN3soLetrLWVs
bbtnK4GcdB1F1kOvvUCwFDVtyyfZv22kfzak0XnxlKN2dtr5qX3/CvgfK9l15VN6M5vch69iuXjV
YCG6FWWP6y7BQgz6EQJF3atx7wrTVaVuEvFlLY2zdfI8HEaxcwNZGolfif16LewB6G3jd0TCIqa1
TaUxc3RBFRunJNISSGxZIVpBLhBMxLqlkHqODGmUdd0BGjjJ0zjIJ1dkKDhDjGxngLBK1Zqjyqk9
+i/BuICZIXTCt/rL1DU8SSGzF+bENpRJiHZtIt5oludL/gwEpc0A+33pfLozOGT3KbCvatQ42Zh5
N9ps7eC73Kdc1UPzc8ecYSRz9mFwaPDXy8v90Qanuq+EMjDuMuckklNma0zF+/hCgy2idF/N6zfM
eH5kvWum6L/mII3wph4QxU+P50WYlcRtGlDTzx28a1h9z5981Z7fEVSYMBuVNQHfCJJLhdofRZ9S
AIKxiGFKQvOCgjMDkCFojJTS2oU3N9LQuGSX93o6Q5LVmbAdf66JV5YGY4wMIEvSBhEIrK1coMLa
rGuL3yLuv9xhG/Wb6ZvmQ2UmTgAUsmToLh3NvL3btaBS1U2KCZdBPCyJl7FP40mSROzlGjcLOMGl
DiAA4N1JZvahq7l5H4D1sl3nO9c2sJXQ1YqwMdwHpufCYYsgeRM4LcjkiAXsm1T9Xx/SRLEfPS1z
bW9U5R5Rq9Kh6RHekK78G9fHqxfXkhIhYFFPoOWY6jfnXA+BCHvyJxcN2wXOrPligX/hixccp62b
ZK/de8RO/AwfJmERsLOU9T73aChGE/C1wYAJexRThnfYTszIdIUCiso9I3IoTW0LXN2YObqQ3eNP
jsVBFGlOHADOsn0FAheH5awekTd0HUXZfUb7dnOw44X0HK8O7EJ8nVS2mgOycjL2nPIi3RRqhNQt
gOxwlD/zLkRAhwYyzaSBu4h3OnoGz0+P3zukT8KQrdM1Q+BXZWYg5jdQyoavwWhJ3xa6x5gRrFwc
AL0q4g3Ng5KUZnnAEKnWJIhMJc7sN06C60VuwC1nUHSnVbDG1R9njgPMhdAQifRqB1Vx1QXzaoWo
IZiy566fIVFgY/QJX0s/8peAf3dfB8Vw4v/r0CnREzkBWFQU8Fq7XpUzqvr8gCqLV3Y7gTZkUThU
EVHF2WVm6R06vVAbFekW2M5bBEuf+7Hfb0PlRgxupBmYZrruddfs0I2+nxPAdwDYohvXd2LmqJds
EpOqtoxE2soMuHR6zwqE31W249aPJz/eiunvLB2stCnk2Us73YlJycISuMF2uzfr15Exx/kN/9tV
ii82ZqhTcCALPa7xPWxJgIBaa36lxQQzi5i6fz2XTYlkyoOn38TZgL4QdV6Pf1HRPdQSwa6IhJJb
C4B+n4G6KTLPG2+/5Sajqzq5Wen3DIxMGgslvvhN/4nm9zcj+MIbxMQdXdZ8w38ofrqRVwjFvr8Z
EW/0LwX2CdN9N7q4/yOOPnXppYWzfTyG6zpqnuo8twrvyoIkFwHUbC+z17FnHpvSOvESahnZqHDP
x316a0apZS6mVFM1YIsgDJ6RP6Q1ZZ9NapH7lTeK/Hxh2PuKWz5SSzsmn41WYU3Nxj8pIyS581Tr
QebQBGeDalgxmOmOLIlpm9qHNHHmX95wgiExi8pFMWDUOs1Ee5F91xXvkC+NMyNU274Mywit2k4f
YSHGyfocUKnQ/ArcBDNgo/90+bVXpgjgj6YIFB6pqk1b87ERNTJkvibMbZ5J7tcxgTM6KQ++7EtP
K0TA9xAyugp/kRVGTcJzKH0qhYjAejOdZRm0e3R3Z1CYZ4idKRMEdmH7JX7RzjaaXg7D9yo0//3Q
YMs7Jv/cA7JUT0XY9EAVAUQsungSZSU3dDIydk0JbiPchu0mWGAz/+DolPoSlp5/w7x8lskFP0Ln
qneFtwcg44KLkJb2i3d6sSQ9fcepRT+zVqRdgn+0qWfmmBAZ48oQqv/sDCuF2Rj78vuO9u32ZgCY
/rySg6WnQWp6EroT9R6vQSUYvb0p5FOJzbYJvjMrJpkvAsfytvBduDzUTw5HZo8Yex1IIfIY8Ma1
hFK6l3iArYhU52PqB0q+qzqQ7YFK8lnBz07bnCTAIq7wW75dvMi3giC4GfMfbXdB/9lxdZcXTYtW
XMKp6siUoJLV6pf4hsHmuehija32La35NMMwsKirnZEGA8lC1vUyrHwSZiPoaLNYsG40ta3rmrfb
xBX6SWgyFyYrOwBQX/PfluvAgBmKk22DoAI8wfoPYhQOX3SRNmSaB35jgQfSEx7x3WX34dDC7ucF
i2lMJ0tNyqdfHqI4c8NThThNZFoE0ovL02orx4lFvYkQfw9BJj5yLC9Jh+64rpRaQnnLLzLJeNcs
5UnjgbinzFwFB4oPx5lOQRvRgA2mHZZ7IDg4FD3idXPxzQcvm5qYqgQWdpGn6KLbZZy9sdwbXQzF
VRoMzmyLAnk0R0wtP8ULe2/GKMrAVtEslOPTvttfMUqO4FDH00EGGYCc8F5EO6a3R9HNCidkX+jq
2hDfY1NptINlDeygEjEXTzHNj2jdSZUV6VzUCK/wGJMnm3OAtbWqVlT/3zISVCDHKFpsuzwcTJeq
E9BqSZbHADhS1k6kK2xqJHIlTdXq/4Tet3zqY9wqKRLUeZPd5hYjQKwSxRTU+aPrOAnqcQIZ2hl9
Y3yhCWrL/QuAIBsGENMjxs8CqUBwvw0kuADsJKM/82nlc/ucqWo0QRed7h5FwtCUoM5FDnvnbAuO
MjqJsp4QYM1F38IucMH84AAmamop4K/BT1HHh3ewDrl+/S4ViQBmCFnvSJsnTHxT2/AvCACMtYeV
KGpHsPG11jB3l8y9bQl/kHbShK/eBmyU5bqGzfItrkTmu2GYr58g+EIfqmTKqIo0Up+NM9efvyYK
6+hJ3hyqDcMkqlgmRIaymwhiQ1eyIeu8Ic6hqyh/BmO26BglK6lVPzg7VZm/OpJQPPq4ljVY6mvt
tisMoKwqRhnxDYD4oWuhk+zr4xk+6Kidr89Eo587oFBD8Bt29YYrOuR2lzL+GjhqLiP1Bb4E7pH8
P6xOE4Gm9VzluvVVEKFIQDc1mKLjadiEFzIrVToHRsOeqh68x45zVOI8CkpPH4DwFJ0GuvOG/vSL
EYtiCOfUpyp9ufsRtNkgoPhZysfxRiPC4InxWdqIdGYFmFAuVT8/BlzxbKuxD+Uc1Q5/kRJxAoCB
vabGUzsUCWqGQtK5DsiZDbND3bh7p5VSQmXd0k6cryG6UxBiWCdN4D/kVNA4b+om5ipzRENingvv
uqx4Afob8J5fPG5TsePhOIV/I/HH6/0YcwWpjozmA5Zr8n93ApIHALBQeitMh7qxJxFQ/o2bgo2w
MlRY9jb91YO2ksqFd+yaPyk5xS4p9dz5sxiw9WYlDr9AWuoxkaD4SRt+06dP4HvCaP+YYI1deThI
dFPs0JTL2xoKkasCUzGxA29/8McN1X8mTCU3c82yD2cbfsaOBYFg1OTE1ojUf98eIWKDF2ChQdyH
anr0aLDRWsjMKEXO2pSU7FP3ODMr6r2nWtEJIzHBR2Jhy4qKdjQZg2GyCC624UC9Dt1+YDvUOIrU
q42AFeQQ9DNpesfVEjaHYFjz7MBJchopiLVyzKzCIXOtSP4wcDmA11QEX+XMLvbZ+mB/7OT2l2iH
oRsCUDEW6gNK/kdITIf9FMsLK1Kb/39CgS8ZwqmYQDTuWLYNBk6Y8mLx2iZXtsFK08L7w3302htW
b8ePntOUCxpR118GFj+l1vEJzeNAdpQF2/Z09yIk7UAft3lorh/TvimQrbDBo3VnSqeLfEWZtsCy
0mRQxj49NKI2QOjkHfkaNYLVTqNrK7G3qKK0gP6F0WCieXpY3eWTn4tc07QDSU7Z9CPBKgpoD2k5
SWuVa1WRkoC0/TvyJpYlcnAjAAiXhTcPuaS5Uqlx7cfqnBA0YZbedk/mCOQZ/GvYdkjAvpor4D3j
bbIjldzuDdZpSmH27gOJQdgspL79+0RJlPZ/txJhxGqey0OgSOQENU9Y7R8vSGc6wsyXUKpgpE/s
8MS7w54tsvCsjVWCk5uLb93E5R1wy8px9zQpBFBACKRGVf71lUAsNTHe8q3QIJSL00u3LAdvsHHW
Lofg3MU7O+ZV2cqkrWE03CDFxtCtJ9rIB1GQ5RsSfLbSo5JsCeLXAewdsZ2/LbE/KtgraM4QKWkZ
WANy//tOJYGl5tHoqW4AEyD7bbzAqjZsGvy6u/qsxdvrfkDeOg7OHZ4eKFS0bM0iBVFSowntzC2W
Y/y0NGHw8B67dPHXkFVD8HYlJVoyUFMBA3ka3yA6+hLaKt162G3vZFz8nNtPH3/zDZOnJ7p744R1
1i9IllOsFGPjo5lTSxdoUOIZgjQnfW6jNF7PEkymlxUALgku4pZh2+QTSZhFt7ENvLPlWzjmSUXt
sC0uFNEbAXheyYNVVPewt3+k+PMv/+DeBr2VaCh6hJOuOO1ixwvbLn09KORAHVvlGEdKrzg0O/Oa
876eOlJhTAW0sI1d7PaMDExA4fck05LB3JudRaCv4otk1aB/JAwQ1sFrI6aZuOI6fjB7berFXQo8
XPoymYJB9MSvRpCf9xvxbNi19S5XdNl89pO1Qysxmxrm73Mrvi9m0mUQcJl7h92CDVMqseQ/Souv
F5HKA+7VRr+1TeuhGypv5ieOK3DlIZWob6pC24bY1EHkHTW9PPJLfcqw/YJtbBitb4ROAG80Jy01
ZCCBl3hZz79FPr2ZvsXCL+tSoqhlUaDcuIw31OTov37jjuCZK5oC+gqXqZyIzJDdKslM/XVqX+uW
yOMPHNMejLGk10X3iC8YJtqMf3aijxfZPFIK2ed2wk5LWUgxEq7kvnU6uHlXbiJZ+XnQ3ND5Y9AG
ODrae5qJvyv2sSkuZGjkey1tkrUERlpVfbNl+ve6/WfVea5KKI4E9HzS2zBphvWQvgncBtWOLh3/
srvCIRQdtYVRuDbIsNybLe0nORYJdrzWaCqplzltI3idnl4NGJJtRRwpemgFFY9YHDt6NmTkFybu
4w9qgF8TwJiyeY2Q/rfeElNYK7lriXEQ9qzXToLilW9idXy2qD0tHKRtcu7N+UXFItUonhli6KDO
DzAXOYUNXGps30smaTw5BJ+SQbo1G/ugrLGe4TMUfFyjV61nv42c7AkbQ/UjOlsZixpFtQgvNE1+
oeVkL12+pOSiA1+RiQcfnaTHvYHV46rpWGII5lHDGd8YYc3kvOIfLv7XcdVb09NwkiU3WUoKkLh+
qyyc8kmVcUfVggD1PaVfu04J5ia2iQwtNn8o87jGvwt0J0Eof7vPoV6/L8rAWHo8jrqk/0FVRakA
nXYsKl3b7k/wuqN/DiRt22RL6Gjzzx4CaOH7rZr/ql1QT++zpG6O2dMV5tej6Ifmr9u+Amz+9rX1
S5H21sxW0798ICEDYnhP6l1QWRCHXOYNPm2j0uWjuE2OaQgx3ge+s6EDkJn5O8q6bOr+e82KotGW
b6GbI+85fHx0uKPKc78zaEi1mhrDv6Z3r+BsmVCW1bLNM3fj9j6Uv7KLt5TJEaWd1Da11zTuEz6L
ymu53VhfDc8v/Rkxr5Y3eQY6xXh5dvNgiNdF6oF+/9ZLLITewusgcInRSBIdD+PfgqtN6zxRrYR/
Elaf8Ps75JvCaIbPngVODXqDxS3S/zXykZ6u/seza1xCAon/gQARfLD8tMwkJ/7SnlinOSUl0a4t
96a3sIZ3UyZlBvGjPwmmNE5WMFMxg/SuAgPSf39WaRkslcQwXwc1jif/bmtvJjfIGo+TEdSLJSWS
BHIgXETyB6/XeKjzMiIa1AlzeU71Yy50Z0AZ0wJFXBKqu2qVt+i7dIFmV9pCWw+3/+Ayp0sn/Jyp
k6S6DlEcXdNZ/dMC6qlk+mVTOoZr0BHJmKYdlU1bxPZlr5kJTxxXe50fSboGqQwh6Lc+EEK8HvkE
fK0Mt+UlnWupY1YqeB+AehrcL6SY2/gc300fE27BXyJRPQ1HgehLLTObPIhMHnzGccW83xP0b0tZ
vmY+Xb9tP4i/9rJYeHtKvIsPCyz4WkZlCJTrcua1jZwop8VDi30mZ9C4z9vY0gDL30azFztG84iQ
m7vlPdQwlso2miCIWqg7w8Z+fWTZ8BAb/HVW60E1VbW9x7rAXySYPRcV5Qha6pGnVzkjtmtCkPgW
OBDe6k0glr37xuHsWiuB2UnBf/XNKu8Zvq1juM+Eo0QCo8Yo+tleEWZREuEkU9RkaG1ZtbFrGbhC
hzxt7I+SaemDtLGajCn1mPUtXIJsiGclB9z4/eZg2JsYGOFV/wWI60IqSOLd8U1TyKmtvOGmgiOX
7JDKq/YzJ3btGrtmglYRXaCB+K9pIZ3WJy5vb5WuYRaXwaCRVkH7B3N+q0I4BsCk9lRHYsMNhgsX
rm1JJKlrovPAGYATQO3bpIPisOXUVBXc/Vn4MmtF6TrDUYXIVuKk6Pe+J9E2vdijf1IxaYip97eS
GbylTf4+W1V3LDtuoo0utkF1LehxlkTtA5tIo9q9SSsQSyDHufjqeay91p97rTRdIic66C96q8qR
JuOB3dYisWdp7NqAOqokPSk/SM1aZaP32TaqliBghrwHSXN2/pT/k5s12E4HmjsiaGLp+z5s2ZqZ
HAeAgGnl3kwFeqNythgZ1r6h+7OxBBxZELg2VMcEYCIbjKulTuBJryY3EHt18u1p9xAl3oLjBoLw
oehNnkuy0RrEUYZFp8EAfhlUmkTzGJ+3r/aZo3GKZWYmSmkOs1SMJaAkHcDKrV8ZchxDrERmVzxq
anFAT2bnEti0h/6z2RZdey6HXG6r+zgbNEjhDU5sKQVNclreIUMHZKOarMkYzuh97i8xK3L0mbyy
6+BpkBoHjqHep0w2t6qQTjuMig0i2GdxC2KIi+sIj9e+8Op0bKOi1cCi3oDJjsRoIXTaZn0A25HN
EdSJwEwghSR/7hnNNI5y/bw51tI5l9isMN4gNp7dxnUfJq9DETbq+EBmWDDwTx1ivM+WyStUGX67
qnw2HR+Jbf/kZ3+a+x+WHSDX18Ew0otnl4bklG/Of8CQhd6tn12hhEII2VKA74gad+sIZ6FvYpSK
2Pt+2H18kz2t6WR4PDVoRVd/bCL0WSIn3Gn5EQMPRPemc1kr9AigooVAvi5aKeyGBGDIm7BGGiMc
OIM6Cc25WAm9rcw6X9+xTt6TBFJDJidXC5d5TaK7sf3VGctd1t28AT9mZ58IhjjW/p2SE/FTCrRk
3q1x+1x7N9M3aTmh6A8l5J6XrShmk4Rv1lzqIgG6BT9pXikIiD1bGuHq56l39gALeBhfkaZD0LZP
afykCmfudlbh/VxQXM+idkRbGcZb6ADEuuqkzfMoinA/j4uEBJorOPscz27q6IYfMMSV58RDF/qb
2YpquMvnJ23jlwsDk0Ua7iDxTP3WelLjS936hBOha5/b7WdfzVy0J6xiGWQenkQajn47IS6+I//w
imaQ1wI1pfSBmspCDVENw9x0EA+sv4V7gNRCCbqPj3E/76eErod4NcrzAgANWIGxQCLn6Yl3tCrx
wbuBO0RH8g1l2mO6rEj1vna3Mjzvb5GWn9oGerjmRsJz7hp3NvwnaCXzF+dk/hsFnNyr82ErBMS6
fJxJKBPJ3zWn5wOvGUPyHDPbo+b95CVQ2UVw9YRtADUjy7ws278QfkuVMRyo9GPCigWh0fs5iJMz
YkLZM8ZycQZyV2B0UxxG8WWceYEV08VoeREt6e+3b6IWtJjd75Ut9Cy35u0VKsRHb0S490XzXy2y
W6zIDy5Ol+E8vF2po8BTReEgEmNt90RwrAzagjCqS6fsHT2UMJ5O9w/5K/8bI6bRoJYbV7tfNpqM
hcF/JkuvpDy+DWAOX4JZOSfA8WP4yqtzmccOWzEfwvGG0Go67fuwbU7L9pb2PVAHCFuI1sib3/EY
shYijCm0MpbMhBhtWEKItNMf5R5bQTU4+pdqxAiEP8dJCIRHGCyR8vgG2fgKe/fpIze19Dvn6nj/
t0qV+FMaC2A4DiYnryDFik5BxMSCjMCq1JPgSTYL4V5IszT14kYRmjgGfuRvaKUhQc82xT2YWm1W
KM0WMt11DdtLrPu9OPwBBcM4Om9/4KlBJgW6XCSLLV+0MY8FADjzQf/Hh3fCYLeYRrjRWOMS6iDP
S5s4MvfNbeQJznzSfkj/IrpC97xgEI9qL2Uskn4vHGiCoMdzOc2GaasySos/bHJyqQkD3+cwCcBn
P0Yx5OdmqSdvvekT4oLVnoxsMrzLty8qqB3ZpViZD1cNnSTpycB8/h2wg+6bItOJhGmps27gJS8H
1vcb4dInKllWz7uc/0o1YzpDPoa3qV6JYqT6FP7vXKgUjEWG60ym0OtIETXWcDYPqacWav1ehyjf
N4hOkNX1vMYb8gr1hJfksW66mawJgo/+zTuLaTLkDT0VO5un+tGqfn2loBnM8V2htxfnKkJng/jA
SI8VdsUl4TT2KDxwh9sXTGC0dIGQpRRs2DB7217gk/kC82tw38FlDHQQW4Ko56auFcI5j/mM8sKf
W+xIjuunQZC46XfrCQMoInvcwWB4d2b/g7eOemmQmWeoWXGa72FlxztEXcYFqTWCzUszRMjws9li
OAlUb0n9pJFxBus2suYqlNJ1scmYsJXI3FSKeiBJuTuSn8CNY73GhtlxetPOPhmZ7fG293pI5/KZ
t2fEg++vIttgMP48URrKmsfXssn+NCAuylWuz3/QcvSxTav2LRgAryJt0NyzJrNlRzTq4yWJKOxM
2ElSGR8n7BvI+Ohy9wL+JELI8rEQhnCb6hL+D8v9RvrM3xd+6nq9D9+IbFBt2tX5gwig+QM4NLrX
935+ngINBqoKRDBbxEcyRiQJ8QbzA/G0SMnMPTOrHLbEndf6KXTJkBLpE4EtySHY1MqBvVsLVLQ3
uGhpapL1qRmSBuaOYPUx4D1mjD8Xjirb23xQspmuDqHg+lB4AkHvUrNAwvv1xBuahw4Ct4nB6XRj
7m3G/DiOENU/WMTZe+glvlEW0JHqLO11Zm2+1pQAjgvBD8cjigK2sKDg6b3ChMZMl5yVmjx80+D/
2ALTIPk7oNHY/0i5EjqNCFhN+9w/u8HXWROFvq+jU6TZiZAYhYz8xYeu4n86UnHG63il4Dzda28S
NaQlXQX8kT5tBCnwCItp4IWlCd3Srk6OC4sb2rAJiovKlOPyHLnPytay28ogp+9O9r2JomfReNXX
7CfYqAEz6j5psoemmzpw5AFlAxm22sboGHum9N5Y2HN8inznU45J4b6wSjZc7AxxUmEwokuIpITf
tT4rRl99HO7UpiN7l0zL3lAZCQDPN2PH2GmU78YZJQex3CNDtT67RitMim3xG62R1c+EmyLTiB4D
6PvVe/Q6lOYNYKcuWcgcMfi38unasgCKw4TxhNqgJSc+0ql06hDygsA107fQxpGDjeOd3LWI/T/p
qBEglSF5XD8tuoXkmSg6AFXJ6bhF1FEa9uuD0lCcdnFY1gHzFb1q7R9nizNKLi6ItMKRIhQuJLVo
/O1+aEvEvAjWnmyHNSAjNT5Kb8evycfQtAzbgMZx4oiiTewV6WouITD5JxbeEhpukHgVUyh/mYRK
vljhOeC8rU8yZUqxcJ8C9dInDfLgHikJxg68iBFsrTpaRfgYqRCocFR7RPTHyGKrHxLbplhOMEfw
mfKGMVhd6E8W+K/L0JwcNQxgb/YOxIZPcNWFR7207xo1KtcmYzM4D/sviX5K1ouDFu/FpHQrWJ9T
AmaB6PXacprZLsYOTGJxw+4u2vDvwbQbQNIU91gWktyNLZJNA0q9i7ujf1Cl/m6h4nJVCGpzn4kg
8np1oota0GHvn1WTYcnX5P69aSpttKtABzVhO2S19V/weu7ut61NVUUU8fxliC4jot67Vw8qk8qi
gD4ODKqkcHc8p7lc1RESFOc5PRpFvGZBSS8L3neHX1BWeyBmH8vQrd8hgy7uTgOhf9vKV/Xi5mEK
CZ5g7njCKgALqH4yYqOHxbFE+7b6rMgIAHgoqXxgrBovw3XdW6HYDU5T0+HCcg07y92ucpiCEHgk
ohh2JlI9fQf6ZEwu9z/0vpYZ4NHlBD3riAkHpJWrg3gOEa661/YnMfRfVqB1zCwmuxjkVlA/YDgm
1fpDcgOU3MoOg2ZyAoPPQORCfyoM9woV+HTCVK7wCELfL1/mGhx16nvW5rMRtd90ZjVEuL0zlxA+
EEwwYoT3vp+qMv6D3RQJfUC+RAIgLZ1y1xFrW85Nvt02ERk5nTqiZx5CfwPvCglgDXnICU/dv0mS
TnVycGqu7cYVywX6/bgO70KAl4Qt/55zxv6aucpcAYQydg7EZLNqwoFR1rs7hXfKxdhA/NpT/IFd
SmzKn7TPmAsmke7Kc8DxvxXsXdO87w7oIkWK8a2XpaF45ver31j90+zzS28gCVRGfEg0K0Y6h/nn
8dweKNBZX2ChldgQ1f1/2sBIrxNPKV/9K7ScI9a9isdU588SuDJyglJJqNztlLP1FDrx7hEnXXt7
8T39nRkztRbzq/TaKWiWTL9r19hwtAhDfRN9kZ/Re6RPZcA1x9XVF3eNvP15FGwbueLBHoqlR2uL
oemr+49x7ck8+8HRFuYZV6wb3Z/kQu6cbdyOBbQth9zVBxxvKIM0RfLV03uRcFipy28YXL3WEIpM
d03UGET+YQhIIyDOE5Emr1tzF/oPKq7eIr3ty/QyRWQ2yMZURXNZyfbLmmRn8J/siSpQ7NrCRZvR
GZMPhNIqfJD/zqupYpQ0AdO+unnsGQwVkjKUmyqQiPFca1Yakg80HnGbz1wSZEe+UXHrJwjvnQRO
lKJpYa9ci6uc0dyL6pkUdujFlRiBRzasvPyvh/2Acu5/uVNaKWDNa82igS30AK1DxTeI6hEYzNYg
v8/llAtYs4Xhz4t9JtOXmEBjma2xSzvyuAI/Jz6o25Az0FenxvmU6xrGUQfmOH5DphBZeoD8dwIC
Al3NrLKoJmdTF86ZwEs63tDexsO4vaZ/dD5HX6mxPb3kMjEF3lHbR8pV2j03kckysBS7o2dQoVUK
hx51cPkk8+Fck2ARWjU2nCBVYfdwvrsAfXR8XsgIyi228TkygEV0bOopGU3w3EXsy8mvN04Xbi4R
5ge8Ab66CfTVnKWLPRrBWbVR0Z8e/+zoUzQt/cTn8CfdABReIARIEFCafdMtKo79v5/EQzyc96nM
BD4wNMyN81O+RHhkgbwjIdZqfTlyIJ8KpIhroNUkFqL6gwSLt0xUJ+d5iqZnOZR6OH684hd22+VE
EWiNCLWmZTcogduh38iH22jLB342h0nEIcdnm2cdzw6fSFDRNW31tc26SgAQMn7uzD2RmYPCgDqf
tNm7ilnxjJdKMzfJtjQz/gCOQXgNTfYx81iIS4U99a6FTUTFfrNkV855AI9TnOabWNzSCb2p010m
K0eyV8khjRegNSRCdUjCWk2NR/zcD2UvC0xr1VVvUMU6fjdWzrNLG2RFTkrVbZwHOs5QBYZEFhdU
u4rMJz7WHuA+jv5UM/swwxWWY66V5FztI83SMJVUqA50xFWfbecfCeRx97fHLiV3oyMkugmd6LP6
MhVDPsDCBcREBCGik68LMJocVFuh+Pya10ftlffk0vnwlmQKXmIQ5kG2Cr8nVvUm+D/h62HFYBM1
L0773O4u0FYFWyvPzQKHqQJ9xyVXZDZFTT8S+cNkFoDhMXyF1uk5RqZVPbnXgyNw3aGoVLRpJBVR
KZsQw1mqgEmIzRalzjQ+9aKQrmcwhlqgRUaFYG0tMVT8//2s0enPGXWMk3NmV/Edti6hO1ttgZO8
bYeVFp5c2SL9UBLgUTChVz+i672t3wuDB6c9Ds8ShuTTGgf3mb57hPOETHHqLboXOuCKHF+UugdI
an7W6Ynac+LdE4/4ymn6IPS08oUMdKBkH+DDOGISgoc/lyUEYN46f7oWShbfcatlmZSoVv1V00AC
fq2mULjumeKy77kpurrVJf5jHL05/134FQC2z59c0aUEQEhHE+lnnpsCQqhNTa+CUZbHDfCGDqo8
BHK8LqGWL6PNWIhfRKoOlaMDlpgWlP6aGeoUmexmAZVzGl78cc6HZ/2Dgpk5qq0a5jv7oBr8RQph
0yzYqzNyws7NNhibW+skFhpkOQMY9pClIHFpz0UjrZwJnxRx7028O6dIXd9Ry3BLZ8YimeSMQN5y
LkCScLeSlwEei32KgqKlREDc1D5sMl7FkHeLZsw8Qd51MSy0Qsi+DmD+zds96afCGByfCcGmsVfT
8jB00tbB3oouOeLe3DeEgb1/+G+uOMU1R/i4q9eaEe4+yA+L0FdlN4zastwYGTMdSW6vGurIyHxs
yAW0N1mVg3QttDskTy64Lcts1lYXEZSzbohyCwzkWO8jwDg1sOu1F0TLPkmmZdcKj36EE7ykLbGS
ydjgHnrM9cNLe4SV4GrMp2XpFiI1MyN3zhswOvr3eVnO6I+UJcMvtfRCe3aTVnU3JMmAVF/Kbvj5
O/VQ1h7sLHz8HPxhZCF9uBXppnY5zZ0/v8vfxIsmshcDJZaMk7XtPUIGag/VhxjuNDPL82MQXtYy
JvSAGklN6OadPWkEQJw7JHNPxfd7KMjQaWChm/Js9MJupXm8kn8vIFd15EQhpZVAOhjyBrvPYfC2
k8heNVCJfDudJ2cKkcXDM7AVBYQn1zmho+rOIcPw1I/XlI2Qj5ckYNkxtwL9VI/9f+pA7oepsS2p
5lrnpGgwCOfl0XOFIholZawmpm3M/82577TpY5QSoVpC6S7k1GCXFW4gjv21Fm4QKlOBon64mDwk
QeaeSnmzwPYeKMXTTk1/dFw2H8p5LzZk3WEMWrmKQkOUQGVdn5FQKZ3RnE60RJmlGIW17OaaAAxc
0vWIYvf2qTc0pgqK/J+/KKR5upoMfgmPYOJupnu3z+o0I2tsNv+dBwNbkCn5sLjH37z/pvWELpXa
Md9yrnmHOXIA0RHCHGeABJ6L2wHWmvPdeqIYclFKGH0zVBTOivGT7dyBaPgW9UnT4y0SoBC80IyJ
yOQXA7bY29O36YStE3LhLvSa3CZxcFPFhc7I01Tymm860JW2v3c8k2lobYnqha2ECN7onhbDLCYN
lj1Oh8LRdjyZ5j6M0PSkcXfTCaGvt58ZOGDAabOeJKHEIDN27enmhy/uSRY+I1MhG+Fw/6TsPS0B
sHPWUU6AoCUWjZtuQwVOtDypE1okMXGhm4WSDaGzQRcFQI/aAfHH3u9PNh3TuT9nt7fetameLXMW
/bEuGa0t+EYbWa0LPmeHlvPDlUALolXdfRa/7tdoVs6NAzoHmDjlQMu7VWyLff5zNJF3SJ1bb5vj
Csw/HXgkrDJjJTYcsYFeB0SixjG3mLQA6mU20iR6298wbDd6hBfVEWybN2zO0t40teNf/P5HsZ/C
Vnk9fj8nZhD9K7jc5GKlIXHBYXo6v+U3mVJ3cIRg4kHsKuPThnySZQLFVdaMORBzd/63XisBzWXn
gsqJr0k1wUmS0it1sDR1Q1hQvRbS5Ehkk4rGB9rnQuaXrAS97qOeijB2UiNRu5JOGcbG1979lfW2
OXwDqI1ghAOarqr6MItHmniTz8GI6Y+TQcfi3Sc/NWxKOeaeh5GHJUjGvbqJ1auDXuPJSRKMmskO
hwtT6w1eN5RiaI5/Hr9B32pirmviE/hRwztvPW4jHTejG3vrcnRjkyt/5H2SHhKH6kO9bL1u1Xxf
nc30w/M8/EkIiZY/oNfti4v/BLIaItymHUPxWhyTlJzHuGEmlfH2p/HetZuLp3PbM4fHShm3dCC/
JD47nJa6XgaRrkxe49ItCtJueSwAevHnRLUTc2hln1eUMDw7csPdmRB9Iyt7h1lzFUUfTx1xiQoF
q1XR1BYDFrnKatmIpteQxuZWCcSI5fcRRsyvoktjfGPmGiib80KHIAfBY+8VB1O68foMd+HK6olt
1zXOSShVbsekuY5l0d18H30YC2O7DpSm4P4A0mMcKr7XReGnJmIXlCVPPaItJZV4aUnb2M33JYVR
U8YQdqSmirgnHXPc+Pq7jjZTLLjoWUU2V5ix1ezvHEcjF8nIeLUTaezFWE70mabxHzrLd/ZjlFgQ
QWiqAx1Udk+6L16b1AJ01/Jj5a5jVCfGPwR1ZRxl79/dFuu6K4yyrMlRjGw8eJRl9kwzD5KbhuEH
ie9gpSUbOXsq/nvYHnMC7yhH/V+6VWlvsGSRY1FmziIClzgWHfRQvy5NuXtrHgehQ7/XZi9/eBqP
Ff/skubfy5j8vPIcVS1/NbDuJkxMdXquprXIJ5B0GD5+E+KrZ9tmghn+iIIYNPK6vRzz1+FRjhwb
VNtIRJaNFFTEBvnx1OoSforMTAnvZy0uZ+xmiwC+skfzwnwOxyXGd2WhgJwcPJHXd2GKDvde1HTx
fmWbGF4fZntPFW2GvgbULSGUrrmvAs1vJaA7sMwJwpbxeAlNeX9d6E8WBM1OC/kFapEt+f9cI2B1
c8bWBWZfN2kgwTuliSq32ET6FPedU8aqSVRwIA0AgfM6Py1zvddUoFaMf2wML3VzfXRoRx5Eo23+
iPjKHCUnUEfiYWZ6W121MS3sdFCGYnYnCRPcT6SDgu8uvdfTo31oQP+KQWjdkn8xV+44rsayP8OB
gnzmv0fwgyqxzrvqYAtxn6p7TQdxg2dLoJ3xfeCTeq+3DQNg3JHOjwX8Dvg4GHJF/zJQUZrlYYhJ
k+ouLTxRfbXYbY6edu/w8VKNTpv+HRHM+5RZyZbMxr1I9V/cv704ZTYeREDQVcAINMDH5KXT3iRg
bBbd7ELCAGznKre2h/fQItE7deoYyd+0U3hWFnGB+lqNKhjZwBqSgnmqQYnHZAcV+KfGAPAIhdVu
WXaqBb5ld51wlvNWSDSQ8lEkpriC6iHu+jlN4mq4YuqFLFlg9pav2lf/VbypQYsCH2XC+3ixrx1e
UHeUHjptxeVPAQkVDxFXiu2n/3nLfw5cwufMvBYy3QLpeUrJpE7HhKyQPqsef0bB2SJ3ZLUUCMD0
fDSujHwRKFtZcHQHH5NqT1fzSC2izvXcZj46x+zyGkAe1Y9onhffWE0VCzTKaWxLKlccvhjoSQGa
9he7Gsh5N9NVgC3DZxRvclEULogNewF+W0g+NaeEes4NYrxdloaMU/b+ghJE2p1amMAc9z7tfm/u
EKFjhm5qfoVh/5WyWhfwJLsnyBAWCipBJIpveVBtbNp9LY2x8cF+n3MwJcLXaFolqyfx0x2LVsOP
31VG65F8VP/sbPuLfLRRs1Hh5n/QTzkj4tQaIy+SsgMfxWq4r5yq8G5qBoB2GwXnvl8zemMnAE4v
VZG0CuJ2fn2R5JE9Bt+I6ndes2zZ9ddiceH3NohIqCjzo7nZTLXUJeLt3PUZNaJ8vEYtC/BXaYLS
5IK7Ikf2b+2SC+cAzM08a+q5hyau/6m/GJEWW5lk25gafB4WtwKaW4WEspIeNDrRM14uoaS2koRi
5dYOxGYlMA4aDU9EjU8yN4M7S+0U0ZK73myXJTez1mPbXl2JSVl4m+jDxBR0H9iB6Ca3LGOEFO+3
J4ofMSPaQlPBUYdFQ+ZerhT2aV0V4zia4XalBc/dzcflb6Tqp7/Li82kDL0TKOgUSoCbVhnNGG3R
IiR9zSx+56GCmYYeg+GIb1h+BIioHzpXr7+pMXW8Bby9BykqQ/DPc1AeIJRQn9oeTmD1jyOKO1ZT
0RlurDtnSbXzI5bGKu3ktENyqWNaQTm00ONgShfJmTIPBbwfVcK8c9InFxkTnccb5IbBIKOVPbUo
sytkgbppWEh6HfhVb4t1Ij46gcA904VvmEVa/FSXlHlz0Etxjme90cA5qAlJZ/efUhDqlFNCVwSI
OoGTwAigw240CirphWU17uUeZGFJMriuCsCKqi/3SI0sr0vQGrcK+kBi5KVdLuA5mmflgX4CF1+u
TSncSrzS2ZpUmZtL4t6R//V7NnGDlJq8aOagg4Vr7dwaGUekEm7+9eRWaExPAEfKM3uZYgcspKo/
g2Q3pqxqSYOl84Xn2+Jp5VO5NRLJhlG99XAZz2OJqovyefPGrDOBPppI/t7O2JsAV+r8B52kgG2b
QLAOjC1te0+9eZ+v8g+kJkMbN+S+FbZmnu6ivBoBG2zBu6zU78mDpiyD9tmtJ8tAxx9nZ4X6vaPc
t6pcN8/inDHvU6O1mprM1jNawymBiRKknc8lLwAkJ5hTqyTKDffKE4dbTzAMQ4Y+FycS8Owv0WO6
jCLA24yEeh79F1Hx2JApAUyS73HQAxXOtpLIJyCt5UFmTwyYO9+/EEdHjJM5yofDiGHAm0XdZEMF
J5g0Blqhd8L2OSYoyFuVi+IQh0AuZzrLV+qT8YBR6YLXjvEKTo2Wvk6mu80qV0xOJ7Q7WvgFJOF0
J/hIvp7Qzre/wAG5ZcSbQpsQHeglJf1ej50pwzhH2N1PPEa3BPWsU5ci31KyyxPcSx4vCHeMfkpH
NuFk7ebZ7c4ASq2EJ5Y3X5dq11aB6c2ecU/FLmIoPtKl7p7vgfnEFL1SV5yf9C3CeIYwXPRyOEhu
yZUPUV6luj3sJ/0a0EN4VcZcj77tog9+FCDmJ+vAvsFtlzF0eZnN8aM77t1IUMx6Eb7zaNay2wpA
CyRzD39mEIo0kEH+7H/agGneLcxBYUXI1eJdTFBOu2hSS8qTGUQoCv9dpCbN64tq4Ym9d7nRwv1f
LtDuahd03RBQkYucrJlZTiekkQ9y92hPKii8AX1h/IWmT8muJBH7lLULrKdVt2HA7LcX+rVwUD73
YY2dbcbyF1FW9MiCKbBiYuJ92f0lY4kPu0iFiGwk91nshgM/l8Onu7kaVCyzmhuVV5pHeKVIB6FA
GYh5CLrpO3VpAllNhyo+A8KFLFtVNIl0WlMjP00HondCd58VlaG8fBkcaxH2lG0Xm0cN41V91xBA
5M3z6JlEXv5GN3YVEBtXGPcjnR1IG4t8NS0gqR9PVzNRcYoAwrCjgNZW17aPOLbuOl6VnHB1sPTs
BZaQU3uvjmi3RV7OWPzZ7koPLbbfb45Q42udN6hyl+cPNoxJSbeQ11KJSkjyG1MP0PWv9bs2PTUg
uruvMX3vwr0BOOS+SSqT8+b+Igbd+pXZVaH/lFf8Vs5+XFxH3IwRG1b5k+zzhL+PZt/zGiojrywa
RUje7BdT6iQYjkkCx4Hbm4DjE64W8VLFPx/BpwwO2hQorNHgiQOziDDdv76gUlC+8u8fKhwJyFAD
joP3xxoIF/7jZtER7wpPUWly/8opxm/2pmclQW/+m0v4golHmCQ/lFQMiJhEVJwIAicr9cyVMXaz
I6HVBgqvUVKwGTujS9/ihJdn8jDK91fN5FVbyV7kHydqVxNMT1xvlb1shKgzawbIrW8n4kgI7lt/
DFaeYO8OK2tgISEHpJYfSegpNgs85EyfzOAaRXvgOIyeTbCWIIIzLvyfF2zbzrc6LzfHNQYgQ17o
WBRgH2X6CY/3OCvCAoANmUhssbMZkd0ptQrtUiNH1iLZ3MKCjaJWxXfIHp6+gHu9x9uDNttZMKpW
uTh7cqM7Ap1VSXFV77+nCUSGUxSUzaoeYuZK13LTjxZ5OR1glrR2cTfwIWA/r0kLkW1iU57V92B0
HwQ5j0MYbDku3+QBw5aoRlSGBPJoiie8AIIR8MVJGzpsmLJKUmHARwNHyHxv0e093f94oWEbqn2m
jt5025aylwX0cC4yyHcsl0EB5vCIX80A7ZgkiwQvPfIezHM+8S4KYnk83+dGIZlxuKfTvDJfTm7T
S44WgAC11ABeu7Ws8zpU7kftLKAV5tZzaPYqi/4DGtA1hxHPBbSpSwl1LftqdogFPBOMLMUrdSMf
AmKOA29YBN4NUXf7loF+NjAzUVYEpW3tiIP6DrwGT0dyJRWUzkeAAg8GA5MpLCo/CWlnXe/GW1E3
dER9KLrBWIOyBwlctp6ad4FWwXg0LwNLoONCqNXgA5gkYO0mqvHySSM5htMmId18TtKaXQXfQQr1
hfhcqkzjb2JIdrsJ6WrkUHcbta/EoH5FqFLb3Pm53pDi5idLsOvgLuErajL7qoVuqPJTlO0OKgTE
itkgKbgcGIARNu5osxs4SbIgh9/TJG2rMJFc5QRdjKhp4T/hRxULgV0CwQeVUe5YHTstQQHfq3Hr
a3zXFVqnWW/jQDtcvFcp4gl6rQFWDzEGou+PLhi3mm638tv4B2FQi9iRlwkgONvHcG1qI++zp91e
WsCtnXQ9T0iVRO5WfK93PeSRG9Joep1RyTEf/Hqe7sUSxaE53f66OuLnZIjwKpY1eOHPkorPsoEl
/qSdV7eTZ6hdE9IdMQ8+6qasfa7kCQfGAhr+r7oRta9WPksmYe+K+uLY1MV7eUYI6d2gbFGACrbi
i2KnkvNm0ZE50avJNufc+jfD3fLLAMNzVotKoJCAARRxyRpIvv8X3oLSGcaQyQLUqrUN2Goatztx
Qx1grkRv5fHjg6SwMH/He5g6lHg2KI2PrehrPYUpRbLaaA80H9Mcz+oh5CpfIvsq6kcPMGn80UTW
XjnEqjKLGKaDIryUDAnoaLG+XJlWhQ4D7pk5JQSwyuNg0aY4C9vWW91xPtH3/5I41y1YvMe2TtsF
A6Kbkq3J5rjRdZ4CHbHGZ+nheFFnFh0O8vZIeEhLSnD7KcKfaZvpxps36pxdoYx9DXzXcSKtFWkB
RKe+Rjov6ADgdQ2ewhxS0XJ5np4MaGLo8y5dumlGQOEv/kehs6F68pstzIFnwIGrFVr9SL9+8R+0
b9+G+x8vDkzvQ5n+bNS8TH1J4STUoaJ0aZTIbR3VprboTTTaMXPEHWUBwC26YdGD3kMOrz5tFvte
Vta6PGaaYY2uXPP4bX+Z3Z9VW9VPZmu4NLIuqOiZ/Aw/KcxTTjk/3qPtKcjrMcJiB5o3xJDGXLtG
tcSDnJjpJwtAG1WBGooIxnTTpHS1Kx9R4v2T5SU0o8+RfKosvPl2ywJM/3zXLhYNd2K3u2z/Mum7
AKiOuJecaqdLMIUQ4c0t+JdzDTERZ28TVaEHDfOp0AyLXvwYl2gO30IAy4s/fRsuzrBBrsl4gfNq
D0Bh4Wf8WGZdpdTidFNKNcnW0f3XFLR1Morn+c1LOqOWOjKAR/cf3uxKyUisqUo0rCArYVpk+Gjo
PWAUQzrV242+zy/sVKXTisKMzeBrymzV4h9mcGUIW/Qzy+qgtqaOHVEIMOgV/rYfPcfzdDL8O/Sg
0k4PaJ+GWxjvHTRj1ghWrLS+Jv9Rri/UQC44/OHvLCRk07GeWZAKnzeknW4nDFsL8jKyzfcom8ap
tvAy3ZXnUw6qG+WeHdmJVwZARGu60FbRUDfTbWRJbXsvhSO6ajeFQy6/CrghtSyfp0raq8RBLtEv
Hu1UNt916SgZTAwFyQC7LhbiDIkuAGC4i/kMg3TLm/2ctOJbV3E8wUgVMhign2KNlgNYq3dkNxUX
xb5c4AbJX/5mtdi3bvvRD+2qiTg2vyM1KXsbrblw3HoBs0Cr86XKtj6ZXv7g2z0NpgWC1zCK+wGd
sDm4Wc8k7Q8eODGH1R1wP2eqU6LmxSB0UvMZp5fVGe0/8+EeZNYWN+/BOLorDHFJpXRvHYDiVqvs
CZEIGcZKkHx8J05r74D49oBqVzE7xoOjNrGhANAiVARIf+tKItOE/iIMzSxryE2ipAH95x1KSnpt
3+1/fRGT31MM1EJRC5VLAmjI+or8vcsu2E/pgXgQmEAJVJLnoJTu1ZnEJbRG8x3Qg4XSs0od6Ne7
AHWYZHK+IVrOLH0SZEzTuuuYIBq1tR0mRXGrth6q2rCRmya2VqMyF2JEph4w3Vp8QJRNIyx2Ttq6
rhfFNvMmP0gaKscpxoPXLH/Jwz0kjuCj8S4TZ5gR5otbF3W+G18vFb8ap0kXrOZtJF6qi9RxWojG
osLIX3mmmSutUznF2zGFRbaqhrahGWhgusB9lTo4lsUmkvOlL69m6mVn6tdSqw+rhc3oHToTLG5f
2ltaNH6E6aVMqRXAWwnntosmGH7OyGgcsgH/VdImdhOYABRpQrp45NusnE4MUro/R6QzUNgkXY/L
8AgOLKqp28PiylTJdIZ0LBuUyYWbXOmytbsRUCEUMaKC8ZwecU99rpNpcUJbFNR5AECRt4lCy7rc
rGtQHVQXL92lErqcIZvAb/wiLKxz4Jj2w5IALDm0U4JT7ZyMF5V5DzumAzGh6HVchilMjwhTRBg4
uj4vxdTdajJA7yjG2wslqJQWeqbNawGmF55mTt45TZ1WNKMLnjsiQN+b6uRnsn0+D+lbwQlrpaVM
CVAdNmFXgFy/j3eV7dqUTAcpaLmcrD08ESE2rkIVCSUsRcl5eGYP6nHrlr3qQv02kvXDz4SJlglr
smnFY0eAjUoyMEkvRBvYo9tXq6pVRJvHruldFoq+bRil2fV2MZE7vvdIHAa5gIt6fW02Ezcpofu1
SxwrHDdjt4SU5rfwmdtmZygZrVpNY2Zt/bLkdH6z84SG236MqF8MCPkLNC/a+Hu7T21wA1XqdVwu
UN6IwF6lEvYL7jIsIQ9VcoXO4LlhD5A2d2lZhwhCWChuaZBpiHTsa4TLCIZRLHVbnvTxFDMjZVk6
w5BZlXuT3/cudPXJeXjutiJEAtgo2HB46ErIZL2Li4rjfdK3zrF0yuagy7V0fMgYWJNlvhWowyI+
jm2KbwWDBvrpwStCFPzoKdEJbLt/yU09jBAunZ8KKYlYMa38AN8ISyjrA+MzsVbqqSXjkJbr24Qh
hNmTstc+30FdorLZHcZ/2C4aCfYGC3Qd4YehJEw/v2y7U5Ad490UT1wmdDeQ6WF59qaVQFwU7QX9
XiHL4NafuTEjUsGZ7dFSRGB7ZOFVCUvs3o9jz1/idN+K9UcZwhRCkJC9YTEuFHdM7VGu2mOLbDKS
35e3LSbSeuqcZcSZyrES0HI5RuB2l777qy6IQYbJHu33BJ/5+861AB2IRlQC803UV3GBxhuTbytw
dai2jV1TLMolOoSYFv7AFQf0kqUZvm7VfNNptnwo6aOqjtxn/H3KyIf0DZwZ3lTKfi53KERKqdpJ
xSQE2TMPvdzFEUG7lfWKbptnEpZ6aUOpQ8Yl+aflW4yGvQpVw5KeVDbC4ZwS1X1KGyOVDPOJCv3F
PEe5vwvc93ibnOgtiWafMZ0/kHhZNdYZcE25xbx0LWOyCi+9PbN+Ctxd1lW+SfBSG+4yk9WSa1q4
78/o1/20eKtJewi8d/z4smAiP1d+WHfO6qj4OKUbrF7QkA/rWY0LVY09Aycm7fLDlcEy33yxgXpj
G5+5HqkSu/pMGe8AagfOctImOVlOaCcyFvv8UO+eWrknZMZ51S8wPpDmI0AmdvuZdnHHyYSKOov6
gJssew+Eb3XYtJp1TmQMwCqk2eZcKLbQWpi8HJNXNBIfWBXkUu/DzbbeLwH3nkGjYbv3wtk222RY
L7wBrF3JZ4Hzbp+tsd142tn59TDXntcBBA4u2IyhE+hGAOCV6OahEKZC1NfRZkn//8Cm/gpo3J14
kITUVwCzBQksykasKPKKgVju4yVMoJOtPVf65I8QJrg2Gqk/SpokM3Az/Q4M6YnhbmSEg4jzjMpk
B8xNmJCWnbF//zKaeyyLSyUeHEHstsl46XH4oBaK1KZS7/kx5yYbQa8qukzgZQ+HJh+R5QgZzrli
kKP9BnoxLS4p7tLqz/0EHwb6L7kR7GPdC5E7q3Sl+ufwj/YMAUhnPBCvHW85DDiSzwrxUDGxVIRC
vQtx4hHtGjjO8wXnyevJr7txFWdMGJ0TXGhChMC2V7MT+ZLWMqwm7BwwC2eZfoawXujSIcC5ePWY
kNvF0pGWsfJiHlELiC+wnJ+m3lvY7Sc/t9b2x84I1Cj0o3EA4pibDTZCUWSU14jFMCY5TtQBknfI
iRs82W8ePQqOdt/MhY3AQPfD6bfVamYz4jio+B5kATWeUW7Vf9ShlsSGmxzMcmBrChSs4U4OUcHB
oVZQ1KlnlZknhS0nBmd6LTMR1Gjh2tANiYwlGTqgBlvb13Ch9F+4gtlXs0eEJi8dgq6S69r9MfEV
/rCfF/KmMnoQ7/G2Lscvy5pl75JoffJeDiErzNGBhZeDB8jD3wApZ7+6ijbX0gECQZ2EVisdJvNe
Arb/2TYXLpekhMC3Zyqo2irpqkd2jhND5w+wVgrftcILee1IZmoGEkA+gxfR0Fi0FGSHYa5wJDh3
3xPZmkqoSLKnYbzxngmf+6FmDCBueIkJEbC1EsuFaWKlZUw+ZzzpZIG2IzkMmAZDfP39A6p83cG/
Wk2N5KkpH4hKNdUDrOzqZsmK5boIz4O0kCHYvlQ5Oet/DHeeaNOz4bX/qlJnBWxrUG1Hfkf1Z6sD
2c29FdCzS5KZZZ7B6E1djRuISaPGN+NAnUKod3Zs3tvioiuzrv4JvSnzntsSeK1T7D1FMivOfQRM
kazM8/ct43Ps699f4K0n4iy8+tzwumNN6gq2LefcCYDB651PXPFujQJ2GM5hrFyIHAbyPoUDzkdA
TW2PIOOP8wq/N2UqfdIviKeIMVWAACc0R5GYlAvB90kk2UzZ0oeC+VMskpXEMJaazcsCE3jCfMR0
43sU4KbMSjpCg9XSNNBZCMNDADT21QLxqCQEWdW+NFnbdjnt6YodTkbRx1IrBBtHSiT+8x+agscz
puhR5Conz749rRZYd7zueSfFEOmgBJUuAkVOdsqQvVwIqZ6q3cUW5m/6eoffWxzl1aaWL8/wmH9g
oKNT6IBPIBPpwdg3q/KzyOhji6G9YcK6gr5NF7EMtdBaI4jT2INAHThDxZMhf3ar20fsCtfrG7nJ
OMjeSLDiDbhlwykWEQEtTZI3wThPBsWjt4Gd7hcbnlIUdnZN77bP9oZ3uXHAFkLhFqiHklLotx7/
xWzR7AY5G4vpnK+PYLa37cu7x3vylst1za01ep2RvbdriqV7rAgI4Gclcigik7etuwU/yUCt3XFm
wksNDZ0KgndT+c2dsBobAWrTB1TT907693lE7bGDYjcoxL1gvZ2JVC9IoxwL22slNH/UZleYYP7l
9gYaJ+aaQch3gOoLMHsc8Iv7vcYpeHuexIVAh0VKBSNLyuZzAIpuG0NSqBgBe2XwrIYkk9WWwBWh
mxxcHzSeugyETPNQy25OJJFKJXUY9bumwnNKZZFo6zQeKe22e5qAxgDvsC9pAHDkyGchlm0meO1G
gPmXLBkdfbLZNmNzcV4YvGHwU2rUy9FYjHcaCBkKgxakIq7mOf9eD1hE3pJJdZ72q/DQwcF7rE57
723G6Pu2jDUOHiKHv7Dxmt6Pt6ew/7rPS1pFfOIVvsrtkn0sAl+N7zWb9qx6C+2aJeIoHhKD+uc8
HXzHn17KmQNx2CL4xaxlKWrHg6Rk7y/cq4XfJUIavhben0dvHSXf3SF8Aa7aYTbDHNNG4wNIdA+9
EEtWCKjcZJmgFe7DwtYbDG6Ycq3mFacfHxfxh7mK2EK8LymPykL/3Q4oZ9XdW5F6racnmT0K70/w
suCpBWPhquD7omgnx9VAaGB2ZXt6jU67VqW8+dZi4Aejnhela7mp73YBPXVox/H2JDdXJ8x+Oyom
3rOsnhfcqSzH/beButu4dRywma5GJG8hz3I+QEZRDCq7U/VzxzJbvhHJs8I2NDk0cAqJqjJSRsUI
oBAv1gAnBMO9vgrGpzwIz/DQ0IDlCbsJQPV8Uet8/qXoyBtIT1C8S2yhzo3pZokakEOeZ7h/umhB
W7nartMoOguw1yj6dql66Qm7Dr2KG7MK1nPXCRHi6w1IFiReR2KbjX/dAAeH+msnhm2K3U4SO7L4
8qjvKgp7Gkcj930cg6+7GC6ea6frdQKlfNxFh10c8Fmju15Mc4KnLAeqfgOfUxXMNmRDI8UYV9SA
HDqPBc2hPjn5m3g+ZmzThNRcevYqtbbELqqVfhjMakZN9ysHx2dU50SmYcKYOqMRZeyPAg2Nqvf2
JYQjiBs6UtymnvpFuZIZAPlU0AM02YkCRkb+91VnUsvEckJiylM/QIuG12o8yWfXe8F3qTiXeWNn
Gf0X6FxLPSfK6TNnJX8deQO58uR+C6Eph6kKYTHL7mCC/FwxrEPcM6sMwTgEHCIcCPhTSknspLop
+9MqMOYKJ++c9t2bfeVl6huhRwqdBH4A3SIeKhbyBkrKOuR+ncdT3sP+iYbpZjReM5DzLL20YKjy
BLH0d/3gxE76BHAPEpMyiAa7Cde/UuPWHiErAscm7oYBRlTKNOqXo1lxZWIdn+DbWIHUMImRNNuv
hUYn571j+XTev5q1YFE1SpuhfXI3uw0G8w06NxraAfACtS1lxcD6P+uNtBWM/081nC+rFd0TTg/7
4j+50pEWAKe4jHoRwYP+couu47qCVBjl6vSumcsQIh72QNhcLweP6SZ8/Q+uRxECl+d1+ZL+x/Dl
OQv1l8ocJZbXlilgZNlArbe6tR+gxYVaAFHhQl8hbMKnxbQXAE4cbjhvpO/Njrm4NpaqCrXMlYn9
tTLnxGZmCf86Cr50LvVj6NN0to3C8AHVA/0vT40sX4J0KRJNjh6w0DP3YHPuERxRlXOwHzmrp2+7
caog3CzG1s53ltd26tiQyygvNjEdF2UuYH9QTTUvJbeWoB155ZciqIb37I+97l3zoj8xSK4McSzS
jfSTvEuWApNvEedUMNhQMh2iWloiEAh7Ay7G8WgmeX0Nosp9WMtPPt6RYxe1ofrHbcLtH+bHjrW6
yDD9Uw+FxTUnlm4/40l9pcPdUiWzygo+LiYrQSy+QD7VIHELkD+pgQTpR52bM2BxB3jYmFxuoRpl
GxFJv/6PBcxIMjAJQK/ANUY/McTm9lJAIzZ+OTQ2+goTPuELz3wY82fs8ZgEFk9k0g9SSAVspSHK
iqkaJ2qce5bFaxpb/MvXevBIvH+TO+ooPzz3GEElazQgVIg3kuzvJ1m38UZVoUzvtTvq4xl44d/+
0z3MCZnNQGKGfa+hzge//LvtLBF9HiUlJ9C2Miq+LOFY+uoxJNgfK5/jjsFEi4Ur0kx4NmK7v0C9
i5XTNcarpIAvcw+KYLHNTKBqM312mx9bSstH+1JLwRab7knPIlW3d4hdsWRkb/6tdy8eZlfJhNoD
ChwM8work7zvKAvOtOTPYmEK4W25Nt7kvsfd6anioz3Aq9vvWNiSpP7vm3CM6vQzW9zp+tx/ufqe
SDyzYxVZhuq1cpkLkUuobR86D+YJqFxVjEz7vNco3VPzquX6IfkISG1SUThCuXQizB5nzKAUrZWl
QsD2A7VlCio0foNY1dnZXgpuvb8IrJFsQyV44HFuYd/HBpWc2FXGwEMoILur8L3YX3SAQ59nSbff
K6Fvo/OdOldsKSb+ZIZIFZa4kBWPWHIwiHBgXo4Uj4H6XKgm58LbjMb2K+1cpsVw0+2e4JeyOZ0z
50EA7BSZ2dCB8faiZqvEdzKwvK67i6yRbOm2HovlUPSDNU3BsRPi7m2xe/B/7ahG6ZSeQUD5kT+D
onmqNGOtjNprIpCqqO8FeId9SGDe0abtwXhphA6z89VKphue/rbfH7Hor4ODHrf2WOrwKe1Nxu0F
jlXAN2+4RYoIYRdbYuM/Chznw2qIH1UmA6jcS6sRdbiwPUxRSYB2a3XpovPzzPSX26K6NZc0SMQw
P26CR+sLfV5z40sliJgkceNHcnjalWMsYJeZGQ0QC67Kpn8DA65ABMqSEHAvnJAiY7EaqHPFaVxE
6BsSvhOQgRT9C6RH51Qi4z9K5XPolT1uexL6eD9afsLq3hMN0HvKyGpx1qa73pj754pmULZSFAfR
dMXISbMnS9GF2Y4KzG1sxtyLk0vpynKGxrGZHcuOk1FydOwn/3KFw9/GEPxllIkESue9jsiKzPvn
siXlweQmfyh7nqQY/tKRUtz4IzJgLzV8qTitI1St+JFLGWLdNXqO5wCokqYq94ztwAty6sVJrE22
H4wEsW8Se+49toBRN0Hjmjihoofh2Y7JqFEsxKNYRAXTz2Xf3u+kxscn/T80NrpgHl0X+Fb+V5gA
F26i+aIQmYzCO+PUWGOTUwuy75KSvl8Hc1r9WcGK2oMikx+S94KYPMBxWVjOkiHaldVLTUboDlxS
EndJfKF1csQyBuVuLyPsEdPUEekZPd3Kl5ZW/9yTSdK+HvDh9qzSZWEn0OwbNJcDJ3PGjFAa/8tK
o0VpqWK/1zpQQvF33cAmgzP3WLEddCBAmkGDx6qzRUaPD22nXLJcHLIiUwe1vLcZIhssD20H3vdH
cANzkvVCoSuVgEATugiOZXF7ab3ubOztQHkwHLYYmqwjeTaZvinRwxXGPSEu75z3qVQyeNMIo9IA
KZVzHH5WH5l1cEYwvkw2ElrLDbC/3A0qzXpYzjybJ4qtIRVAbBP78kVNoE/IQa6U3rQNLW29TL63
HcVdKz1kmfwsB+SZBbrAfc9BPcTgY7RhUUCKRcD6kynjdaVUu3R+8GAXTwh0tZ4QRJCmWMyDqY+J
fL2j5NOyKULWi8ThDasffcSncvlGTSXDZ6s4d3JeQd/GMyxUmIU6DhDg7TBRJQ7EOCZLNpHtjCzh
cuuWxY/PgSUfkP1q07KGh9NSHY93lPZ2RfI0omM3e7EK/lEzLKCvxdVJoE/LHpNjYMVfxFAVsaGA
CRmXoPu0G7VI/AghXeE8n9o5EGyQNkeYWS2DQS6+AN4tEVfQY/HIJ5afrCSzZ1oN2H7FikyNExFr
PCcq6kuhWgcSbfwHf9tEdwiN5Q1+t0P0MbEEj6dR18PinKQ9hqOyYky24aIcHqMfoljN1o9HNXbZ
D8tXwlABVlJ3kW6dXD8KY5kRLFa0Ut6123WwlJohWZJJ+49agriexfOFsFJ9Obh3+P6ST3lGlvvW
KWN1p1b7hNsbZizm/sVHFUzeYyqhbyHqpxNEhjc7cQBGJW/lmpzDqPc6B1DL0DPJ72ZXOMOA00et
lRUCIhtQ/lCeB/NKNuHEzh0qp2l0W993kdUl3HAD+jDeGGBxzC6PmvhDaQwSDLSzPP3/SzMazyIi
/g/0aod2n/cQEdDLqm800P6cjgYVYjL1PNrx1DOIkqccRoxTl87T608LAFGg4YaNPkVwrjSDMTT8
5hebBhYcjjPKe/7j29mQnn62j+V2ANIApoX86k/nRXBZVjpIJzo+H0Q7Vl1cL9WyGu2bGEfYN+wA
2ftOdtAeMOSErWtJ5IXQBYAYEBlqNrZLPmF7Q5c6zw+juo5n9/Q8UfQX+s7w1GZZ6vNjNA2L5RZB
ImhNOrg45T84oJYZjD0K1i4P8IvGG4wsuDDnMVTaGU0FT3fohvX8WqlNMGi3qV/1TCFF9qpAzwPF
OEOanbjAfXTZnol73pIod/QeVjh+chm8CgqeNua3q5b4ZREJTrrCSR19ALB08Bq/blgbfZoI263u
J6dKwgUX4FKX+A/+RYpk8g5i8XWLfGkmrFNYOqDegegshQQTe7YnTiLow7dWUkektPhcGS0SK1A+
24oRUYWYncA61zL7WJgKJZQjjBqYwtwtk7MHTVZNSVNv4AJRhLMBv2gB1zGxWlHcNw0xf4xMZmas
TPFhRzP4oysyH0brvRl+zd/tOOLL4hw02l9lJFHsT1+LPRSVhDrwLv9lzTjJziQKycfEaY+dy7EN
tBv26x8TuOAfjcAXXiiQGrXZSXF0Vjovpdn+qS+0iWdRjFWyK9Q/K6vU/y/039W/EFSBS3sqGBU3
JwchkWu4N25z1UkWi9dgQJGbLbI3GX0Jx/FQZn+P8XcAzX3tIXDDkdoCFoi3Sv/IEWq4n1CvAJq3
VgeaKwOWQ0TtVQ6muhrxlvl50jLEwMkxg/JhBIbtgbm+1FnkH2WSsXFiYIP7rJzxSGrnsxhfkqBf
Q+8liGeK/tnG7Z6FhMzG00AWvrRtnHnY79eQr1PSa3u9tuixec1SYyVHTRQorHv+HkH/jLes9Dyb
V8SS5F/vghhYLj620zzjI25FzCmfIeailM10GYPFetD6Iu6qaZrebigYnyADu8Fu1ZuMc6vlIwmR
FhB5pOEYXU5cL5+L9K+FwF+qZpxYaJaUn7sp0Mc3YDwkDoY8O5ne5GU880mEq/YHO8aAIiFyuyMl
/Oh5H8ctPwiNh8E8/8bh8TmuF27solzIxCRbxAtlmo2qTNHYMtZEqgZ07UZfkI5WZIWS7aZje3ep
rRjm8KCKUsvofI+B3Z8HRKAk/lKGURNOTsrpFgPPnKzaZHyvXmNqW475cQZsuGIsW6d0+37nZ7RR
EF2J7ssQxjbp3ffBhD5qfLqI908cIcUhtMVIcluz00EbbMdQFM0XB1rc21lEb0OUziplRkyKGx6f
dx275rLIG9EyVYRatzWkVHe/q+n5DoJzEdZGldZ9NCwJUZqK4Wa6GLi50FpcksAfLtOQeOXg/4rn
aADFsyRcL/KBPVtfvmgP856ummTO84MaTe3vNmK8Ga2unSrtn2QnjBoPKAUv087hdBATZSKPzYiW
vaeR/lPnHCie1qvo2GWlqplcYmM0+zO++KdoX0+es3NctHzoHfHPd88nUD2Ja3l1Ax/c0syk0Lt4
ukhXJWAf+F/EIHPDxNlfyWi8gEBu9ZfbmXzpR+06x+Jr8q9kkFJ82I1A3Pjyn6NVPbad0mYzS4rD
soCr5pnQgkP5A+gg+EP7w36vOmMZIvZFqM2emPVEIxwZQgCHvE0LXWHhZsVf/LeqJlIaJVTgDuAJ
ZLPX0FyNQ41N5Gl2XRom3HJVHFZysXhEQGVZ1i2zlzGbtuIEW1KjSVzu7F330LQAb00V3Il0El4D
cmvoz9I8Q8/+NuBE2MgbYwX+IucJY9wI7BTp1xTn+W0L9AUn7jDQjL2UngOaRv3OIxj1b6gY0oI6
K5eie8vLATsWsih4BUOaHWlsNOnoBDShBorZfVa17sGoaMx4shn2pKQiNVd0QS/BuWmqGKXVcjJv
2tLTOS48F5j3hDd+qQ69GzXrOaacZCMo47McYrbmRqt1gnU3Z5h8yEjz0TrykwvYsy7oRCyIvLt9
Bw+f4sWaHurne82vZSb5ztmWHDHG+nRKQ8yDmNLJdxiHplJ8z7/uWtK2zsiCWBJP6tsKf7sdoXwy
FId/Uswu11SHXlVB9WRJlwuHkfVW4zRCEW7Ufnm0OC9FcP3WXe79VOKmOvx9RLrPvmsyGPwocc96
pyO1hHmYaIwL2gYkcrOK3ovs3hKiET9W8WiN6rRJnNiZX09zyR3cDOmmMd7j4v62xT2fMIMj/oiF
GUh8BEbORceI8AErf/ADHt0ozgrhikMoorb3AMdqr+RJJW2GpQfmzW2WGIEcEBk6sysz1dm5Gz0i
xpJlwCn1FTNDXuxe0V9UzxcFAfQSVZzU1TECIhvFAcWW8l2mtL/S5dKyuBUg3EaKPQBvlEBkR8kZ
OncFdSs3N8reEJxIB4VDjO8xkoRYlXMiiWBPuin4V5Pv7LWOYFtr5sYCEYu1tdi78f6bYaLLaoTR
Qt2yBxkj9ag8v9eMOog7QJ9dbdJgjYrVIZfddoE7D1LMxbhshI7STNmIe8wrlLVlHUnqkoUT/Ayf
fCWa+9Hhz+Y/YliCVyOybKKCyqu5VWz6M6XeIbXEYDypTOIjuNUex9K9gNlKJ71MErNH2nALo4HU
4y8gINHmawpLprh8eZMdZGax5nXz7Y/hHqBa8PVDVL+hLzJpo+0V8wEq/Mz3G4HmGJEsq3RBapxF
MFxo14ozphFzUV/mW6pDjYQV1ySMSami8rHUuQVwszfrw7MT3U2UE2oNwxL2IM4aVYrskhO7j3vx
ddr+MY0DHzY8CTWxQF6GfN7Qjr7YQbEMzS9ZWK4biu9XCLFWVty6EdExULH84xBWYT8aPhLVl97p
YPjI3rP+WuOahChnWxre8S+AT9p/nNi6nIyAlgx8xD+g+8LI6KTZW6wNfJY5lBnGQDxh04p87N5f
pC/My7ebn35G7e3HtUgDuQFl2vaBYKiP2EktGh9PVvFmCf8RV450ZZOd0qV8SveCL9h6Nn3YchXv
CUn5nKMghtPDcz0KHFwFGKWKJJV/FzED5WQFb2TtqwJ2i8a92hlA9gA8nmCi+alGy+8zTHY8Tr97
ZmnCOpM1ufhypg8OrEuZOO9TQ+zyz6IfWeWuqI3LmzsLEoi1fh9J1IwFREF+HS+p9HQymbhKMs4f
oF8/QOpzKvRtO8sHij4te4vPPbOATdzl/EQ5RmWoaC1DUjcSnQyVEvpBrtlaztxezKjEA0sQjL01
DXl6UemViwyZvQmyXu4GaRWAqEvcVRrcF61JLOgziH/CN2muC8n5ryvk33Mt88fhUJ4OsALhcxp0
I5aPgkndGS9rypztDaNaLqTm+TI9SxCshNNWwUu9zcYvVY+iGn2p5kIh014CvF5uqUMb5XFDTrJ2
PyKk8CFxkYeHp00mTKmkkHsWpQx7c9iKcr2ULa88lySda5XuPU+HnPf3ztoMQzmrRz4Y12Sycex5
RP6LZa0fFsAR/YZ/4IgU8O89gCYT8R0rzo130rHJYmcMZPKWoPutd6Oj+hcyj56FUbe6ko5PjeRX
yzgr2tZTUxB4Cuh39ItgXDU+vy4rRKnVqbtzOhrl3rr540HiTVXb2qx1Cqlj3A2NBKWNjNY6jL1I
bdP9vMjtv/ELoJXYc5zKotFEWBy2ALpzDxtC7X+RSWofR9neaK3VP78cgAbW5cxIdi2QM78ch7TQ
DxR7W37aXb8Tnjh/tlBXJNduZ0MOP6OFgmAoFY14+qBZCWJinVqb/6h0wGfuJ/QT7KhRoAiUqIy1
LCTeMB8zxJZM1J2XHbSPt5dYboTaXT2XxDfHXrXVsEfguCQ+NN0xAMXgpjzX0ABhKV5v1jebPzXm
W4nx7DV8F9IYsv7T9+wlufko8NIRzmgqbgoTEo5+I8l34UfQFMgkhMbdoKiYFhPeblApFjbWwYuq
8EzfTaw/Svs/aPJREfG/PkIdQsHTInU2zhMpRC0jhjudSAjHOa4vrNta655LfmN3NwbUiH4NaEVh
2P9JHun337GyEEvIw9Cgg/kb9vnRbYcGnFprABHH8DPe3GBVuhyxaUHOoXorqickHlNHjVkOsGl2
IakZ3iQjnKTAFYlEZBvBvy+zd+WeEA5BtUE4APLRRMiOjyL54EIc21xdq865WkKlHvYLV9Id9i4u
pkodIh2yGvU7gp/8QSe+1ttvceRz4CBTudptf632eV6w+V9bSf1n1LMIgUkX0umXYPYBgiyi30zM
mLV6kmpTyK982AcxAzcOi6OmaZsGvIR5wwx3rlfWCIxZcs+DTGXN+HRXvpMfqhYubOUlXh+51tOL
YzQL7k31qo3XZJEcjvOB3IM1THosdCu6KQlDp/Gp7O10OktguzzkJ1KJmMa1vXKydQkUozLfYPU1
LiZw/57xNHiYNdx3RB+HkkmaP6XcnHbBm1Sds6zgHiMUed5IRrDtV1q1WjUxNJQdgNedauA8lYPc
HEY3NafciecBo1/MybMexdFmYA3AJa8DhKc2AgTgQok/QRGjwzgZL1pz3sWFRWx7LyyMeAkVstVg
L/blYhO+MK8Gy3Fd9GtfsQrdEySTpqAnYC+FlFHEiBfgpSjURRsdvwhCbXuOsTon/2tqhnbgG2gf
naXOe3Tmv5BsyN14oKXRpCWu9p/UOrdeeVIk1zJT0hxSo79gJ84errLtx/61igfcczhRQSKNnruB
07nqIK1EWc3IkWjibDKfGSxmpBplrevJZH10cxtGNmmja7vmbbY+/efmeGL/WcNbDq2wlLZDncxl
6GNyLoPjwIU1MYETauQ9qkCDfUybLNXGDY9rQMfyGaoDIbicOhi1lYIu9acjSfjayRm0AKT2Jzye
mf0apJPXCc5nY/CYWx1I14JVI6XnddUm07ileSgqgXlwxGl8DoIxapPs7XdnxFwd9airPOtYqBR2
mUPaxUMtM7WMli7hGQmBodLHS/SoMvd04slqCEcMEfsp1+GbayyEPJV2GeCp0hbxFYNKXG0lZgD4
hFQyWkYyk6ovZ2Au5FRXMKGqDf08Zm/TtjRUOv9kc3HyA2dZQHndXJPCsVuJPsXMulM1EHbdHueB
U7+Lg9JSpHIK6ncB7Idi2shYESuUiiBxwyJpKM+xCD769fEYzeCwIFYQLF/8A4AQyriY7pfA9Wc2
bG26p+fcoM7vQHut1qmQVNrfQuGwfIkqvNHRlteoYFB7prSc+hZq0zRPVCYIYlBFWhdzQfDfDiP6
0lq2Z/fcqddrO5qBPUvNUhEEGZ0OLqqhfTX0d2Hns1YTJ0EDOTr7oPPNZsvVOmK+brIayyB9Ahc+
0v6mh1FO342el1y8YrgS+gsgJ9Vm+i+gEyePhKwVYgy2L5c/wVCwe/zM9O/CqGy6ZVv5w7npummP
9u99nozerRGNk+92yrwmZNA1JfvwtmvdoqIDOMjoGFcBOeFigtrRtUGCPb3kQEWFJw0K0iXUTeiY
2cW+E3ZnaqnbxXzDtar1P6fHuXj44Qz6gPsV8DTNpE4QrRpjhssOftTMdqe199TVFOAvgCQ4hdDm
kWrRgQ5+taG8P1FOkF2NOhe+pCw3LWM7sQbatGwon9oZ73yMrfysL4rIwg8XgYpIW5/1yeRr5XRa
O65QzjvQL2+YPPRDrYVw4HXC2cg3Oh3436Xk5upsWrMETMny34t6mKyYdoWEWUa/eQbdprk32NqB
PXJ41qNME1go+yMY58qO9PWNZt2oclkpZ8tVtHdS7OuNOEAVoHsL5FwjbsKixTIr/y/uzQlAzhfM
pJjblFiudM+Lqu+LOFjicg3YnRiZwWdRFpQ9Eu1PsJVGsUblIkQ18MSG3MvOH5upOZzBpSDLwj6I
yY/weGMwKkUmx9fHROrh3cn+OCgqbY0BagGjQUC6o/GfCusUij1srgaM0BUyco57RGvl54sxA7pT
nVzNbVXQbUs3yW0CQLrOMZt4qFYOudNTryA483BezpsG4BtNnon7TnnRlaZn/Mt5yTNUv3pdTGS3
DdDpdBUjgvgKcKEBXicwr/OsAnctgEw7CVqrHv57BhS7CQwdDa9cbV56kI2MZ3pXkp6XLVJicyYn
rcMOGu9ENJGvmbTvGJ5K+xnBwT9lsJ5O+jfbm1TFNErxm6dgNDmwES5DIoXbLBHBQ5F1mABV/23a
G3jMC3eIjvKUqcChw2g0tvPJgEqqLh65yzKbItTOFofh9qE0y3ajHvb3UDR5IIcFnE9u+gnZGv/G
pJ7YWZ22Ltc80rKVoi0PSqoXGm4Mj91v+8wwpT3tnBKFmTiBb71ZDgRH0/zXN+cGfniNbm6T0xSx
ZcE4xOtjwf7PvFAKgE6galfYVLbF5ugzpnlxQRiDLTs8uPT7rKV3eTYQ1gA9mjxzdrsSZ/UV+qOa
TTdaQibWrixyuTAPPJqsGuFzu+fT/e3L6gZDnVzBRMX1pmZJV5HNCze9B+jwp+tshjYVFCEezztu
zPIPshWd3s7FKUoMrXylkYPysH9CkT5kYPDrFj0xZt7Bt9WuXeiUzvQ9/jwRa1e2qvZkzOP3AuH2
2zu6Xj7lsSz90fKKplcz+9Px6qhZyUFL1ZOsiujJBAZm8ncwUg/tYmSPPDhcomCDR7s+WX7OWjBt
pMYD67ePAYrgMV77cz+qFoLA2/GMDy5nje2e8qbspPxen+pg7R0fR+ccpzGuKymZh3rBANNZX4eW
jkERTofbij6BUAjGtKOX8B5ssxf7RlJuo/nUtJs1OVH9ijcS08+trpDwrI7um8B5H9bHzoYfqqzq
6tE5OhYDs2dlP/uOCQuuTx+Obh260aqhkJB1Ta83JBMGNIO6yJf+Pm7ZFLKQL8OqvWVXoQa6cqj9
qhCd5/dHZtmLbwES7Rb5CSWJtfoe9lRjN/tCJfhAG1knTY/cbTYgQwmo/BT61bA8YNOlpZZk/S5o
zngLct8LSYKrmIdWELbEstioXh9Otpx56qDXtLLTlBwouGQxNQ5C4kbAf3Eg1obYZaxJUcLmV8Ih
64KyHINcQnsLmABq8UnTkvVEQ2d1zzdJUB+dL4zhaR32pyQ4l6v3gsSkiyAjHrHepkOOkSZszSzp
NzOUxO41fyupik1wctAt3lXJVXiLACFwW+PLolzjyuCF5Oz8MO1Th0AfnK+sQKn3q5KkOLMMta5g
DZ+BaikEmKnXmXXg1tOM/KhhwJQGPj35PjoAqBO4BdNT7k9fvh8ZpJFxG1MzFSPE2qpAaw5h+G4j
PmXKwZXqrkGSHTVhO3QpzMCCVAgQmdYPRCCj45b8iyjtRKyOXBlzDPhCzV6bcAf+9393jTwkuNVW
eed8HfUv4K9zCbfCGC8cvhYvJ3qufyMhM5+uU9oFRtO/QKmtN4iJY42MSgEllXjPnekKvOK3w35d
sE6NmLDuGgSCpZr/hIdeWlVVnEQPcerVE4MxMuFMFx10+WiQWtBzcRzv1KwhmYLYSJiMOwS9TQCl
kcjzF/LzC8eIWYUja2qjAhfbLWgf0HYSUG7NR96SUO+Emp96hLuu4ohlPG120zXr+Iy1kUySgupJ
PouRK12qOJvqr3ul/mAwQcbWBxhyYZn0I9/eBOo2yYUlbHFSbwUnRdyhKgYlASrcSVXPbs+wDywv
Iv1P9Ihr9+dh/pXkf1LE5NyX1cUZsPnqAZTAHNSjLpXIT0TdYmnSv69fyKM785hXwspodjftM5fT
niro4RyGd8kjj1a3DJZpP27djGIm8KjBJZx+TSEEKxpN/IidLsQPzpdCF8U39l17org8Rndzt9w/
OPmGebWhog/LAguousiNjHnSRV5oErGV5k/oBbklCx9P7EzVeMeaV7MjzTO9X+WMaS4PYl0mdPRZ
Tw2yvUECeLGPwaIXhjePCPOSd5K4r6VABpQGE0Ycj+tZadHcMcB8akjb5NI4DFVJjEWShRtIGjLD
z6qyemnteA4oWsfi9FOPX9vSdsrmNHoY/hhdepaNbo4GrwFZMAIAXvb7FU1ZRG8E14G7XAj/wg9Z
4BufaV6tilNufTpEHs3kmKTZT8s/x/6qdzBcPPjBbKBixtxxqjvAPuyCYAIHvj1Ln1RyO8JxdvFt
V+HMKbSijIQWJxGWuQ/HfC92CJMETxC6ftgSMnbR/wiiZTlKwXHezkEcD0vUYYYRpvG73Q8nrSiw
DGhhezJfgYUw1DrnvO7dSKiuBAHgU9IzLV86IBqbr6T+0AaJuWQ73EszHKNr0cPnHOeeEy5466sS
WYq3Zb88gTaSbBJ7Y6nTloOIV8BdU6ExSo8mSCgKVYwGASjDytTBXRMzlPsPxMWzidr84RwiiMwJ
FGn9suzO3Wb+QOYAs5ud8cEV954edhqmEgDbaNyTuweCkupypfCkW68rUGnuO4hHGQPXeWitaewE
b3IPIdjpdGVKMWEhQSBx/FOWoH5WpVOhyMsVOOMKpZM7xXAtP9OW3Cz5oZSLEKHroQM9X+6oqw97
sVbMvuxvQyAjzGyBZego9ooRO07JRHdoINQtmtrMDOC50/EuBsT3N+8PWZ6wZjePsz1OTmrslFnf
PqcmkUc529erND7WdyNmSS3f6+Rc+L2F60QLNOfUZau/U1Bcrn6ZKyox79ZXIdDC2WRb8Q8/PkWi
xCkN28bNfo0IiYcuHZXb6lClWaWXwYCdgqQzvngk1DNdt3wcDfLWeFG8C0fuy1s3/emJbxlgkVCH
AfE/phECNNPL4wyMaoX977ywrDlIA7QbwOqHmx1OHd4/betELDV49g+uRid/rewVZJhLO2/KxlC1
JNJH3CmRKhbIiV34Z/YZFgDM9O33lEGM/bX6vFQXcdTDtyvbZj1rs6IsqArlrFHJalu3w50/+D7C
RK24BZYEi5KrMmdRFRT+MZUHigDvyZRg5c9UiyPVQxhqGSQ5b7woQz+4tQR/iXOHYMRPbNSaS+QS
53RlWgCWLOUYA5TXVAT76Y+NDwHib9f9BDAN1JNz7q8I8R0XPYza+8EpAThyLmxyjdEPsSinA6Ll
TZHp/Wqr3OAvUaNwTNyccxEeAIynax7onxr9aQ2LjhnIP4AEA16bEC/NspLtEwhb5H4VSmcPZOoR
0ge2KgY/5jbRxzuWnrODoBchf1OB1oJnSTrwy8WGvN72H74X72apXwflUNOhx6oEiSeOXXbf1r/f
8dZ/ymgLSKX1mHNAe99ZdSYexUbtdmpau0A8zJ3Y5noOy4q4OmhrR3zEwhw1EKc1haNTqbggebDt
ZZmTP2eA5z2+/T8PoJG6ioQumUx5TO2xeE6iIEDCSZT8PMB68Gdviir8Qvt7yJdVlqYf8jxomjtJ
jEibgZRBEi5aFryWxT+y6j1RtutfnRiw3XjXCjRwmOQqBe+t5f+eGUBNcv0ULRfcdr/hdipntw73
wbE+r4NEzzn5zwTSwq3mkHnhdOMeKmRB5Qydy2MIc4iCT2t6fwYtIMNFnn/eyXI993qrchpc1hM8
QslUb+bDg0FhWs6u48rGJ4N9rpNsIHY0haWA5v5lLF56qwRwTGMqGxQZkOkYTIb928XTlcJmDPJw
DI91sQYOx0ydIxfdObyO/LbWgC+amh4jWAIZH6CdS4AJ3AKbrLoSGHq/DEWwTbZP8z6I7/ewhiRA
LToQCV0dWXxfUz60qfkaSxcuyOESvQxtY1k3h1cB4160qhJ1YtKZ7lP7VVJDpadAnqFihmdhsCA0
Fwn4CCx21wdvf4LTUwQVENUdnWspMkoi/WGh+/4vV4Rs1vP1VmBu7nGvjX/D9fQzXHMv+ZbHopVc
g/83DbGUl839r4kpD7uSYrcCB8wpuUPoVpEGY/ZDwb2Y0HtlMBmmBiruWJylad4qyN8v6k1Qda6I
LrFMQrF84VygU6g01Sv8tPeT2DMZJJYH8XtXSzmihupEHPUY5/aj3VP/Yibx0cr9fbopBjYNzfa9
QKKyzL5xbW3uflwh4oKi6tewX+hPS55iYhbmBiQyxipNxjsSBfgq+jAQEA8EroMBTKfEYvy5O+/z
R6a8y3VIb4+Q1kDjGTBpbr3TKTkZA9OSbBjm8AkIJUqRRX2HnudGDss+8LA5MNA61JmUKdLII4Rz
rrNHozpEJ+xAo9Vhv62h0rZ1+W6rRi+qhYUu/0wtE6L0S2y4bqFarIj9cZ56Bs/k+EcLjcdMZC8c
b7crIyIfN6YAAbnWJ6dPmHT6aTM75Hcw1yeRJD+qrtABQNshfyglXd7RoZI7YHAQNQzlZH+pTEqD
u2SkPd1S48V0dBEM/7nOK0NoXDnPR9DeNOz52WDhoJA2BPra9ROS6GS/Undp3CsszmcM6svfTNeJ
wxp6PNRsvBh0myJhHrrvPsH/mQljpZDyBR61IW0Vtwf/4MnSj23u8v/iiFJV4CN+7vEpsmoCO9G8
LOoGjGqJ/+1ErsLUt3oyRZ9aHy1b5llTPBBjWssb0JT4ufLpLvgyLxSd2gISbwMDdaOO6P3C3EXV
k66xmC6jmMS/QU2PppoQMipF+AD/ldUzRIoN72ZLRIQngVKcHw2Em12vLti0b6nDbzxNSDIQzrhb
+GlWM+2+Et3Myp/tK1+8mUSxqglQX7vmk4Rk4JEEOexp0BGUiDVpZpHvza872Gu0DXq47UZRmtJj
XModwhZmf3LKJ+23fEu+O5jjWLIqZN6zYWINoIC3CDE47Lh57xV2/oHH9AFreODJix4XQYeEukp+
6svnz9S7NjBs67iRhkxGVFSwyMZSF3o58MuKbrDKHSgqcBpgH9ErpHWuZrzu+Adg/fbpGOI9Utal
6W5eckZYZMGlx3suLzFzVstJipDd1g9JFavdkwzzoE411uDpqqQp/OlApe478xKY9Op1Ovlfvf9v
zjVt3SDaGjX4cUa4B/lfTRQaqBxuBPVyNhV0PkvPXvsPKeXPZkYXXMI4ppKWuQnv5sayMDWgBq1Q
FJz48To/6Z7d+dI6qeT50eIoC/WOhndrLuR9ch4iVBabHwnFNkz7DZRRBCAwo7nxtJK99Zxo/2O/
1685gmYTv6+P4zYIumW2cZVRaGMwZf5dzngcCux5e89/x/WonQrREpk2+qQOGMy4Un90500o2q4c
hVQztdStuup/PIkI6hecQfvo/S6b/hPfCryEnYjsqUkapKJ7hbjP13SKfCZWBXx3x6EktKxnkc6L
627K0vo7+rQBrClwfH2aOk3UjCknGnaZaE3U9H0yduBRAcVAFjcuCfYx9gvViTy0GN1jMWq9BD6z
BMH647tXZleM1lZ+xSXhWuHAQ7z1+Hwku25tx3b5O/aNQ+R4wVsXrVBWKV2p7RVp8R7LzTFsmUqI
kNYIrTxHHCf8LNy6xlDaKecWbEUotfknfkbzs70QujDyKUbTfcKb++pHPv26BnLe0lrXOl23GUxt
vh9VP1LqodxwxVA3lBN0hzJKZ1fCIr3B1oWkpdXRjNsMbCFWfo6uRhVDafpjNcFPZeN9L4mWc8B9
KSKtBW2hkjMRpIo+qYzUKWgJn02CpPP2feNhW5uew4OhETDSTcdBq7qVt8w+HmgC4FWe6UiHqG5n
EvYmI8jYZmC9Rrx5BE12t7F0aJkzRwnWNPv7WfR6xYJco3CRsRFuad4D4YKL+MwTvljqgjbLfBGI
vwqNq8k36SVB7N7UO33KoOdXqL9viTo8ZREoCGg2CALUTNV29vu69n1ZlkuhfIWos+M7ac8/TH/+
aqK6QI5LLLaToPl3VtYY+/cxFLgB8CKW0A3/Jt+lQGl4lGociCJYOQDFM9xHnY30DQXlmX2cG+6q
5q8+HNUnyyVB3x7SO7Y1ESnbbX+9JGT4Up42ShfCbmXVNWHJxPDSyAYMa2SczYWQHumpCR2gA9mG
qha2o2Jf552dKx+gFGkQVFl/AqxWzqL1Qj0Gz8W2aSihX9laayDzo3KNAobaZk3eABchH90saMic
P3JLGAIUbAw5RddjJEUrGN076u5k5N9sFrYp2KTNKeHtiyKd0MWipoyFBPLuGsZZh55Ie/KnRC6K
0lxctbB15ct/bcj9FkroDiHsScOvdmAGk0nZ10ckKge93IewWj+qfIWASkW8rJQjQZ3x/WoeCyUM
pLU5lh25DmzkcnAHg4auHzhUToaBAh6Hg9pTr44yxDC581LYBxD+1ye4uLX9ziKJLSiN5FqiFBmk
dfr7ezArW6aF1PRJEMo81ktsf1s4439P4Z9aoYbhwUdavpGj1bzEyfDGZxFZS7ACPbb96JIrjzEs
5TU2lF4NXOsUgDRtO6y81aPo0QqkY5ynIGZ3KTiSCfAhCrLSl2NzmS2uqAT377J9AhkUsGj7CY/J
YP5PGdvrnY0WQz0KmEaxwR69A4R/F3wz76KiECjLaJNqfLME8Lzbay5JSEwc17+JqjtLF0nYJZRc
yLt/qZBo7zf0mZacXUzz0twlqcCD8mSB7GgUR3gDD4fZ7nNTrFKnJF6MkqtBo08jBiCPTE3sST49
NftOj3fzZGlgJ9BoXaM3pj6tIZ47wi0ScMVoDakv3bbmpTg5YDASImVEpAF4Kz3EzrVpWOXUZJ2a
+mruWYMLK7f/859sj+zCcVcg7pTdIXlFml9fntqtkFlGVwd4S8DZlbVI7tM2kLPsEi2YFTnFzFuM
jh7LIsmhIicEVGhUJHC1Qp3dJwsBQTNibykUmasK43B1OYwhoIPGyzRybIpSRnWH74dwkpP+RjU4
6c0IFuLPR9GqYGhJAmhcD0f5AukC2MNXUksKlRuUEtPIj1HJDQR6z//6II/3zyxXGOX56A8ZmvFx
r05vbJ/I8/3sAx84ObRfLAoHAXpFq6/lRQDpZo4S6GT9X9jzOy8o1eS6FfOfSujOzo2ZaF+vrZqq
UiYsOb6jdH5MKzj2QbNVo0b6TbnXRKzhYam1DDiWqUzoaMAgsFJz49e6MUqaKozhdBAq0cpF+7TS
HBidVnrx+IMMW/HgGg9nf3yYBpBXqtWus/VDzm/t7hm+zodOmq0QDF5cCFQ18+pOASvTaEtFpzUZ
aY3RD8eMkECGsBAc77xePwE/jFnP7BZOt7v2/VRUAT48UfuS6lWkYCb1Rqy3wJ5wSA8xrfFPxYve
Z++1Bl8S90VxxvXXuzzynESa9puGIt4UzAnVChPSUrqJpzdWB8N4aWmPWDfOqfbXODV69fF8tk+z
c4+i2X7iC/fITbT3VJ8CCCzpbjgJVGqKxh/eU6KnpW1rRtYiIV4atGCuMD7YWOwLHwRY4kXXMvXp
hWgS0EM8QEYymboU4pSJ0CWOKiIcPGVBRHSFIiXsBPs1fa6+bQuquUHDxDdqiv5wBPu266Tg4xzv
gc0hR4ffF0lsFca+zXcEPz4FF3DPrBXx5INXVvNh62G2RkwrwmK2gsYpp+ArqswlPbw2Le4vq6kl
G+Bv//Q+UBwRdCvfZ0t/OqgP34JKHgVRnGh5KSdh5xTyPJg/G4HWq9g8iwPF3XuWbpk+oi8gQ3YK
s7/nVW49UkIH8Qgt35LTqQI6W2S03fBrQR5HLmcEITx0gtRhJrp7let2t8fOS1TlJxizcIVAzj8/
SwAoyyvoijYJCWKlrTZA0C+X5PprmoeKXqQDXwXVwMonvRPZ0Gl1k2k9ecveuWpiaE3Zg/Fq+QIE
Cj0nwO4hrpxNiV6CgLfrysTvcsYj0KMF8MkQb+ejuVkNZx9ccOGN8FOmVnulHVOvnLH8LVaCiJs2
aziL/IY2wsYyZqhri9TVAOamIRtOYGzq1HQNZQ/atlemsGeTUoaSri6plIDrORFIdXnE5SWFD7NJ
Vsdz330aaXUa4gxwdHq5a9L6+x+kWy9QSCTBzcvogD7QKdsMfFQtatHwe8LmIgugoHQnB8OjJFJs
q62W2CP4lC7AlmMo5HeD9aEjC/L7ZyeZcGYtykjwSWl+unj2RAuZMemoyG7xSaUXDSL8LNeZCawW
25qHQMAUW0TaYBQUGRAHCmaU11GptJsej9YL3UnzIKlRtqRO/4BucoXyhuQ4nW8HFhDajM/yprzw
yyd7rs3UDi1OkbHRm3xBnOsR42o24JOvkraTDY3mlUzpDivlP5NHaWkagtdH5fIoGXr8Ofjxz/ME
Xycu+He8aw9OqWPlV3W1WBoM8Hg49oJPE/rp07mP0W+xwNJlYjv260nJoht+0JdvaICsTI9/ouKm
GuLcQ1VV/wwqLVUD6wHkWrTOPaPVFWJ/8ofaKhgdOJdmwsQpInuf9YsU8g2YBs7o+fOKdgUasA3A
bhaQCtJ6AMVvhTiCZ+2r0HML9gpMZMaaKBbG6hkizUNtZeL+0hNsVondYdMQcBZEFZIYeJVdF6Rx
dmTF/AvHj08vOX8O2wZxAC12mYhIuCDRysIj+tVmxn5XT3rYo/6t6iNUeSK27HmOi8DU7irhd1oa
Zn0g8OhENCByjeBkwRcAKnN4+CqZ26SyJYpGSt1eN/pUPI3UkRxf6u183+OrknVxQT51d3tMYJNp
qgOw4npF77lf3Ra2+ze9UXH3HnC2fCRHsLsNHSgS6baLh4nPECfANEqDlaQSpz29cLq+tEBBjxxl
AoAFp560kRWZHKVZezQV8R3lZy1YImNG5/Ddf7rKM9GcYoU5F9Rm0KLUP3Gqz4FEGnxBQaleTcln
of09eB8BKZjVJowJMCvuBDpNUD1oVQQC2q7pcqckXXzjMgpjpsOk520GxJdsyPUJZ1tvMBPQWc7w
SE4ODTG4Q7Q+rQrMA72brTpuL8xNYHT7XH4GpQftajIJ6H9Lm0nZh6v4LXDSlUugN6mcWDh4r82E
DEZZ1GmWlEqRB+thT4PhXbc22TLiQ5l2r4rg8HjWT3kAL0Ba+K/NoeItzkT0jf3wxC3ZMvpva0kF
9jPC+39NokwdK2nGw+X2hNYHPa+Fqlqr966PHQTn+18LsynLWgprJ/iZbBNCPEG4HDXCHymW4lRp
G9OAaQFxWtMk3OhycmEss5rTiWkINrZ0SvsNUkVGs8XBIsIyfqRDXXfkPht7Ky0bYdhvUDYkmAgG
dZRqkH+R/HQztUFHC43NlZS5lQY/QdHNuVthC19OzKRfwF9diSJKVZiM3aByNF/slFi+GIaB+PG1
+tsPpUFi3FSMZT2gF+A7DPu7X5KgwaC2C/CZ//AnMUtmTBphU8leO6oKU+IwXWLe/I8xMb3euK6k
zQ9L/mFCQvAHWItRF1l6n11BDkOiW09YWhgQX9rlF2YCX5rBOLxhICaSojycpe2wD77wO4K2LrMW
55H9cSsOfrhO1FxnlP+5b+egBh0mxqkioJ4BjRmE6uGy/gBbkzvSuJyHnNxesPQqyVpjocGSgGOP
JqhnmfhoSOgVTXYETTq4m9ThY5U0iTQZUbdRp9fHPW6kYjWINCIrvAft//jbG7F9Xa3C4JAbD/d6
3uXbVrirE92w3Peb7sJSt3d7Nl8lyvQCOJX360x7ACu9lkDBWevog9GDeFrGok1qC1b9UsPAMlIC
K3usR3tkyELZItYyINFN7V7Ovo2OUh0ubGkSPu27qb/L1DwujTSWcXD+GFFr/81UKsOiS1d0yDHm
PRJA6c0OdMoozBNW3ARd8g+52MAdxnUzYOpcdvpF2B3eEy4CtrCa74/ARlTm97C2sSSB7oE8YudH
sqdmgqBbmxWI/llqqLG3JNCzhZ3om6KAzuWOxM3s50HPnzlXlXN2D3HcFS1XAFgUx+rhuId+QjYL
kExM0utX7ublPWmzfadtSSBRoAN09adubQ9tsbJHCrZ5m+ich9aC0eXFZaaWcjOj2ifWAIgIf9AI
UwV2a5N/byCucuRzUieE0RwXkwlH2rv94fjNTDWFXuS7gk+JYXqf9IYIH7yvw7+2R+CT7RgViLcT
LlSjaw+wJxpjCPFssVNEbZfzSnu+lc/G4VUP9MBIICMrT/LmwHVnpcZPiq++adGB53dXB2KR21Ih
ikvn+qaT4PJO7JDFw13iFYj4H0468xrGlMb3oIPrE4k4PfrRnebhZc5PRUj4KI/zgaqApGewSzyc
j6TE2nPwl2txraYTJI9xPaNOTrrdJJWE68cYG+LjAiZQOb8pvucIEmsP1m0aHnEn/tJvTeckNeVL
s3CMQadf+a71+N9U8rGFkRxxu5qmo52Vd0XEk0IfYDnlVo+2JFnETkbFxTmew4dSAdBrX8R9Oi0Y
pXB2Cdp1YSOFZgkMnE4wdXgi/UZKHaXHiUZi2p6wvJf+rmxqeLRTrR5jD1rscdUExW26/Uqh/vhc
tJqVLSKK+kj5rcco3pjyblPh+FKnoiU55XS9U6WC4NOqd2mVLdFk630Gw3ZJfKnIY+r+5DyhoXfT
AFe85n6eRjJrsN0/BKB8oJs3a3SFCGAsyK9HUGrBBoSNgTmyIjeoCOKMVv+7EQJ9+XK5Q4U0FNcS
bo9WPHFIh6cD+s7sGJ9AhhIt7EVm1URmurVUJViAAfGL1v6pU6vSGAzAJKGEmyiOS+W21SUqWOFx
KxSqm/qtAB2fAQbaZ6ukE/mfYfwszAO2+txZEotn0N3mhKFcfSGgwHsuRFwSwlWLEHcQBB3luY8Z
W8RCA1nmQW7qctZ9JwwyvvuB+O4Q1AXNVLgCKEAbF8OxP6fRt61PTXRQgQYE1n0UwIUxa84CKyqV
Yh54S9TndXi9z51xZFjgHBn1CRmeZ5kdxVc265rBWdohEGy1EBq5bNvXNGzbDuleh7UoNT+Im1eM
Tgxhg6gnVanbMK5jrfdfInd0bAeO8OQKPtvUI2JCfTn5KGGFrYOayz2apH+AOwKXLtkulgvUkpH/
e9Z7Tl6O3DjFhVETgCQqygfhBdOxVlKvqvaZcQysw0WC0fb7RjEk/zLx8zd0O1qgQG2RrwKCk6Ey
TK38MuHicsgaAr5M1IoMnAkj2QFuYeEqOgzwODfrSS1DWWLjp05h2lv+YR1IzaQUVIiH9h5FtU4T
Y+ieSPUGZh4ASQbAY/MStHQ6F4LHxXidunox0broB9uy8aRhuGl37Lw86iDxxZnt7ALlVZsnKWcm
8WpohS2tHMzI02W5Hf3KO6uqhY7CPNg5xxeCVLJzISbAqRWUTVRqwMsbU9IsVw6CQcy5rk2a4tBL
acSd20L7T7ptZBjFBY+6StlWt5yaL7dl3z5rQZBMjCHh3txekqgBs+LqcvSb5+5e16r0UCGcieQH
9a2xpzHBQqhNwrQQt1/7a/Tawan2sBBcUVhgYhbwb8dbcjugE1oI6xELFin2Oo+zUGcgPYEAJaKt
f8YInRyf+n3ZyKpgFY8fPnijdg7dqsxWVBazaQQzp0p4TNOQrcABiD0kqNcflH1tyUq8xS5z24sq
IedsWtb7HZkDTF5ym5LyK6j3qFub5BQ+5qN6lWlvxtMgL3U2bYR2ffgPx6G/volBriiIFsKRkaC2
1UCmbFnRTbxSUfu0AlgM2uPOx0rncadtMzPdFBv58DqRbOHSihl7b+yOAiT2ZhegmEt/t/mWzt45
5V7dCLHY7Eat5J/VlbBvjrM8NUJv4o+G4aKLvBVplplbgXWQUhQ72I2kGLiizP9gCq+uHDR43btw
XeW9weuAJry4X4MXGBo7FnjNETvSfvKgU/lCETgD11Avm7AX+JFsrVhYIlKr+w5ZzKJ7o84YPnG8
il2HHdDXSduuy39VUP0LsJxff0FS5qshTh8asEe7CRyNnKKTm6YvUjLhB/NnXlSmqqqqt1IN0OTw
eE0gdjDu5RRqEooHfWS3n/VllfkLLVe5gF2+c5P2BCQtOJFmr3p72fNFlA9oh7uIYL4NMK89elnd
6ilCA4NJ5f50ramwoKZvM9EytNQnb5DCz4DaBlq9aif4uHdo+QhJeQp90FfB0VP/CpcI/bQ02EzT
CdMLOxHdb+gLWWlfA2YRkN+n/a0tLav/Uqdflkq++FQ0xJ+EKQOchYlN8ClDPWmXyVzmtqAflvRW
gQZt9MF7PWthk6ZS184YR19Jf2lPA6K/fxewtEWfzsoPZLc8dA7l5dQWkMHepEC2R0P7Vo7b/hXu
g2SxRiHp+erKzI8Q15vslP9lfxnAMmdB/6DG5vMh7SYnx6+eH7rBburOOJ2jM4D86z0tdQ7QJb1i
wq4Ij+jwr45tVmQ0T18V1RfEeQ+nS8KHZZ+nx4pWbvmiQgDnVujEEwhRY7a8dd4GH9NROUAoEGAl
p8SJbwAKLXBi8t2/95+Ip147bXMTr1OUri/3kg0nMzsqmEUT8MZJ08V7NMnRnqPQTnKrwFJsfQ7e
cgEYPUzxv+RSfSphgXEXThZK8gXKMjdsm+kxlfUOnF0fuPOx+TJghg7nCSs5Cbc1OWJnTqeCoXpo
WbYF6mW+vRxtffXPnaYOShd9X1CYsbJLjBjNvEbmSnVGRb+0tHIq9BYA/HZCBG5yVGaFoPpj+gG3
6YR6MIyzsDkCULeyQG7c03W8LSIpRpjQ0o6hjHresBzJ/SCTj0mvfqW9hkIixrfZ4gsit0bijoqP
h32sDCFj0ZAg0iyiWiDcqFZ4wqDZw77P4pj6miI8kZvMeoyYCaUeKfDOAu7M3PP9NrHBRjYWypRL
49eQWpWiU3VQ8ILwn49UGd7FKDm/oJ+AxCJXbGmnz2bVlr0QECprNq5Enc1dE9K2K1WK80a9FXH0
u/DYcl0XwRRtwoM56oZt/JNkUQKRqqTYAqNyi7eD06Gfh1ssWK34ugjBafUo7OxKxC9wNKVmJRGO
ZV6KJwvn0Yz6/0/KTKPeq8oIjaX/9igtl9ut6dmHKnKS96cOYumSxgvtMwNdLbOBfbsmTvYM/rjz
qtt0//GSLDL6istdSerwMcChPCPMaw2rNUiplb+AXnnu+KMip+MhMi9IfLUGdIS6G1L1Tm93jNGB
opOak9GvC8PT+PT15OA2hkbAXzRhdgGfePR2dcyN0UJa3AntNLzSNGWznP5YAQEHNJU3VspKtzHi
7B41vhXYNuMEwbV5ZRpIcbb6I0DkpaQmOtIyLVCHdQ5xVa3442CAr3FBDWSlITj7QtsmHRRRC0CM
qPRnNwLfBKYktd3j6O9PbNHMXXGK3QV+KBNpCByrMk3apwacdnSMCZbxt13cxRclOYzSki4CQFmE
FaxgN7ZGneg1Dxq9DuD6j1fh/oV1VxlZDLCV65UO3mFeV2owi283JJrrWM3BbG261hC92tTZGKMj
f9znxEaoqJIWInm+Q8dBCsayUJlFCmXCNamH0IHYX5q5IVVi28amTK02FU14NPwu6Nv6EG/rn2NX
8fNQUW8578OXp1g7mTl/DwjXGlBL4B4u/r3J7TUo4/4H3Z0Bcxehu/zFnBsRBMulIHvnBZAdXaXd
j6SmVSFJmZE6qeUsuArmvuCrokypglpn55RwOHgVbgT6FLfbT1EuSjAcqDTdqFq5HXKKiVjBWPAq
jWD1Q2ru4oXOuROlmTF8/I0AuvZcp5YHdcEwX3dQTdZIvmRnORPVI8LSPnV0Zv/hZ5CmLB0cnzcH
03Ty2IImJwqncknCUBspGp1dJTcYpiOW3+3/J+mrlhIi+Cy7qPINHEdcBdHCI28A5jQfKoe8GarD
fy+b+tMVMkx77cg7AB5y4MztJo3PJYSwTmlQtJeilGkAuYPbq8yGGDtRDnrog9yGCnEJbJoLQdsL
qow/izvzkcqV04RPZFGSjKnReTrZc9x2beGM9Kw0BzQdzVgHgXhRlKB+u1fbcysXIRRBhKXhOFx+
JnuBMCyJNnfbURWzC2XRooZ3rOt9tAn/DE7/sxrYu/olYwSFdoiAOMcBUh9QYxwgYIhLREFGrk7v
aBDPZE3KSzDeoosDkrIsai4RshQNwQz+o3+UrHuTcE2ubRZ7JtASCuWd7MGJ5d70qhjjBd0Bj+T0
7CN0KmAg1cjWhlEtuPezKYCeKREgxWEFWhKgL250yOmVPnYT43wqr8gm1UUDSfB/oEpE5RKX3N2a
Fwh8tZZn1SXTWf25FvexNstxY7S8Cz7tAZnfCtpgAXt8QKdjhL9BQggly5XycRyADTWdjZwi1pd5
h0KEuowuMuYZWmN+xjJfXB4Q5KTOFo0CZxiWpder5tYC8GXhTUUNLrwQTrYgly2CqXK3aW6JFzJo
eJ+0m7l5MKtfhYw5+5cicUJsPZbRRqtuHqSGUbOrdlWPOIPn0kHIH1Mcx6r+mP5BNFos4lbetIde
PPMXeF8elrCgN70/jxMHthmXxbbm6Z6fjIGaNmT+8sEEs3C/58GPapUeXCoNWmIrX5JfuUJH7221
hgWm71iX56WJ1Vm43n4j7eZK0YueWr2UIMBn2iHyqgOJsMhAuzrvsaOrdniZf28HcTy2fRMMBdz9
dCARAwUdLQwxYczdp5q2SMyQO1tf3fKSg8RT1eOELtG9qjKmjclTsilp+sah4qqvDYXNQdXDFZc0
Lpuq7jAIu8cEBgpK4IE009S21GXiT/c4M0oqhtFbbpPtpIvEOzX422khn4w9jbM6MvT3fv0bjcFk
XTQK6i6KzFqbY0hEIj0tD1tRXTzhnqkvldoqUDMSbYGRONXI5ZGbuTAu2A1YFA4QooHzxq1ont6x
IsRoeUNd4kbpEcpkEMJcRPgE6cF6P5/fJ+D97wIuWlN+oKWWl0VFVaKPvjjq5AcX2cslSHYxbLyY
KmyWu9viwZHdvpddoz8MHFyixl++ZgYq2fn+UEAp0CUlyrLVYYMPGZR9BwLAU+QWttVxEuJLk60e
aOTVT3KhgwVu1rHyOalehyrroAAShCLm3Oa5pPzh/MXU6GNmer78V4DQ9jHQAe1ElksLWRMwxXlD
a7kYM7I3fcNVNSVj9jqZTMtQx+sEzBZYbAkTk7nNqkmmpXcKeeOJ8yr/JyxZ6SsWMO/585SicCiP
knbbpU4jKo+WBzFBG0UvyyAgH5P9KC1f/Ym3fNeiM4XU4kJLSHbljx/LMnktpbnAiXIoBOu+P0qJ
cRvwdMaOqu8p0cyTlmRX1phM/KIMgLrCTpqRt1ZJ2JuRoDE9/vOfqHw6IlI7ELCq4dmjit/ilGo+
A0c87j0A+goLDnkcXtcfXiP8FQWzg+xReJUkrmfrr1uRXqFZUWPhZpSi1fO2jDeTl2kKcnfornuY
I3YhzN65WJFfYFS+vUWX+no0ZkArfZmKVM9jIn8t4SRQIGkReb2F8IaW9Jj68reO/GAcVF6jHCd7
YIGU7N4VZmXRt0G/7Ht7Avp7DzugJ4gEDquizeyCGgTxnySJuNDzT5ebBBF3cVmHCyuV5ilBbqsh
xcSVtO68oghqda+NI0mMc9qPcKUof3ObTKo0YrVPWyVcKWBAY/tWtWk9HbkabENuALNPAYO3oesq
n27wd2eXiWujeFCN+uZq0RjFAq24lDsgsS7mWC0I8o4ClBR8YCtaB6fuG9d5ubPN9ds4x/jfdkx8
cnepfrZ3MK6t7LFNz4f3DqGDT+AITd7RUVrl0sHfmgTjBHKsRr+73Pj6Q+tWBHTQ5vBBkOdaulG0
9yTaVqD7OG7uDRfuZds1D/OAJg5gwijg2SoJ122VR2ZwKsmxtyPfO+oGW5uAq4sSCllxxMUdaAXm
3paKo5wwPGdiOfzkxbZ46GjVEJODWoM6Pi+jNDiVYGXfX4NazxSOOpczP5Q1zKdmGjBiVO9tUQP1
MUFm4ryK9wvGrhd4irTnIjI7mBAcRNGvWTe/Iof6A5fOlsDvbdBFscbkYxaWJGFCjgoww62hhril
+t6lBBLTeSsE5AAnIx72sx4ZjYnYpJnmSN5Vp+W7Lw4HBbvp3k+dZisbxQijUYPdHZBwoHeuck7E
wsyCTFr5YNrWEVebgUbdZWqrlnVB8KR5px7yoiplWxAAUA/Yn5vzYOcrqqgMce8oz243s0ARTu9u
vUlJaRwbI1m4fLvQrOPfjGiZl/bLlVbIw4UplouhMvIH0TYlyE7vLeJohb8DOwMyPtYWE+ymj24d
XbvAHz3qe29JIykq28s7ipJ4eh0zayb6yzoG/UPCGVNy3N07caW9jVbEHBZk2GD7cipaXCNSLCYQ
ehA+LckpjtTNOGUYui2KXvN3JY4SSXAxWusNTAP+pa+rtKuvYgcSj+smf9lydOUFN1CEKbDSYbHD
cQkQEKoYeFLF+yBMVERZTgiy0eZ4EVnwMPiLmcQXi3NcZXHxfavJzBKjTVahV7+CPsLEAonXIvNg
E6MgmQI7HHQRS7RIyGFhwOtDvRMWU5lgVPPN8JDIYtQKxxJ+k+Ik3KTHJzD2uFnKDtdbJkGV03II
jpGWr1Ferk8RijBuAWc6mEDpoxMg6GaMLHOhaHUDShw+NTBL6XgOyxzjLBSyZPteiYOGvY5K0UbG
szSU8Sn9h5kTAaJR5Bs94MSoZiOQv5hM2IucOcoKycSEu3GhmN5qtBAlVm5/BPok2cZ05enjOKz5
okaLqdmVyL3wyWSFWSpvg+iMwZquRmaUzOZZqVWiU85+tctOCsWqqp0BQfr8nnx45MdmdgZLhyAv
Ylzg4vBNjCZNVagQvNLnGLL/XQIRCnQOeUW++pYHpzvp8ZsjEwc/jQcsfpMoHI1ST4Dlt3eFoRLC
MtlHXZt2JP+H+fPoNistHP18XhbuRO6WtOo9KPzCfZKVd4b1WkdnCLMcQXYMtUNwOtT7fI08KeFY
diIWMHavtewUEmw1Ek2P68b8O+d9oPpZIDyuQXe6h0eRIq7898jG4Wm8lTC4bTyzvK/hCupMHDlo
XEFLS/GXFU10Iv43pbJccbuq4rhdsDbi5QW72JjNoJeLiTGf3YCABLuKononKgs5lwH28wN+E9D9
JsGkRiuO0RY0sWBJ827PsBibpghkqo32vne82WlmmsWCz+lh8axn70Flr3VKHVQT6CZTwH9+dp1X
jGWEa8/8XDyWM5Nb0HZSKR3yNuz5Yk130pnF7XUoD5wwFauLeFMXzWlxfBs3QvHfRYUbnYmu/6mp
3CR0jz+HKxIRyGuWNwnu16tH++0LYAwVRjT1SktCymCK2Nd9VyIKHf3gAJsHQ1bxdugFCO8VmZbQ
y2CKV5jBXAKNqZo5KpuMvakvQOYPS8jHbPTP5mE/SM8upUgrS1zRzQ4HIdioSpFFpKRzYvO1Y7aA
PFXVNkd5vFukmd7hKlGu5d6i2YwDZX4WwELIveGIkiAXY5Er+kUk7yA/DDwfBVffE5zfYI7Sx3Mm
Zwhm4K4fi4VVEFFT+pce5GuZoSuv2HcJW0DgHoY/sGIJEVJGvbmzFByVPHuyh+TdVAKvhfLpjFoX
UjhluuqNzqXNCPoBcgEUzG05LHBjLDPPFG8abBatiQ/We8yiDNakcZi+orQCYbFXioJZZaXr48U3
rmBDw3VZ3InWFDgiLAd4oTdRc0vVjeq/pcwdlyffWYm7n2UanMbQoMLq246HMpm1TINcC+ObQDYp
CZUk8fcckQKwk26CwDEdsNHULvliS+zPvw9+DkAAn+s0xmIftj8UfYxaldoe+9lLeE3W5RMqJnUI
3nnCjT9gtrPcui7DHPmCpxM9Jm59EJUJ8O6bYmpuTQ+YDQe5aYYxRJLoKDdkZYqnIkcYIuvKS3S6
5YnskgGyU3N5YK7x2Tpbw94uMQCC5kC/s8ejc4BXcT+nO3R6/T0yCFmfq26KanXILU70dxacTUDU
/ZGvz2H0JCN4jNfF4kZYDu+uMLAG+3I54Zu/DVDqUmX6dzchMOtoEkLHg9hoRoff+FNREeY2706/
jBARba64bYCwZlB5btHAIWcmzUQyOlZ3RNTsdksp8/E2A1BB2BEImmfuMB/7MsvMdRnuDwKv0qb+
zwG7/t8R+2j9gF4XvNb1HIxTm2v6VRQxQ8JfAuTSA+R+bNDo/X4Ysn6bfBF9GbkJRoNob+QvSvfW
+iyS9OGIMosaHXhNxq+B2Wbt2YshNmU1bYJyYkGQ9uOBB3RhTCXmE3gDuApQZhUnIMn2RfstWfCq
timEmV6xZ0rfQVYGvTxt1ccub3dRvcoYYKWHl9cdtC+ihW8eoMiayMcpRDxweq5yPcUSUoBAg1wk
4Q4nTgphYmXgSF/iYDjo4VqlBRui+xh0D8hPZKclF6KJIsV0OIffjQaaZxsa70we2PxqnV2qW92c
pNhWyEbjm0qfkErXCdSIWCowKHzUmjzjcNZUhCkg5cz2sD7ktnJFjLaHM7LhC7w/v1/TQdylahsQ
hLtCzmTOc58UPM66vy03K2xmPn0yLec8i0fFsvY4QXuB/Uk72cK0q8FkhmUQhbvNbKFH3eUZSz/Y
zERyYw5xgJ6zJZdQJsJorlfwsOW6rHeVK0ylt5hbeJl1JEaZAFiGrGhpyHQAi4ay+a+P2va6Qrvx
8CMMl6RTlDSWs8iQHrTD/TGd+nrc8O2+Mtfv2H8hHXY1kdjbY1rprLOyemUgk+xnR3yOFPmOzxhm
Rx/41CjDaOgar7PEya4CsbgE2uhe+RxPOePZITo4mYqAaWXsBhPLNXzEUzJxjwGSmb2O06I3sW1g
fhOMAxwyOMLs7F3iGmUchWs4O3M+PyLUHVlavjS/qnYlp0g7QshFtfgIlPSLwmdJ9Xg/CAS3z/Mg
ApXKnawIKQPxzNOCWlXzMqE0J+px0sAVRGJ8IQN2lhG4D+iExo0i9XfauMXbvk+Nsrg5sBpplFFI
QsRVrUU73s1D9JrQNQ89ZJKVnmasMxpLp5EqllO06fnjVJEnXX00pWAaH90nxh1MJ4WiDKAMJKi8
aIdB908j3nCns9LH7pLyvrYnWL3oU0vMVM8blNfydcUzeImyKnh9x9+pGWWVz4YRD18HNmszswla
0wjQfhvLNPfc+GvghAxQS2U1Y8+Y9WtmaiOZDSxRlq34SpQk50sRKYtK4kCEbnzWSh5XOaacIRfn
UUyZpIOjTnSL7OMrpNuIGAL3pQrkybCLpgc2+u6kkSpom/RW6vrsXdt4zev22zZEwl57uJw5NG7g
Qex3meLaxVmAxigoUPbTHd0O9U+7xy5o8Nne71Xbtr/JrncrZPZ+VS8p5YItLjtRFB8Azp9Pyrp5
HnVP+rbiggWnLzoO8WAp/23JNH7NUF80vC8hqPSex5sAKnsKr+W7x2+e6SJ2FlGMEL0dMP2+GbTH
lAxkdgSVRGiuEfGkMA8Pp3ndGUyC5+wytJgj555IGJlgVNMKLLj2Og6wYPD0GqGg3iOF6AucikwR
SQHEKuD5b5WCPVnqUJYAlThMfCDwjuZXqr3tTk28Ll0Q9WUs4yk3FCvEweH/6EVXxlvdkxoz9yNY
cL8WrUlTA/JnP15SSvYL1wT8TAfN8K1AQ2LgdPvmCvnZoTYEeLNe5iSWhVzKeOyI54dxFUUDyrV5
8cYidRbZqGTpaVtOXJL8Ma4Kl+FKGA2oyQ2nphohEzH2XYsrMTEkvxsRhHxku9Ewh832XL4EchWE
mHrEgCSOseWWvTzhIo4pKYXT1S2TD/JLvTEL388jwwVWjkT7kF55RIP+zzgQoIo1j7p4etcyr888
6Zm6UO6CM2PTWCPVkGTrZPeDIaal/GeIkQXbM8eLQBYopdFzSr9LYkysMN6BdfnKefOXtHJIYSYT
8MUFaetAgbSrmw3wnIo6Q9QcnWHkEOB2cUApaJqK93xYxfK9jnFmZ6Rd4Vvi2mXzJf4JjzcBmblM
S03W+CsBkaxHLNkCtrAdq2bnZS1PhpSEUddUeD0F6gQyJ71jkcxQNzYbe28KIx/OdGRhjRR1R9Jy
DShZycVKVwCW4aMkpj+u0TZ3fvNuB3q/+A7mrO3DRpibyRgOrzvkn2vAneMT40YzQzVhEQXkFs0H
8kePp8pE2ejSbelepnY0FTudE99nNODZuRMwLCBM+w2g1kukDxJtxXoaZqZ2BexnCQSgwHqAc+NZ
YMH14WiUtTwFMzfzxRvjx8hPzeKto/+6X5VvbCbMtBUBL/laJNEY4KdJXtV+/kMl55DVlzc2TW58
WiIbqNpX7Vu2In7BkCZBkOdZZDDFvHlIVtn2k+xaQfna2fn5PunN8WPDrR7Z3rqHsomQS2L+enEy
MvSc0ricdpzGIuuTjS/ns64LFMXGD6TC+La4ZX6K6ae8/s5e8Z2kmWy58HzPHhf4q8KHRp00bosi
/P10kN6iMeLrADLMACbqUj3Khlzs4erVVtql78CzGYM5WuBenOYfYEy4Xb3s37iLgvwX/uuEnM7A
JzWingD+pq+T3eGI3XXDtKFtu1PDqjWlx9D2i9cHX3DseCSDgfoi8zwo0mH924XptIGDmNxidwKR
lKx3FQokVu0MdXXmIqG37ELlTTlPhXwwlj78gXeE7Sd7eOuDYdQBH0k/GOq34fNHjrV2HqvPiUeA
n4OFPQLghDu7dexWcfQdpqXT4WN/P46VbgDHk/XSev8ZNC5GPBfB1Z12tG+1z/xLl+Sb3cmXhZv0
JtDOcFpyH1xMy9uLLCu7Ij/rHPOyTkgl2PkdDBN1DfDIXHXU89+HjIgH2GFAf4YCiOGshXkKX/FX
DBSxT5xER+Vqj9HeToLDoir+sSEU5M7jifggg/lWnCJkNfZVtpacVPd9gAaQJp6UIln7bxUy2Ii5
pi/U5ybclbd0CwzfmrXH58ZtapjBkgPLxD+9evTHH50CSI5JeFIEFCmeYaeXgyJPK7uccN7MRAMp
Bod8YI1K4SpQ0NddWYnc+78/ce1uWR9gKHP9Kuh5Kb+SHOWL7c0vmn+C1zQpz4iScLXq/majPz3A
SZvlvozophiuNuR1QJlQBD4SjKfvYCB3MGr/ozpVwmzzIBgkrKN3Zmw67++dAc7XdvEAOUAuQfc2
kqIJSed5hiKILhwMzfvRqRKRgleGaiLou5frfygpug3j0D34jKFp3bGoiXU0spqUxmvf/nNNNaDc
6EKnDlzShQ+PNFGZh9EdsDalymKPklJQ2eMXpzo/6+kJ0dbBZZrjkh9gQ4WgkaeSSwdahNHxxQWi
J5sFRj+cti9KVdBv0eL0XIp9dfqbMD34gScqLfa63bu7VGTVHNqljbK6xnGrSAw21UV56bWjq1LU
J9pNtgld0O52kQWuzUjB5jAR5YGl/dhOFsRcHHDX/Ot/hXaVVLWRpwzyiJDM1DU9kmw7GhTzxq1t
5a2Veihc8SMxOe1q3WxzE6zr45PeP9DCgJX7vnkYw5jkNL9HAp/DhS3Ay81iRmYGu7jTuzaxgtkD
rkXtEYf8q+X21DEKVedpbT3ORABJ5DQzzg0bmb8D4zyyGdAvl0qioicpm2aEM4MjsVcG/EvORd7m
XS6msxZkpYJQm5ZMw2q0fsvmehZgI1D4pBVL9FeP7znNp/IvbcqQhiYAtdivHvNoViiKTBtoPT9i
IGWkCP1MsBcdUmEP9yZ8RdyT+Ag875g0hUpe0+xty/26BbXCbs+Jt4ln14+sUv4hunQsAbnsIYpE
nioPeQE96SzAyL3nBISTfCHbqCN+SDvWzXnVwWhcr89VoIGh+Q56KnVRVCx2NHaMWoAYpTPBemZQ
1p56FhaGbaOxS/Ln5X1GKqkcwYgGXFtTsH7uJ1K7726KMhXNWCHhMtYYk8w8XUGeoaZSzS4L+9Ng
PJ1KU+G5GAD3vMDTIdN8NsrFUlBB37Cunhr8FHvqL3k7onH8p4tgTxbEvL6MCbXDPCTDMrkP3VSK
xsoGkA/GGxS8qW4pU0jPBVbT2pf3azycdAuR+4aJt88e/V7Pr23v/a9B0VawuiUDFJ80colxk1ar
iPC37Sgp4gZMg8yB3BNVX0n2KBTIAnYmUGfcEoX+LeQH8yPVjusYWBCr3L4FSA4FPYFV9DXXzE1G
zc2vUrrVhaWpMR0m9vu+BGaKYLnsYH25TAj5VsQkGqShcIPM2J2+vY+/R6IwpW52S8flDDlPZnZ0
imWRTW7uaxNG5gwzM6uMWE+1ZuBQnvScAVVzEuIgVVWsi0vYYYwxojCItFoKryxvuGTox+NbwDI2
s+tK+OgbLV52il79ki+Pmt7EhBvWpTpG6DM27bYMy3OURWIa7i/cynOimk9cSVN4tOnOkUActGrT
Q1IbcAoW/qYS889wIKHag/Cda11ntKkaygnzdumm9e54ovpVG4t6NnvM2+TXRBGsVUhD0uiwHdQD
pKLA3HcL51C+BmrLbGKhFxiJJvkIrXnh/CeFnLtL9DFV0B3Kzu13Zz7Jx8KTi1331CNQ4wJ4NcKy
nYO8eKLEuTyeinx9Zzpa6d5s409XbtJjyoppJncqBYH7Vvz63jBUzijkTMKkta5BJe5zqX7WRckl
hWDEJPyCladzKZuSps4sQtHAoT0HuYERZUwIat07N+vH24eDaR4rrfTcpk5nL4yaxG8Rci6J+9FK
+IKfP+jcSz3BJPfTYFi9lfTm8RszdtCVnhqcekSlxVqlg7LHcvlBt9aNaE4T7n1GbhACJGah02BJ
vp2aI+k/2THt4DnjhoGVEXlAKw/08Lt6EXTxhkOdcZNy2EOIFM7VFPVUbMxFmr6VJM8jhCQrasSl
0hHj+G8mcFx9WnCjFleMEuQBb+gvRUQEYKTJLgNu5rWy6Bfttq9ormop8TxG+yygHAkj7QXIHL9J
XtY2uEOFz7QdF44W82GkiBZt0Ujnwk8h3EYin713b2w+Xpjn1dk5R77Sy4ZZCaGTv5jia4+EfrrU
gtCluDx4/liwVCSMQ7YUU44DQzZBSmRhi+XQBVYxcrYCv/+DGVb3dShhBb0+g4ck6pUWDO+6kYux
j7QOrYn9B1+lcKIp8BO/AZ7pmHZ/+9XkBbCj43t+qow9ONakXPHItdbiGFCmZNNcq2mHuFhv8c9A
/bG7WeAruYdC4hZThvnGMbT/r+ciiIMoyaMsRg00Wn4/ObPZaKhcqn97IYTa5cw5mTn3fgEWDE+K
GCKiaHZ41cD+Z3hqiiXHY/MrYD9OPdV2iqyy+k5o+R0VqHHX9KCQjspLzVc5ozanQyGAwwS1BU9a
RieuvnRBVMoFGjFmVw7bWs2gqA5VEZGlE16aIgpI/gwulXn8WGorLH1wxa3yUgHaLh19FsLwSjFH
dy2JDyaSe3j+IyPl7SXwG2vatHaj86gFZGb8flEda2kStparB8ZFaJVfvP8UjyW8/eyYnWcG4l31
TdX1g+BJV5c8wqcewQSXJV33CZYLhdZsBnIZBib9Fx3cvC3cRVfOpVXbCWhlMeZODrL/JKrTts8+
pl1NlLNRjPccPO+zZQBMRLRtnofzwNPgIVuGsCO1eFiFa+csWhEF3AaU6Q6ad7fYPMlUaReW5Ovx
U72lp1cX5c9AjRHoX1yLHU9jOxDxTKMTeI7v4YmgwKwsNLkprUrRH+O9mb1+EFCSVu9cM23jXAaV
qqh+GCF7UEnLHpkYY35PthvOUrt15qKUw7VlUIjNQLaLl1nyjMOve1ltA6F/19+qj+hxsJo4yNli
jdUQexW4rZn8YaVhoHvF4yGfq8wV4C0KacMXCGdE39ucnm7V90VaiUMdX1RjOR7M9r+icm1nkM3t
kZrkfKraIG0CZDi2kFt/KdOOdvd+INb2XAMdbPQlHIDkGWjIO/MyUHLPp31EkyZlkk1jkz/E0+AZ
rbbQnoFzCtUGeX5LD9tjllCw05SjZJ3DNmq5Eq31k9XvNb1AOoWVCWyi7GIRo3ySEeQChXd5lEDX
d/b20+Qd9tfvJE5mEh+NpSrRCpSjZBfFQlF2uq8nBuqqWzz8QOJ5kDUIiT+yM+da8hFO1fgVEU6C
aZz4vITGOtQ8OBwLVKTgjOhrg3vDKW7EpyRDqR1dVYyoF8XZEjX49B6wqR9RNJS+zIu5TS4VpZCL
OLhjxu21/WrybXD7R9efYcZZb48iGwpQ6oxVCKjMLLFuQe8INsDMX6JIynsKtaVnG/V8brxN5Jbv
yl7KEv11akB5q22QWBjhEJzhk1jndxBVLUuMe5w6QZXJ0Q/hRoDg9IKJYAcvFmpwzvASgJZF3sv7
Ap5kU70A6sUcrLiKDLwy9CG/aYvSyxqAaqm0iPzBjymaYF+mYzFhbfeYqjAHmqgxLvD7wpaX/SOK
pA4NWiFQpPXIkM9me5ZAHcFxEv+6sfxxVGP2/Gd7C7vZlsQfnesZAKqKAfrXHvng3UqhzbqX2iV/
RPmQJ7TvVByKydXWNTtr749QybZhQzDY3+4tOSbCn8p/Sz+BLaQGpLydricNMJ1r797c9pph4LWi
5g9g23bv705CKMPvyiJXaBR1CtsG4uHdZ9PYiFr5wkBIlEv26OTO3SfEvPbjLpkgo0cg2UpA/TjD
N2k2v7C7P2oQqRyfvu5ko3NxdLNjC+N1dRUzT+uDo2tdh4BIAEPFjZp/dI1t+KRbYnizoSfY+Nbr
6o1ESaWiswGvDYift4OiXCzIsGP8UlNFo6mgqPxMmZGPqI2E03xiMXWcqLjVmUhEV5ptOlUQqvJS
XS1ZWu8FKRvuDhPQjzlmzsUMC1k9u4VQNOK9bFtSviv4iqdxwmWoNus2tuESUDroiFd0+g81SRnm
eB4WDIn2yrSUzovyMObCW42K96Ya8MDmkGWAAC7CSFvLY42OvLzCF/bh30echUOq04Aw7xDTwbWD
KHGgPebMXKAFG5BVO3To6QLlWaqZqWCwcDnbyhMX6nqeBPr/qvD1+gFeNwEvGQ6F1dNihzBoZYoy
p33zpzWo502NpTDlq9Co6QZqQTcztxi5sVCpQfO9kPNhnsyDwjhVlpjWCfJR/T0p44yjP7sgvUm7
dEmF4NOt4AT8Ys43Ls3jEuzdTm0JGxvi8hUZ8KX1z0OF0OOIGH6ewk682W8D8r6MLb7Pwu+/K4EM
JF+gvPbKuRT3zgY0hUb2/r1WpIK1f59iJMkFhaIyzNnzSxczD8K18deBbYxoJpnGfRMn0MWzchcT
3K+7dDfGnTuzgspFDFDdTV0zzcNujssGVYKtWPvliBk/8zOFxswOhh5GBJobwdIcngmnbe4fECeW
////KBfTJn1pprpkxM3skoXHaE19hLWQqVdlXGJcm+fw5cQGjTf7QYizmlzEatsb9lSsTgcc4OsG
abVHM/l6BIiytz5mesxQQPV4pWeC7U2aCw0sImYRVoMAnuKdPfasFfQ276IeeGRQ3JcwOXYrju1/
JPOiuTvg7PFWH15CzxpmdQZXeNZAgHBvRVS6obz5Y40psvUuwveySqA2tfJLFDHLSkZOn15Ag6Ia
tRvSMFfg8zuhaW/EUWTyGomfJM+REVqyFZ+fT7YXPoT076AbESdAvA3s1KwXnj2qz83ybeVpetDk
4EvlxsfK+P6mAbye3GnTVwdy3kz8GOQlptXycLo9mMuS7Z0g/QKggD7pes7fr1kgvTQddu/z4mpQ
QOXK6ftZAEonbzhd4wY0ckMrShDwrFWRjtORr1IHXC2I9qqh7YVjXhc3O3B7boCz5Mb4sWDZ5/s4
4XtsRRaGJDdO5zzItXlxIpxf5f2YgVCpw3I7VNpnWlZw+yv2VZ8ZENSXxJptiEtuyB/KFHW8HYG6
SyYe1GAgxkH13e7vqbZu3sMLylm+4L0VUXbifXsulJa5mAPWYp6z8AlHSowu3kOvmLhKS64qJXkv
U3EUSvGamb8zMmeDBDs2G7KI+ypIBaogFuSUtk5R76g3nLz0f9P0dmAKGnwUfAHnUxxhMHbobMqz
qsZ8I8qY/VTIuiOcXceK8+QmCwsZEsgOo1pdG7AkyKJMqiEtgxaODrN5YE5E9pZY9W2viDMBCcYW
XLA7nAGFDmo+zW1Q9PLr2n4ameLB0r8Eq0wPOa4aeMQ4+Jsy76Kyzw7HZyUaVGzdciJziM6hTHUI
2sC4HtwUUNuTBl7z3oOYFR7AHMTh/P+2infdCuo1im0DCaq2bvWrnzM2cZyuhXnWatHMryaKFGgF
TtHExfrfDal6x3iVVEDlTuZBX6b5aMA3EmttpzWejshG9mGxLb2usEk8ddICnyToSTKftEyOQXJM
qtT+u7Ucjsh+xO/bMp4h4h7oXSFsM0Tne4JsfSBjPJO3NEWn5N8NLR+w0gB352Ctfa7HyF08/eL/
z8LcCCX+ETjxHQl1wU1ITvHNMnAMFc95D1x0QqrM8zXUWAdSCCPEpgqGnEobNj9JwCZYdNfnnpxc
jqv4FSo3JA4a04bQZ3OuZuuc9lG979NXj1apeVSq40rhS7YYDZYja8nm54JHyEkklO08OrGDwfTJ
Fjm6wvASgzZn94WU0wHgn2oKNJB2XwgvjIn91ZKB9j2jPEUnlV4afpCDDyAPXRN7sk1yD+Ehm+JZ
MRWsCjReGbk62K+E2g4f1RgIFxPs21kLyJjLI3aPnfNvIJ/00BWdMi6ayUOgkCM7WDzQYwC1dlKH
hDZqy1ZgwkdPRM5dDhc+LkWELhQoRiPu6de7z8k6EswZ5BRu6i+L1sgaYu6aAhXL01XVWt0H5VE1
YqkdNIoT51ydHfxLfWVjciCfD5vitJga0yEK3ox9XMJmdOSyfO4wx+dDTrMmc2ZP+UIGihLup83S
QgKYYkMBKsD8Y6/n5F7mQ3X3Wnf9thaFc3dvAn4MwQLeWaF9iaGMjiyer5eerGXFuS874FPGf+WF
sOLxDoMTJyk3BFI7j279rg+q52dMXNnLb+jh0v+XEozksu3VHKSgaOjI2wuhnMU7RoV8ffhK5qVX
2iS/Cd0sdfgHISbaj1SISn0l793QiFlat8YdDD9PQne2rdyn6rrWYcWCa2kExaYHCArdI5oWpjwz
7CuSx41OAfXTGdeMwWFZN2FF18DWR0aBOn+7S3InHhxMEgaxyiTTTvp2biQH54i24HN0SlXoJdPZ
FDEpp6u6g/vh8cM2D8zYcG/4nuVugrELee/767WiRs/20+dxvyutnBZr+XxrSONMtHSqeVo4oKUt
3kqhk8vfFgMqNIsku7tjHzTEA4L0A17jqm6nf99Bvl9+l1bEBIF6e6pK6fyHunsJ4coaxksmO7fw
41iG7jt1bIqiw/nyoF124Q2MJCKsqvMBlcjyN/5VsEAV3RNPY+hwiiWlCnyAOgPDzE7qPy/hJ33s
F1LX7+p2/jIKB9h43kT1vQHm4hjR5Q204DxFg4t6mKXQsMtvQYkAFTzOkPVVQeWv1CZugW+CRN3d
TRGnEDeaNPnMm/vwk7AM58P8KRCC3uSylZRpDvc3KWyPqzE2dACT6z/KceJFEm4IqrcA2FuVvfcJ
rIVGVEFPJBxyW/XUoWwnV2/HbBRavxnarS+umit+SJLltdEg/Kbnxfku2Y/yobPx6HmVyGrTHlHU
nWuB2vbW1QlLm3zU09RLrf1wRvwOqgx3KrtlaVz3VycQuslCRT9YryjCKWdHI5v3MvP+I5EoKSNv
oEZrqgmBTUlIp2DLm+7A6TTcFBQgVqn1BO7GctPJMSBe3/8FeuKUv7u6X+56aiNB+tDO4OXbYiQ8
CuJ+pkf1XF3nzKNgQcndwflqki18NbaRKLRk1OBzFCqWcTELMAPrstM/E+awbzz/MmsEc4Y1whwm
nisKIdvRrK+G9sjfrDxBK1Qs3JfKoRiRltrhPcy7PyNkXWwH0UKNE3MFpds57GX1j0eANUDgUZEi
Glw/fyr4j5oaYww2oAzYHXtuNMrKQO9oCW6qFqxryc1y+zYM6bEzwAPuXyazX1LKu322Yn4GKDGI
oj4jlcvjEGLVPsvrURGwrrahWJkaJ3b0lA3QdcENSrCSZFWYd9PACVr+1fg66aNuraSnTadu6F0Q
e4ygwp0lIWYz3J65gWQxqKBl6EUsxR8jn+8l69VRPJaAtyhosToUDh7VK3jFO575cszLB2E+tj7n
hULanrlp2n9Bozgz6UmUC+Ivi4/xvOMtUmlEu3cDWWRzcve2HTAw8TRTVRQeVXnUoYV/wEi0Ulzk
aTiDjHMOF6jeI12cP20lKUtYnIha8Ito9od8LfO2wtkdoMfFSMiJXzsyn7BytMdZ5J69gS7MYlos
x5A17c1ajn5A9n/JmE4cRXETuH8x2vhd48YHOAfbZduaAg1UYt1olAcwH/BbGrLHdfGnumlmgz8Y
ck1nTN4szJn4Iyg4GzkDdG27K2jhxoMw5Mz+rJXxOAd6oLc50MrmENAgMjoLmOHvRp0ZcpmP2ecl
n1MjsOqnDduxbVxd358P9MrH++E+eJWxOQbvtvNEXWdgf5eBMr1KJDnKC/tcQ+ncctQH1lBGBGCv
fzZMXqfssNRfVRhMn56Hgu0vXm92L6cj7asyssxO9XWgKGlBe4AJsvoOyifOCHAVKDMgd+ZeQ9BW
vIRX8QQAcjT2XjPBJSiRhMmDxn8Qv2QMbjVYovxXYIAUUmOtP2Niaa2i3ybF8TPhAEJ5ZHQGJGsZ
4TCAwE/wPyovEqyGmZS0UMB/Ib+Z7h3dUgnTIRFt2ZJG7LujjaGGM0V1r5jcXNm7Wwttvw/FCOCg
kseuBbuv36lJcNczHjRxfRVqmsCCTB2J8sfHhf1Ng3OiiEf5zAKWZSZ7IIjRF7c441QFwbYiRlrA
W62faKdVkSrbQ+XWd7+UzbtSt1CAWxG7kVc1/SEVhhFrKPFrlyWyA84RgjtlDEEss/6uCCx/qF6H
jtUBV5zbg6neZqo6E+5A1R2Uze8T/eQeAk0lphpF+f6SRPlsw3Z4IrKOwafTSFuR6Osu4s+J7cOw
Tq9VrTSmYIGyQV+cLrNyJ0w5PAt1VkXqNTGa/4hxt8UNj5ydIlZCMI91fuKr8OrkuIEIGQ6j14XZ
a1Dy5LNWycK653vBXJA3aLOdrAQaLIc6m0M+nUy7yWcGWNvyz5f05BxGa9w8/rxWqbQ0idFidOOp
w5aNeGj+KfGxlprsrJ77mWrO4gw46v6ytd6frFLAipBRmhiGoRx6rN0i4DhSkSTmdqrKFJau3B8c
DzgSTnzFUyDMbpEnIQlRQPbBqOMDKk6spToht4lhJHyLTbn1Yxz3kPOYhySV/d1pvTe0jygJSFdy
ue7pL9oujt7Ko23WROvUV6SPDzUOFmJ7gk+GM+BC6CEVHmQTtOq78RYH0xbnreBND4LfC3h3a0ZP
yWlhz4yr6DhKNiwfTqIAdEB4073SyJOJhETZhj7lx9b5N/BiwWtUt7BpY73Uzb54oRSnbfXF5Gce
ecvwOMHByewZwowaFTmLEwWnZeBg9skJBQ4+IPWMw7Zu6VhCfDnmg0Xhln1wWEAPXYrWeSxhnxHn
hftBZps9VfwvbOausrNmvim7FkjPpc5ozCqvdaGVALoeO+4MqXWihHZZ4Xu4bd2uI4flL+/tPU5Q
o3ylvfk19vjhYDZybma/hCHj2h6pg9+ITyY3XuXxKSrq5Nf/B6XVAXVy8PIZcCkUftjcMxrtNXbp
w3ClvVLFyonSm6oYlCdGPSckTjVVfUzAqXvnuSgfBVhRTLi6NAo4ERCoIrbvZEmLOujULtnwJNDt
zLZ7Sj4WNwNogUst38Tfr0d0AwiU086FBdOQbexQXQlQ4IolKGx8X83abYwm6dmRB/RCGrfx/s5E
VIqBMWwa9yTFUYeVV/5btDQCh03N8jkVhFygkQNVNWwaNjSs4Hz44lvQ5ju3zBjpgmvOxeR8cTjE
zUFYkZC4UpV6meSenP/7fx5xkZuj6bvsNzRH5SF9cpPLmLRomK4MKcwbdlrDlwJWrfaZrKNOs7SV
VLfAVEi4z+A0fJWQT811utZckXs5Y8sQArjfSqFwwF98x7J1DeTJcA8V5sF1bp4A2gtTT0GBMoeo
l3vJYaSwENKK+Uz7qA6D7a+F4+BvWxvUoj2AF5f9oxP0T90rer9qxAt7pD+obzjDr4/S1njIv/Sk
sjU2A4uEYfePDynfkfqHkr5N+igcbhWxf6Iu8V8yLeBmI7jB8eXldvHaCLEDj4CU47VmEfQ/C6jm
ebLwt81RbaEnF6eqxgU0ZDrtBjo94uaAI4Kxy0DGoaY0T3EdMqUDMIjKqFKKNtrMo09rj9zZ1MvU
p/QCkVRzGjQREWvsaongjzGkzyxzHOBuAoBnhkuw88laNy1CXFsjAS3jpivXExs3LAmATmE3jlSD
yH5sxEdbwwawgB1Z6HnwHFk2JSezWdxX50kN2MoONOyoDPBVo88mdKHrvJVf0VhHrqWulvN+eMLJ
96gdlokOu3r+5Xmo58qCTBTnQo2JEu7dLucbQWzDLg7c1B0IKPFDxQMNXBi0Pg2EGTPfzX6IhqGH
AvXkIzp0HkhgLyCEuLGXosQNltYU/ylCBXvq/hMaHh4e+GslU+J4azzYWdJOl34I40iB6tByRwXz
EIs0w8Q5xgKnN/7/ba7cbUN31AiN6es/xbCE/y5qWVYL+iCkROilQmZYV9z/8XUslZjXIHfd2Ai9
bVuhtbmnCB0McpcB3Bj2TY6CgNuC107gMdYaTgePGi42jAOeiUJ8hY7FJWtFQSsQXo8z+shjFG6t
xxBs78xEj+zsIysTWDra2xyMpBEzWhNfeutYl9jY3EWUkDo0gj9FpoaAWkvrkG5gnnIBvBBcqnOR
0gnu67d73QHr8EQ/Lv9l9S89p9qaLNkDhPemfIGFl46Wx6nDBkF1bMgGh7Tdsl4c7LmDsEb/vOTD
HLh3uWfZM2X395EY5Ug8A4I3KcJJw/C8MVlAz2U+sJOFR6nNTwBSboV8YfNSYY94OBoJMEjp3sHl
WNroAs1a0HgVmyvuXSTaHD8Vx2T+mwwg721kVPH7gZM6prH2LaMtPBpXxCqQWmsvwzxGUHspDHDU
GV5zvg6x1FpOV+ruLbb9vjmo12dN4wayZG5UPtK0XG2OmONm3QjtBPxPg8IWF48Vnx1muXCOms7a
yda5Tqh0HwDqTXh8/KjCLajDnUgBaoTxgK80n5mIdUqrTsio/dUB8ZwfZoKJ8WwOa/qWgtxk1iIB
wiR71YElSjMPyC7o6aFnCNeFHsI/fVscCMnkToVnyMno0/YTVAM7c6Sq+oLBluM4imEfKTO5O/Ed
DSp8JK79Q+Ig+i2HFMoKQ3iLmiVLFrvWTDHoPzORxbH2IQeCwamKQUaP5gow12vZLUb9YMgaXuWh
I9KRGpY8lXauWDEkgnyfhkY/cXsSj+3xjBcYL7kimUtG9kmOOQBHgiFJL7h88M09l0KcKFRgTUC2
SXG9aUpp5fSSHUr0iE9QSGzCKjCzuGgiivuHlzF+WfqSsza8UtgHNZY90WOQaxtk+ph9EQt372/e
tEVFTWqmzFfNSfJtj7iRk7PSdjYX5OwGY5oILdYqkQ1Yb0eRbs263ZV/oUN8z+EemK4k6k1ABjsG
Mzx2hpN0UOX4wE1F8tb1aDfbXiIiBr1t66dFad20X1mH0Vt4bQPk+zxwANA+pJl1Aa7MVZvCF68Z
pNC9FmoJss8nCIdrnKq+5KmbmPnMyj26YSa1nGjwaIr6uKLoFN8goHAkC1Bz0jxfqC9E0HX3q16d
6kLvUHD5OPdqlxsiBHL4zzDCG6yDyvdCUa2DCj7yimYdf7nb3zUBxVZTndq3IW+q2h1YoWqB4RZs
PCnHYz+RGAml/eYAIZMavRABVWL4IzEO3utS1AN0G21bdNV+se4Lan7ijPNgOFASMk7iu6XwkuGy
3uHnIDEz7XLs2kCFX6JIDQZYsMu8MWB+XgHkNPDZADN6L/wixMjJol25f/W9Bks5k62wZFCm+K0g
orK3R4afIz/y27sZ2suB5Y3ww1BdnP/kZeG73XfZqnwNECMR6moroAkDE/A0EIaBtPGnGit0W+BI
tw3mrjrrHQaDhTNlUNYliWoLEfvmZktS8OaDuvFXDp2KethXJ7nlp2iA6RNSqpU2ujb4JbynlzL3
bJCEAxF8AgjktFVFjZWBclicmWUHfGmLWHsZkjPkPjJGra5mPbGA0FyNs3hXPNudQwtLji+ZirlO
4J3KLQy538WxmUlPjpFwdYNSflD+o5HeUyi7LtnWsUEKv1V/jSyKF35k65qnSFT8wsiGjDCH1zPP
hKLVuV+yLOliwBzbKQUsSib+RPS91H27U6wTs77/aVL1/0O/mCeL/t+CTU4JX4h555R8GuNa1GAn
KLg6q2iFZmC+YvRc/74Y1yetXUs/kl+z6E/aOS921bfipEufLR4kBPBW55Zwch5CE24fmIIMAzBU
tp2mzVbZqcDZl11lNoDEJqmOoAMVdpvDSQtN+D0NW5J/mX8wuDyrzPAsNOniNh4Xy2Umq77vEzFy
52BMz7ctHYj1OwY5NImT7RyYrM4ueeR/GlrPLqKodDkFiVW3oaf6TCxQPn3LScrMjLhq3x02anlp
vMFI4tE36Eytnw/gKHaEFaWjB6tK+3m5P674lR/+kJrGioMIneTZsTN4MTvQcfg+HOfmYikrffw9
5mlfmo0YzO7Bda9YfSdE3ga7zrZ9ibsAFfeNQtVY3MFF1dXjEVvvtcC9w+Qj8T14R2rev9j3F/df
yTQP7ENrRMih7nZldbruXTss9iUwtJGjAeyvYlwZhHhQRwFARYL2c85EUxEVAQeuNZMTLrLnHMfi
oS9vM4LXad+hF990fTK/zQfmxi3+T7piA4coL8XReE3o7gyyoK/WP4AVFzbS5w3+W9nAie3Hh23n
RXcsEuSowPllO+twNCspUbOVVCy2xJ4vy25YRJTtuV0rS1PCz1Z7jxK/wfNlLJGgwSGi9/veSPpM
o+GtgLzgCJ8XmOqKAG3rzyknfh4QdNJIUrhh//4N68OErLjJ2JLZ1KGxbSWJTmHCJBP5j8Lxrnyu
RcUVtpVftdt0z+IbieL6sYDXOWVTsEJp++q/b1PydOFVRd6HA9Og+nvXShXmnkdM3t21iXx1PeMd
i9oTFo1NXV2IKyxrxVZtmYzv+FGAfb4ru506VB87Wcz8xt3hRQT2h3Zih7UkpEPzMkK3oHnwulTX
nI7drSt5FDENR7sVZP19uKV5TiW8J0BqnM/ourbgNlKQ5eDK4xOC2MF5hrHe6864mKtrIKFohIs/
rKRxVKTGILztUOchffx/pYwm5hXaJIpml5RWgZ+qnt5H00W+/1zVHzEveYG8rEYcHh9yJr915g9o
LHEpRsuOUzqVaajThbd81mlkGvUySS2mBguU8jSQn8O6MR7opbCGjljATSE2JumlNoKvHjYK1Y6E
26eGR/j2rWyoBfRLMY50AOQ/gmPERp4z77Dgm+clHbts9iHhUUNUlLtmIEgtJSZoXZ3ey7ciTp9p
Btua0RTroFWIVJ5qrkRINvYYEjRPm3qXSUd3K1IwRhHVDFG6gzSZnKS/MwAJPbWqwWibB9/+IPjh
XYx7/Vx1S6jem14nswykGjsJnIVKIcstlD2HbvTcyX7kI8hxPeMq3pNojw1jhHYc2sYcT/FId7X/
A7WCg6qeaMM3HIlCIMCQEC7PjbE+Of6D8msdnkF2WhmkS12P5skGLwxNZ8n1vxrwhckNdWghazfw
mxoKjkOaG4oIQWl7tqHkPJo8dqRTUY2WYkNmSpsEVRwpkuWL63dENd86/cBoPZvQNPAC4a5Po9Cb
q+MbPTtcC006h9bSDoTEYGf0h55LElzmv/gCcgKPZvMKhqBYFutOqwCeGrjM7gxR6V9Q1hDdTJTx
Jh5L7tc4izvDjXw44reLcKmgz3yqhoDQBygkwJxLJ79Qk1cu/xs32NJJwFF984HTHOBhpt1n6+nx
5BWcleDLU+c+Rooe09zYexIeKwzIaf68aLzFUBtpXVzr+KIcXYJ/uZTJBQKeZ0WcOlApK/na8rbg
Ik/HhQBvPQYHwp2+9dqJsxaGC9F7ERe6+VrKXYq0GYGI0a0SX1NqKwTDuxDstd79hDGfbR8ht3iA
0FP2soku0qCDz2rTbU6woPDrgrLvmRfTjg8EFPnlFqccubmrYz/45RiJABNL7H/nh1UqRwKc/Ita
joVEbam6DWgJKkGMVUjIj3JMhqjMVgIO37lW8hphEI2fJJZ8px1FPMqk182zyzPY36Fm1Q4qeCDl
/iztdbt9xiZkmqabW8Mx74z32ztHE0KwK2KCCdpgroicJRjpAHSw4SFvA9YBaCyfzqROmuE6kx9I
Nd5FIPfS+4tTcai3Rpdpt/hAL4yEfVJe5kD5g/8mISXIau0Nlufnu9hQBiIf87aoAHf+gltiq4Re
/uQ6i50fkoNETSuqHVifggTUzLOYUDvj5ICvTfHTpBUOndedlQROvz9DIWBwDVPXWN6eo7Af40/a
gcNMcqRg9r7bI0SA3RaXL7wURIQMQkqzR0hBZpHzXligT0+SL8/kOSCmrZCTUrEOz0x9YW/fIluV
prbOJRPJqUa/C1D+d6uQoIyx6vHYiN56DK1NgJ7bGXa3bSbIK1nzVPvoeSeJJCrLTRWpF8nLYl6Z
CTEwu16YXUh1h8RAffp2IzdLC937niV8TWmwrh5Czhy+J/IfoOU2HkVE64EfNnL1+4wuW/orElA1
7uboaaIlAxI0aXDYP3w4V6CJA3KlwWxF4tAYfh5/6doKoYTyiJEKka+hEk9V1aisnjljJbH0r2u9
kpFdhiku/gcrkvNEZE2Y+ADG6GDjYKvUXRou4MY7gCunsVfQnvuxx6CUpU4UVsrICN2don4KY2/3
2Ec/sMbM50iJIB+vLX31c5iIBqSkNdoIUy1HwCNvGpVLKNFKZJpiY2FCZs7/qGwHAtOMRZCyK01K
VCJVvqpXf5qyz4zF0x1S4fRUnIErwOT/UOhmDNF+NRoBVNlxhFZA00S4YX1lj8cGnrE+oAdrOoY0
Su0PGMnHEC7hxSqN19EIBNYpKY7csYe2pklUigMnIoeHgoWdIlza0sHFnTaz7tSzmCkYPtLhxcWl
6Qy59SEHwLW1nyJqkwYUvsmpKih9LJlVJ88m1R5idPrIDydU74Fxep92gBGx+r6x8xM3FmsnirYO
Ujp0Lszv5hDp76c4BII1EM1cqFDsBEYK1FnU45chzQA7ipxYF2wc1CiyzZj/ZDFGBHC+Jg49GdS5
paxTB9xRQZcZ935WwDTfC/84ECWlaNtDKK1Zh9ASwY0nwIDJ7U9p4UGAAuo04Ymd79ImG1mw0jk4
Fpm46cic4PdY/7zgK8dHdjajfIp6lZbgKy7prmkdoppSuNZiMT0AzjkR2QtmM73XAy5NTUingZ/W
jtxlwFaAn0Ff/X0YtdAtb1KGAcLItPgG1FbVTx5/XJybCGLwpHDZ/JX/dxOLyJyqyhHJNqMptzHo
D/TgcU6j4fKaZktrWhC3KVC1ZbUIETMCWKhh22h3lqsRn8UT0jBMlkm4XcABk5uX1q/PEB64ScIX
bq3BBmEFseH5F2PXwf+2tE+u1TE6Y7iuAuCUyKh0QHOElgY3L1RhWblJUngiJPdAc/VkT25B9oFI
Wdgk31LGRBYLfzO/BCjR4scD5V+w3Ub0fZW7PFJn4tfsGmcYl8Aa5WOpkyiJJ1F8Lh7WTD8B/ox6
i+pUObtDEouVgGGP2W72dxTtL89NLJGDSavstDgFHyZSeWyFTDe6QAzGYJR+0k9uGiQg8HfEwPpI
REe0QCn+xmGl71PuFJTOtG4WFcymEF6BU5AQRVAt92GoP53r9ORmymbuuC04k8tRwTaJcfGIGgqZ
zfBbqAfOFCXnrUMcCvkmjcjGO1gJmm7ztWwzRCIxbqdGnCG3a42QFY1f65OFY7KF8/zjitD87uCK
G7FYga9lO8K+/F6TKk8fTA/HAJCG1i9WuNvRVoCmg6MBTW9lWRFOltBZ0GZhZUuN2NjA2o8xM8mt
NwLiwqaiyaRHEMpDTe28rfXxxLPaCt14smQ+B2L6f5P/kPsRzcnWFRdhFCeQsyM4fr6k0LqoZ4Tn
sJcNS3gu3MUwjlqAkds0P5s4Ne4yNwfRj60LYnqlY7Uzj8wbU+tYdKLgVQDbCaKXCNYx3+68gAU8
7YJzGiYfLWSyLrMTS98PvGG3qfh2R+paBHQfUk9Zs3Mnv/5yQqFaT16Cinud3WmrAQVFuwkcOgWi
CBfWaRj3Tadbk8yLdzbUjGFtI9J/dOTM7BYohPJIqJYywx8BiL9yYXpO2GuM5w+1jzGNcbxbfv8m
WiD1a0UfjlISW2BoZs0aA9EMJ+t7V+Vzs+xTevDV3aMfhipSL41KLq9FXaUt7p1tzpRjUp/Ui6O4
5pxUityeMEJTDhh+0cJT9ezW8Rgb4aVjdIj0u6/k2FCM1hwMKsOBAVJpJnGSyMDLzGE9n7V4O8FH
Z0rC8jQxaAug5CJn3I07qQ3pf4SrySP2H0laW2wVr5w6W3sKDfKIgeN3ed4HB02/l4KcfLw59EsU
oPrmT+zVuCvqI2dm2nBWCu+fdqxkx81tgrrWl/9wHKQSFR21J7hFfV6Tc8YgZGd0H6XGpubReKL1
IdgFpmRkymmO7I/EzChUhBgl2v7PlETretCxeggIYaOYtd9B+HpSUm5jZEseHc8Rp6FbXtg50OFs
X0/I4OxLDUo9FtGVqglolit/vIkjkWWZ01p5AiG1ef4eo+PV7aipC22TO23eN7WUtFLBYuGC8vHX
9UZXuShYSwtjwkHZ+2sqd3I3TJSP6F0SFyZT1yev5Gafm5hJIx86aj6awmUUTMqwas67KQo3Ww1W
iyCAq3QYEedjK8qBq2ejyA0nucqrwMgkXx38xpriqmEKWz5IdEZIpZHA1Z2xIlJgScjNbn9B9Z9m
oPhg2VT2S0eMMYNp3RF1WTwp1B/hp5AtytDbpY9OgFQZLcYo3MpbyZKDUFObjXG55azS0IeYM7ri
12qL1QsDNthjMP3e1YzKdzOy5V1MIciKMozP7DXshWWD3vACKDHqNRSr2goGMuBAsp8B1z+k0732
hu952KQyU2j6fe7O+0lgibG5CZQWlT1P5CqDQXLrkBvXS9q7fS9yMMy676DIzRMBwZJv9pn1Ev37
zhsOrBX6Mlo/fxdlnQ1lAo5R1Kew6Afb3A+e74MZTQCWl/ZN+wMJ9/R6xJAYxMMoccoyj2CNyvcd
9LV7Cp2hyJYm2X6w4SKybGJhOs2kESoEPZgM+7q9UOeqlsuIhzFfsjMC0aPQSJELFfCyCfAaNbnl
crCq3wSNF8yP7rPR/wUPDDLA69LRNgIgtMC3MPGUGlAlmEuFOQqmgbnw+7iPhhWkP1ZCNt//8O7v
hVbXX8A74IRbgzfSN+Dz3ynFAMJiOuGVqSxcyxi9+1AJb7wRH7V/x0JvmXTN4lg/b2UMp6pUmOA1
wgFjm51F5rlcr+w5X0Cao4sOfFQi3iENNYowP1MCpv5SY5xhKvkZ+uTbLvoDNWE41VC7LJR7PKzC
r+TCOjzlq1Qjch+E+uXd0wlIOu9d+TE5w41l/ME2FX+k/itSRQf57jsbFG08NeeQ2yZ0pEikaOoP
9P4QUCeIkiH0SReyz1uBXMzM/m/6ZyQJYcf50epdZL+u1d9HZOU5B29RMAs42+YRc10aVclbwdmG
yJVtp1CVEM8RSyAem13KQETVLRflqiDE/A8UpKWU9DWFAKWWVqeyt8aw72r2rd22Z9n1brK49+wk
xhVSLpwT61as0W0vvFZS3//DMh53ls6fNw+CDVH/mAzEp3X5MFCLg50n2Mhk5mXM3KGT02XUSbgz
sOyeBfxnqgh/DuW+ZJEorqRM+zlHU5WoSVo8sET+7EPId7a3Nv7Apv1TcGt7SaTEFIeVF2ZvIpep
5/W1px9NjU3z79R7GA3Mx0LWPPTq9zEzBZXha0o97YlMcENePj9ywT6FpWp6GJFO7A78KweVLYIx
f62yN6v+NruZwkv4oRyAbMIM2kss1sOTHyzvbfHllRt0sBrql5YFgpnD3iVuYpXVoVM9+EmGqXE5
sbYSEXhoQYmsYJo+ElkEkZRjGY6DYnzW8rMkZGLrSKHdjiZ9lqCJuOqo4Ly8Z1lKWGHxQxr3BfFe
LH2jENZPai8G5HF9pPumVmpwo2i85YTsgd4Mr0Kx7vDkmqs6ON9Tq3aPnuTIHqrOKKp+GMnCKbzV
ZlRyyZiPvI4lpiEUB8q4DnrCqPatr5Fmx77/GIpgZK1oeR7c28PQQXPCW4pakcGfbWwW89DaFOlB
Bh3VrA8jOHUrWheaLFZAFFWkk8JDJ4zEZEcyzuaIn+uZSEzolvOMN06hYwMVGMtmvzNTuSGaozZu
kuTPrjw2fDqt1LBzeUOSIcZE94blwDcCmgfxX6mEhgYQbu4ciuef1R8yK/u1ToOz883eZO3gzt0v
eFqhYrlEA+kaTYAtwFs+azxN8qgFgRmAHL9aqzuzQelH66El0/M2/EanBYMEBKU4R7dYeZJY0ixT
5eSEUc3kJmhtpJs7ahUR/UhJMp5DZY+E5w01tznop8Hp8juDdPIoy8Mlwy4bm4KuZnSx3HBxhYXZ
lv1Q9bViG/ovbOM8IyXPnu5rK/ICjl6OsX6y6GTCWKrQLi43QcvVS0S6cZMHx/BHzAWaaQnvB9eu
qMYQZyFAYfKhH2FcD3BpvCTnDTgV3EVOfEzePcvDw0v/A7AKBIBy14CeIXC8C6kuY1wNgiukOSGu
qBgOMB17y23tQvtO7pILDL/hU6SHede3BPjW9h4q7arBVIpLgJs7r++j9BJ5BnfErHm1IEN+GSK4
war97/oF6L5Q6ArdoJRjRgGP1P3Bv4nm6VcTzKclEMAGCRZAxTpuI53yLB7tkgpWMZ4Pd7X3smyN
4jalJUFcIO6Z4ZMhwKafokbONnwjpCXsq9QDWA9/bbdSR9Up70Mo0/9zUX9Kc/NKutjuzjkesNp/
JjbNgQNE55dfFKM3zih++/jAvTttFpAqAnLs1AGcojNdcKdHC5vWfChWs6KIKiPniV6WbZXF+Bgb
s3IYwrNRAKZCZ+kTDv4f9O9sDe4miCjXwngZTbGnLjtLGZ0agRRf6SyNYWDvy/DWA1aHoX++v6+q
ox4/4Jp9uDLSejRuPYSiCrbYQV1X77jEpj4mNmUd5ZXfA8WpP0AmRp4MWGObRM4migK3JhA9sZzL
F2sp7ezyvcr50EealrYtMC8kvOz07BWgwNCnQHbknYoOrKp/+pN7uGYUFw4a+XFTnrJdgyK8pvS0
cpLVXUtF4BMBuXpDzZGcYry2xvjpEQ4vDDQhRrUW4UojXvW4U2gJpoFswsqx+t0I1yY8NUxiPWC4
VZxLvXnpRLpcE0PTfiA91k5INLyLDmOs6SpoE/GQf7CwzSSowDIxKvvjFzlTLK3NgOIFoQyI47dO
zArCBrhixFqbrnX3I7/jR/MWD69kSb1QHE38r4t9VJqoKIX/aN01409PzSVckO6A7fybzdcjKQjZ
nW8TwP8h2tkE9MKcfZDKPwE61mujjxuUxRe0R9IFUzO1LbUDK3xnbkpFcGnCg07zCH/qBegAS+7b
U5twxQtz+18XQDqZPpI3BS2w29hTMZWORAZIpn0cdQGu4mtCTCAaN0aO3ypp9rbJRHbOUmFWbF2F
eo7e3iQDFRPfFaQrSU94ibUFkPvq7/nd+nrUsdd2xRogU8lAgoldVQJXGykz9ezK0ExR7zF0QKN3
iEe44s4NXqqoy9kQ2JNEpS+NQDn1swy0F/sG8qGVUUoRv4+c0G5A8CAzfw4eD+STF2cYAnFVsrf/
WQudpVcaVldDy2iomSFdCClJgJ+P7QTIKH2wfXrXXxW3XEJKcZy8JLTobJMTQSHrGrCTDsq+Ot2V
Gv2+hHjznDGpyfW0cNuD8Wqkb3jCvWYXlpAzGUR+3q0dXx8D6EAXQSDODWf0oF3l/DK8WqlZp4WE
1Cplc+plw5ShT0qghrCgZgcEB7JZks1nCAtq0Iok0g44jYlXNnbm3BGHY8vTIF+EnNDQVF8xL1Ye
2W9dVHTE3aoV7IlHsIPPKZkAhGQADD1N0fYfJURiPqBSEguJIuOhZ47a8I53j7IrbAgRDrrg7JPf
UiJhdlJ1IWB8G4vljpseEUCdJ4aWaY0LeVS4xXqYZDKaIwnPSjUzhbxyse0Cds774OzkrIqt2xhQ
CSlyyWPy/g9/y3qYGuKJAyuSA3Zn7QZZFeiUo1Bu0ayDrLOK0RkB06LY1c6bHIjnbUQg1R4+c0O9
eannGzzmSL/Af7xv4o/dc98lLBM90Q1AeSh0jJ5nezTvw+fmmuSCllHrSHc9KD5F89KrrPNCnNAy
YDM3CoxLT2JG58rj66cdXuG/U8pMDU7QeoKamMOb50JiXNfTZuQ2NCoYe7SDwCP7T40RX7GvvTSr
Ofg6KEPKSjanG1UYMRY/reVp0zeEHlhS70xrDm//RRwFi17JftlBWkzfq6l0C9P90xPym9l37nG3
Qk7XOqJxDKTGo0fNm+7PsQ9rkYWJoUgndH93xr9bT//KxLOdJhyHQwWmk6wAMpLjYNGmY5fIkWzH
LjH5suD6n13eF+QcQu3WjJpoqkcrjNDLIttxSKJ8iexiYQYNep5vX+2AtXRbyYB4t/j9IkjMYdIW
mQbLPJfdjgaVqpttXsDkF/reve/MM/tHOwWMoaFr9HsZ9yejNbWbrWFMlUVV8corvx5DxMDRVXin
/7HDZYPSs4CMJn20EE4jZJrvE5Z1Ion0nYRx7LwnY94P2Iy0fUemfNGhd15n8lYGqOE4kAtm7mfD
QphslTA8iINA5TxZ1zMp/Qa4l+QWBXKmPZkzluou64uhJ/3CT31lELOPvSpKnp4gCehhlDY1Kdnf
akoEyhlhbe+AqrUcA8EnigF7E6bhTp+tyG2eHUPsO4IOIzcq+RwR7qB8e+e2DLYYbnxDIaUQC02+
YL9t14Re9C5cJ59TfsGV5widxHOtH65DGWXP8Kk2WsL4ytzFSqTcQ5weduBIkJoBFV0jVeBhhRoA
+AdofbM/8hALpMhdemQCCyNk6qwjahxmi4Ld3Rop+LUVrrseaJpuVnnyekKyYm+9J5XhidpNuPCt
nL6Ta+YzXZmK+njOxiwZRRJORV18fvifwUfKFN0Zr+lPeARbcL4GZiFGIzagVN/WFoHWohoGQjtZ
zDz3Wt/59jAyke5HVshw5JLBzjLeRDH+iQATIuCMWytGfQKI2xyOJaV/RVlSBSXISLjwL39r0DdW
6EV1v+M56lM0m2rEVrH0GI/DtsjIUrMhdNc5V4uJmHgmQ4JhYgGSM/a5IIqxnFfFH3ldllyxTKag
m3+ZFQziU9UtpfGdS90S+6NeRgziHJS0KsrFdUDHfziouza2+SjWmGl/I0g0a74a17/EOrfBx3F8
Br3YQjs50FVjThIUWGWCOD3Rh0bbo3zNtprnuqBmFrZztgL/uHAvg6rYmxjpr8W8rwDpaBL8Nklt
1Zi19E8QDjzQMnwt14hJ1qCG+7qtQTbflVvJEuSUH+Wn5NacFae0CL2m6SsTr6XIiIYGKWmsrVM2
tiZsjRWw7K0lJUAU7b7wv+1/w+4Vsbfjyln1aE/WjczX8ieQz+VZgh/YobXYgQkOfM/5Fln5cUQ6
F9lHpPoNVeFgkSO4lRA+i3rpVM6zT9txCfwfM4lPwinsNjeEOqESbC0vgeLv+EVWkAcEiFbUutye
FKZmbtfclOtQsZWtRXK/eEMl65NelO7ertWBzFCsuC9Z0N0N7qsVSq0gRsWMrfjdOMbDycL4do9T
TwODSgWEwOjMlVnLGsm90ZKncbp252UMNBlpTmwSeYAFasf+3AoODYzLRxgZO44Oh/WAviG2Wzf2
Gr62zWMbR4zvGfbbx6c57+DPzWCIKEsUwxBDXa2Q6/OVVQBkjCaf2T0KQlfJcRR0nsXMhH/vYP0+
JMjO4lnap6eEa6yrDSZqtV53HuJd6wRlFe2Sfx0W0OaV4g1XQCD8sC5zZCtFXuO0CJAZCxy1VfMw
d6aHsAKmBrJjR3CsLnrFKVqts7wOuf0H9w8ZXDFAbiiBsXhsdySAe86wf5Shr1NrrKFy2KZRKlJN
wYOjrnQyNzESWzTfnAcjnO6qXg4f1jRg7o7sBjJurz/A222V4rXb2qIvkh1h7dqaMUoYYnCTyQ4V
s171Ocv3tFeonhfyLl7WMbrjz0tuAVjqbVf0+OUiJQL+T2BXEiKULP1h4oSZ7InRLqLtuCq+7w8P
nc18mptlGig9LgCzKYXW6/Vm0fq7QIZ3pRjmJeVSNfJAsPfP2EQNO5vL2BgiU5Xym9qq/IKi68SV
fPBZoV7diFxYu92Jdnk0sZjpNdsMji+T7CPT0Xmkw4U1oh0+YLhgVLTfdIbK2UWUSTAc/O6dkovU
gA6sBFK06RVwoKHK3Kn9/8VrBsy9p3tPvtJPbSbzcw4OrnOnZzwiby0i0WGh7b9KFa/Fj2OUSs9z
BWuJEMGsF+4qFd3LcnSXOHG2IDxFtovYMU3XbqYsU6h3pFP4xVMcpbZ/69O2NXIFjiYdwQ240hk/
Bu4EQ4C42xJSAauPPaf8gowmq5uI+CD3qkk1pa6XUO3ImU8Wwv1I8tBAcQSb1QqFXsin6dIWVvoI
byKSH31IPsLTlZBf+gXDcg7PhbKo9NUc/VFN7w38kdMBSV3UMVpJux3c09e1GEZTJFONfRvpt8BE
/GHQBxTJic53lly3gQCgkxs3GSh++W124Ry6UhitL1SYTeO+CqPBjn/22IeZ8mFnXrz3EjSjEC5n
4PGCnWhLhOt693bfdvCjUSkK26F7AxF/XfCt5cH6kfBCXgAruUy7gZIBUys6Mdc8+myH1aAWs0O4
S3BQ22SduGSn9g4CwW2X25ulLXtG2BACFOKkcH/AdI1RIv9YkfaR/0nwqCRc32wdxn5r5guWX3KZ
Dz729HHjfxvR8qLpEDSC6KJl+DHCUk44wGjA4t8vuMIpNb7KPWatvciW8ujZrzCUU0sO+suL0Qyp
3uIav5TtKLoRJdHqn1RHML4Zty3zWUVO3mB3mXkUmH8PtX8f367aWihHDXivdmG53+Cjeqckzkvq
wZL7h+x8shDW3jnxHxKagUzxmMiDUtmNe/3fnXCgHMqSeYumsJrSqp/UR4mezEAjgXapE9swgCyX
fyCqVaDqdMhXDL0RI9OzbdnijYDu/NjMlBhvF4+tYNfxd3Rdld7dHWToYZw5HWTs9zXhbWwD4cF9
OVH57NlPX7tSDFGzBtWZ5Hjg1jIhAxPZomLlmy5qXzVfLEzLOlqlT1ra6bNW1N2j+AhVnk0XcV1P
aM9uyLpSpq9txjF7xu1IiAmCwfx85lGlIg3j6y3RXU/hWkcr8vyv5DF5RgO69J++9AKwUtTkgY8I
gfPLA1uNcQY2r0Ru2Qo20zw9hyXFEakhdIw2bOfu624IgKWUYbgvX1SykGLIcbHHABNZX9YzWzLm
PZzWIDzBbQYLp2f6k4KoV8IIv90K5FiwPzn4qY/AF5zPReo8zFAwdFAwsI+wCtW51/CMZeisV7Xh
0pobi8uh7ioXWFbz89coWiDG+lYUbVD9eP3P9jNkc8r4JrykMtEax614PC4wxKCvGMlQG7BI+sVj
ue5RK/+BmeL25tGB+d/elXc8T9favCaXLbFuB4InI8YzB0py8wAidws9xHxK5BB7n2Y74E+g8Lit
/PNO11toxmMo4IUUtdXkYd2vA3kgNUCluqunofAG6c1MyGrKRPgtVqc0afgv6m4AMnYwdQLhiHGH
DBzSytX7e3tELL4/20bC4L1qTv+OwAoaGT4ew5qoasxHc1wMoaCFBonj4jXfCCh1vqenlz7Q5LbF
RV45W6e4hZbCrZiF3Ol8NNLMXpVTT7CZga10JGuk7ctBuqjf1D2tOb3JmM5L6RfIrATcJzbY+wn4
RyvAitmd1SD9xvC5SexwxcV4cFf6Ae0pSmxRseVE+et8Jc61LwW1APUAN3FUt2434LWfdc2mb6Bv
r/9SK3Vq86b2oKSqLuWCnbeFH5UCIjUpLylGLlVEvE/MFk6qssYcfTnDc8YRyN4szl0aZ7ueD8XM
WgwDRxhyUOfMJ35NR2lSb3VxciUUogG6b8nEwgxWfW8BFMklW2SrEhQVfOJy8/wU4STnZdnTfSt6
EY7m7X27lhpJCE7Ks1cBW7eIIBt6WcIpVJhWS6vfIjUdX8dE7IfQ1/mly/kv7X1dfx33rz2U8R4P
ZVQqSFIBWvnS3dj3ZcTvWUxbKDrADuFP8tBRN8lTSv5+IoNuChAgi+25r0GvQAZJQwV2clILk2MO
RxMZPhO73lraDrjKmu7ssZNHD/68HyXoCOTlV22ZA+b+tf52v6dUk0QT2CfSVXT/B5wa7cM9M7GZ
PfoB2hsSWLgE81AhsQegXl9Tmk7jQd3mxh+fc8spPcs7kodcWJqYWtQpDke/Uj1//vurkbXp0mQ7
Tnb+QvZuQW9IQGhGFQvdkdjTpsVVRylY9CM2ESoOQ26JxukZMuPnqKUOhKzoRNAOtG+1BHA7efEB
CpidPlr5FM59hsawiGtkccw+50E8ob4U1tM7CcM5IxqzVi8s24fXndVmf0v/7W48QaMw+1Mo5W0u
usP+jkIzmf1jCT2Tt5p+lSr6pDOLrORQ+WvTxok567I2zkyRk+USKMH8UVErjaqA5QKHhHB4ZlaV
BBL8TmnM8XG1DAkcfAoZptVFZb7snhV2aeZk5oaBA82WB2uMDHWBmzduXoUn4V7taN7ZfvjemwOF
QQsMMqsDK04+/yb6tefRBOErdybjR2KAuC2lIpGyF7qUy14K72VdGUN4pGmWYGB4TnCaSghHB0mf
tNrKxvjJRkzUUNfG1B338kfeAYVxu+J4s8NrkkXsdt2cSoVl/QvnM8mREmqCkkSkhk1e+xPplj4R
xjaiXTcMyhqrY/ZTVZVHjl4tOhZHn7iRi5gmLJoe6oFBPnSIMDluoyt7LmCxoftWvqVTJAGvXLvw
+qWjGBLEijiOV12F6xDhqn5ppBQSAJXUGEF8aQa5cPSGd9oOax2W/e7dilrjpHWn4VPaUbHP3aZI
AQctwaAQkS7m1yXg3ansCKvXuteyNpZVTKy+HNipA0oNm6Zxp0r7Wq3a0a/90ZVebITiXBs9NSQ2
kuOSOCU/zLq9Tmy2plWifCKT7gissidBnoL0TXUOd6y2nOKZR3siAH6WluffNUu1i0iiRuLJhm9d
LK4t+UgVKKC6aMj42zod8jnpH2qb321qyyXFRGM4E01XFedlcjL5r/3FucwUWaBeNnq8037K4tSH
dqHcrhPY5ENEdz7K2OGAcFZxRjYmDU0qBzpHKcsF/BzgtD87M4CeM4M5mXfCbPKv05n9r4sKLP7U
GKYJykxg3xI7lydoOSaUvkNbpTRI959oGKk8wuZ8gWzUbQGW5+/r5+Ytf084BHY5qEFGUVK3lGbI
Dk+6Wavci0tvDyT3d00f+TOrZkBS1ugKb0YsOQZGFDznKGKRF4lC+rYxBw3xhw7V9i9ATb74FHrp
/q1QeADvpU6XapJc6EY8D8MnWyzOOckrgztZ15GDFMUe716RW/yeoZoob2pmdofpLaVcgl2Y7Q1Q
4mZURHxEGoO3+xEyNB6Tso+qKBIBOVl2Thz8LR3PieSO3B5uJnQRz8betYEgalCPOLNcHOS7Zyz0
pxHcGZUtCvBI78mts9xjmvS0E6g71EZ1zc8EoA/p6a0mr3fSyZCl7qdlGf7zgcZ7nbRm7g0AJrV1
6Pua2ZSLLQs8ADAYoRzC/K66dXqObHDjW77E3pnZdHrfLvR1MdFBeaOSQaaeglO59bUPX6G396Ct
EO/oDS+MF05yWvn3bAvOj8J4A77goTo61DzO9/KaOT4hY9HE6ylF8R71zHa7YOiTy2GcLCh+ak4Q
uCDTeH2I/t3NKktgMqDAXdLK6HPGAFxTvNlc/MoMWvlSHTtv1BoAyGFPNficCYpxzFZRLDxrdTVp
f7GCqHLi+x4GJT3YMiIBbHDNy95jv4SYZQBaLLmtPEEs7QPGgo/tXBrN5j9MVeFlJqPxFzdRUXA9
8DUOOaROwszbCj7CNEwEELGFLHXzGobSha8+8m2EVwkWHlNoGi0/ladwNe1u1mIfLxwv1zXXnlfM
ik+DjjAuWNesj8bG6UjQsLt/2G8d5qPZVxfsnf9nErBr9NAv7I4KkRfgWTsc+9QoH75pk0909O44
JZ26V0HZlls2PiZezAtG1nBqhmPjRKfAWoI7ow3xJyeFilFbSs4SNFjGtalepI3ElIkEi3Gz7c2a
ymhX5kSIdGlQMJdD1f+zPf6QaTasnVKTvBbDD9mjgIvQQIhbt/zmUpay1a+wK9y0h/jslfPpqbMk
b97YgmodWcZzy8fLx5R+X8omLIFFWAHOaN3STOLVkgkIhozaG9J6HtQcPzzvhhky6IW3XpvF2nEt
mY07fzAYhQpbFlk45icu0oxppxWd5xLoIZ5eMBA9TNYzgY9xmklU1lym17+6aeKKrh03oxhv19e+
qMPT3EnAPjiWLR0kbPEKZEwtPazMg9rUQLCZs4ed2j75wsZtNkSj22Af84SZkf/sl31lIeDVTXrO
7pAzd8/x1GDQFeH8gK2M5JXzeGcXMOuOK8rcNCdw7QwzdOSmFQf39lTSSHckjRZhWdF8sE7LupsZ
5H0c4W7YcWM+Tqu26nu+mDhGtIbwrK0wYXPqFJO1ktJIfXQLVAEU34r/KmrM6WV+OhUo535pyVmg
Liz2f5z3S0x5F9Z9ew4Kfm7+pRMGq+m7XHaOUJkuMkO96/5gqeTApWH2oqJPsUE4qz7iXggGhRuL
In0fybxqI62Xy5zAqDw5gohFStpOZEXqIf9ozmF6ihCFV1IsDAAehB6+5RR0W8mhMHmPXop6v0mO
iMUvKX88Mwe4OKKovu3xbYByn9MVeBQiMtUu1KeA6UJvRMUF1Y1VP1ada91iqJOYut3I9ZdxrjSU
yV3MXpPqUgf3w33xPpkEMQxT8LV/D/RhZpR0jpUHD8hzPezZbz0f34X0TVmsSxUoog6IlFBj6QTo
dAE3C7LCvgqamuODsmIEOVOjVOu09szDztqXGbWlVNKmg+YRjYqEyUaIJ2HoBMPHoeDNR9UTLJr3
Try4zj0uG6AsmMr+ZE/V86c4YDux2Mtzvght8VzCmcuXMgjjFVIUy4+KBNgUj+Y70BTLLM0D+u1+
TSoAw9MMv7Ajosm1dTDronNiU17pOZnrxDl8huGEmmedPm+VlrXfM+Y+izOqGjzcYXXzcvb9r5P1
FmtJ7+ExbL0oEV0VZ7DIRcxCYVZQl3hqBvPn4vmsspRpHNLCC1Sh4iPIhmL+zti2dzL6c9DiHEDa
2ZII+4KBE4lDomke6bQBP3wvNb3d2CZV4VCUzGc58RWX++YBT0f18W5tzWrkZrftYXWT+WbmCOQL
Ky/FTjOF2xbeeLJ1/zRwcVfq90KN5fc3rzQ69HMRGsdPFXappR6FVPJYAmgmQQfG9S2OWd7MfU1C
pJByph56U1yOBlp9CuTBmbmsrgwupOowb0p5S/h1zuJkflz0WuCM+BQoyqz53fP8IQP/F5IheAqm
eecF89u2ncDuqhoceEI6OZf9blIspJ/J8IrkLb9t1kFRNMhERSU6nh2gX+0fFi5aaZMcmYB07Ty9
DJI0IU+UxV2wMaIi56GmQeBdrAmi7+7/yBWMHPDRkDIgufEPvE4CVU8CTsCcuQ3ZsRjOkoFP+5Hk
/ucfY5fvgjPuXM1LoOKwr/KFiUTA3/Le1qYVkTYrCvqfIusoz7QA8bJFFM2F4B1nCGi0uddWrYrE
ng5tGsAMjyQND9f8SRJZfZpXcvFY4BroSgeZP29WEX6ixbNkfsmaS5joZNfVQ2U2Yt0bC+P1/pF+
o5UAg4WLvIKxlOuXZa18AGtYsoT35O8yKh/iRQRUEnqLCixubNyd76/2KTKcAdXNlk42mwMU4mOf
TNcGFofAfvhYNhhbCNoNRi8jmjL/uFCsi4a07jdb/JuJ+2PF6rUHn4ZxVn1Nea8PGH4O5WYJMEw0
4mHfalrskl8QNELcog8/R4ZPPna7MSvNmNDF8VerVlHqZ4aDiGPwUFBnLtLZBCzDSKnp9SY8Xrp8
AiBFXBy0JdOwC7i4qRk9xb9qDHROVkqtMYvBb/BYlhDh7j7IMq6tkCTLQZPR1lkrj0pzmQMnQPC1
24WiLrH852ltIds3izafgKLMT09TFqiIEVhyop+QAcSW5wdj2txwo0XpfPnwUTlTOHI9uH8CjsnX
vGmm9rnmL8xFEpDafoFfNHqYilUF123IU/zD0fqYwOONIH8H8msJv27fGpjlUWWe4IY8qPgyeTSu
naCah5Qq2EIyQdGoBmtr6o8DHCleJt0kqBzyDXkKDQnzKl6AURdEqQSA3NeICa8ZZFo1/3H2K60M
7jcJ3PPiRMOIJWfW/nZbezsFqkGjFqDet2pM5ZJfHnfItBo+hboUDr9j2UImsih9la/Hvhy50kYV
Wp8XY9jPupxD2hWQpMpsHAubG0dL+2wJqTnh4/2IBaVCa2/evRlKI/hWEsl3xfv1ua0dhjCXHzFR
oWwYpr7BxASXJ41+jgLJ8l1XfYgJCdnO9eK6oL0rqbLezL3UjAKVn3R4fsDBSocwPt/OHTAFb/Q8
lp7OMK9Y0KMJFUdZ0Z8PDRHtV5wUtFXq2Ks8fx2pm7wdFSTAKTWD4Dojqwi4JygbgxEuO9TEzRlj
xaVvNEILOOULDywR9Hzaoy/3zikwwplHjLi18QdUmvIO25SyVKv1hlGKVagqzGBQ23iE8GzpaiFo
7P0dU/wYAwqZfbb48D0OJ1XXn9/K/lfeoZ6NonNYqh9W8ec6jyJGXr+xnABfRmoXcmg7vLGjChh/
XbJuMl8nSpfvWldYDRjNX6+ZVS3hXvBCNpRU0Z1zkVRoDHdVv58DRX36x/NaznSECO1cJuD/QTW7
wN/xV/MOBLRmjtzdSHSy4pxnHxgg9rLvbG1+q9u0za4QQljB9qdD4+JvhW9dTXGiW0iW9D8S1anM
lyhN5cu7IaVpCCKX1ybqB6Ds9SL11KUCOa85A1i3agGEUOe4fJcbHA3/d/oRbdRkhJMFFz6V9v4r
wUQhWABmSQwvqzDDxpuNQcqpZHK2Y9nTr6fIpj10v/m7NG5g8VIH/XHhpDlewHN50v0GCb7mcoh8
GHMXBaka5gce4vn6w9v8scDwDb4GeRFIiVJFcoYdWrEAIrQj8EOgA1fG9xDntvSXu9xnMhvG67mz
EVzPZfFT9x+XhRN9wyZYJJq24P7nLi9861LdYCHnXwd3oLzXsUkZhZy62B5GBEtckuZJPJUlTYcn
TQAne84WgN5jFpi/5eIDNjGfUvyF10ynDCrlQNcg//VDJTcCPknt74SDnwWmwy0MU1BGSxAItMzl
7og2Qxf1BXuN3S+yiqXbeiKHivVf/zU75w+kiteO7CVk7TNmfpJp6Rc8AwRX9fVOnU5gXbUgWfVG
iv28TSYxQKHICk/ZifKqYM4XFnB24AyDOy+ablXLIu18lfowjoJblBTA+F7CY/D5FW684Fyd+wNE
DLBo1vgsW2PI+gZIVIJzhC+rUlXvaNFbj/AoDy7zdWgRcj4UH/H6pb0qujii4PJeLGkGFv2QJ2+B
CkQxzFEgZqnDLd3ife+xiFPcNsOm3p+jqTUox+GQbajTnjHXIS3MoqkQGZ7hqC2/PRVL9ujq+Pxm
aEANr9AM7AMh1cTNaASMIm4pey+UEJlrNlNn7dPz9mOogrccjOqF3toZ7OLd+++BX6SpH2+Tc7aj
lY5djJEPoQ3m8cWPP9wmdZ0ryWSL5QuwtVnzFHIt6PHSYt0bh7OvlWuPVetV7rBR377C3Dl/8QRA
p00bfr1XafTA2FXRdBcFQ+SGhhV6dm2MANYH/3C88/Mv0MD4Ib+///AiOyTGqkBZg3Eew0EiaSyr
R5PA6uVA2aoXkA7hZLpNV67RnlucIRceZ7ZTdr4bq5C9VOQxfhkYcHGyNBDuTuKwRyJ3ApUHweOA
CtnsMPn9cV78ew/ixOn9GlLJ1qzNs3t13lcFYgrJlE55D7KOp8L7jM9C4pC1wjABJGwOqkGKgCRH
mj29xJfs7D24J3DT4jyrnwVhiC9uSfYaA4T/bJaoiBXRl43mMFxcowkwq7Y6nQB/JFSVoMDpgS8T
LaVa94SzUl45Dxc/w4mrbjTcLDDRQYmXZZx3zm6RQw2B3cvrJX1OcoqN0qZ2SEYqjP2Ptu3iUTu7
EY5lImHdc5hghsE5sy22czsvex4ML9PlTYBU1yOvTn8LG3ZBfS86ESDoKcDBcxgkp4ADh2QoxiXD
L3XOHn/4lV0nJ6/28xzwBDHnALrt8deSoa69LS7H1Ii3Y3JmhloPjwngpnZT8bpkFcCTmJ1ynkEd
uEVw2zGGwqjNyiZ6IBrQRbiY9ZaxlsZ1eySzw78MH4t7auWoB+ybhXCxOHIKrwDI/0eLu09QPjkT
7D/wm0P3LqXckRDfiHkqZvngMkqVK16xoT9d4qgBuheGuFaplTnyXCJzMuV9FVgg40BlMVASv5U3
k1FAFVOLJ1EXcj5brqhFRSnNp5U7O4ZOrw1Ea4IUKMHNlwr/8jKjtYVLsKkiSNg9l5n/FSLTgubd
Tsx5pEN9rwHZJmRZoy461SFstHRt+q7JJUUSvO8rmTVC5IJ+HsZaAK9BrN3yLyvi0d2asSPAxdTa
9mgh7pZ2KbGB/Jtjj8KwZKtiUeomiv0kvfR61lOyLSwrHuhau0+FqejYhcdyQvWdwwbBK7BjytOQ
xawnWfCszfv7wcWx6wdzWwHZpH3t5CvYUjz5rrDBHxaWsFEx3/JEgvOaMbMkGAwoFnqKlW+o0wB5
c9bWVv974U4FqSECP/fP+ouNva7I7XJmKDeunRbQdgZmy3F/9Jv0fC5yrbuV5ilEUHM3pQwaYGZP
J0f7sURdCML/f8XdWbactQTYhZW5DZVudJ45aRYgzpPGC3Z8oA7Gu9A3KxzRqXtorOb9l3VtylKz
b8Fp6jF/uIwWpsmv+ey7iTOKFsygzJ7ZXuByo4CT9GE8puV0oJjDxqTcfxpK7vDZkeRkNJ/5pWC9
+0v6iMzFbu9rmkuIbCY/BQjqH1qfdYx61gseoERijZkFTHxSmgCqHW2sxivEd9mPkw1PaPm5WUlS
4eZUQLQqFa8nH0Q1te5M6P/0JRmDThE5rUcU/YI9r42ZUEnghglwffHVzp7J18B/j+ewFw02J1Ms
w4mFqsgVoLugymX5PO/6PpeUK2GQcvpMKh2XnhX72Do3hSwmFJeRi80S9FhUgkiTC4ocBSVFVNJJ
VG0qwOSw+APu52JzfpYMH0EmTkiKvj8wIa23OicRfmnzU1v3WYSJpBvhsEjRoMAT4HyHFIO1Oc+l
WY2ob8lorVFWfH/+sPOrK46+Rl4g+Mb0ItaccGmFMx1wZSen1GKR7Ynpxe/oZeBWWG7b5gci0Jdg
U6GLlVleAGWg83pQDJHndXyS0/kNiZm0CaDK4W0XBqk3ADvwtfihOYAAv1nhRXu+nMxJknbT2vEO
xqcUgz0Fiav1qiKYdwBC9g1M57cZt5FjP+4oyh79/cQVmXzW9ld3lur2boPfdgFZzE2gcIW21my6
VIZRODVxsy2CECseL+rWCAhSVVdIg2kFidjJ64ELM1yS2oTJNt83aPxrQHf5KQGXDoglxAH4OUI4
MEBBsBJLwvqwKKeI/vYXE20kPF755B18gTUfH6JRWgAz7KqoXKxqmqOotyh/OFGY606jyohlo62R
gTcoqdW3B6u0oZc0eWqWQFVFY7aTBNoLNybgU0z8zTYG+C8WTgBRf96+R34ffScUloWMYO7Q/De9
iva8LRsHoUWxEcXlyEJl6nZyHge2nEew4VcOiFfgZ7XV3nf4qEmDBo2cTN2B1GCXUsgwsBx54MQH
cfCQJRmxcnfKbmZd5LUfGXIlzx2zo7ThCbXPPN5zQN7KxQobCXk3Ksuuiqmfvk1w0E1KjgoHrKqR
lVfvt+EBLO1S+bGLf1zttmZdUoz7IDPNAsWCypE9y9CA7W9F9RIBMG5VppHBPD/iETPz7cRn73nZ
eVRsspw16l7cXAqb+p8Hi8TTKc2TBLxQBZuXXJiE9GD2O0U7BtzvAM5iRqpS8LF07Bf6dGc33g++
B6rmSRTEkENKJKKkLILHIoq/pREcp1kbf+iYJ/HLCGvKMEOdeVQ2F7kI+N2BqdCQ8KWdysT4ZXZk
e5G7rppy31ic9qBQ8vWmGX/rADuiJt1X4u5RSHmrFizmXXnkKjsR9sksZEolE+Gm5XzgpkcNlOJY
a4mBf8J6WHLJavA1p1HW7i63EneYgGJTCzfFO9tRd5GmLlmMONCKbtVL6d4Lc0ZWDJmiO/NrBsFC
Mi/pucKZlZrkEgL1Fk4Q/VsSgElp+H9mI06hlG9rDVv+NuHkkThEzfBFm7Rn9HOVgSCObVkKA2ki
1mmfhkY+na2GS8W4pKEmE1fXmv3m2KCAVPh0A/jhjjy1nqyejiC9/g1x3qzosmzqn//pNMmMfCNA
W+koWB0SOv6LKWgkKCwL7WHMGH1h4wdYAYS2rW0hRnFZjam7QTbs354m+/YpEmNRA7mZJqvT2lSX
kEQ5e2Tqei2Cy6A53UhHzonQbeHi8DyJXCk3aex+dAgogqwDE34RR5yy0ztj1Ld+qwxE1czb+C8W
IGa6DjDSO1wbnMUMtsfK1cEui8cokyPWWGd1AqMqX5mvHyCckd09pmwxV/fsL4esSG4PdgC+p3of
WmsbY2l8UxoJYpqVjahKCVHP7CaLdc2gPP6Jr7mdm80G4DqK1kntSGFs4VE5m1e8D7bRS0a5nx7+
cqdY0Qqpa8oTijA8mIjErumuXg08OQnrbkeTalrQbjFZmdPamEaweoFXUL1vVYjZS4yPbUCuC3Am
8ZVaBto4NzRyBwRCQtZh2cFQH+2RMB14cBHDTNXZMbcFIsvPBeLkHXW6tuyX9ypQPoz83m8kMx5q
rdvxCHLqmiuSDJLSWIONpAcbKniWIiWImXfX0cgP/NgISAwojAcL1GwHQ77Q0kTB8jYPvUqGNpzU
jsUA0Wuov2UYpKoYoQZ19fCrtJPJpY/DYN+opNDB8ACO67HGgv6xMJoEpaYUjgbi0FQWDyNOrCSv
xi0qqw/i+eAXInSYSKiM3E1Iw430fGwqBE5EbUHyeXvjqROSVwvzn4KOP/Uez4lIcw0WxqjHBFSH
P8WYjU1Nx9eon09MF9cn41LjaT8emUNfJcD1zd30/6ksrUldcmTJNtn39BSKJmHMNCB6BskBBAo4
j5mU4mfBvsd2xNH/SFbX89dgzDJrK+merb5WeV9T5Fll450UGaHfyFXF5z/zbR5+H/uz3oqfZCmx
lMhm2kNtQ8xxjKxWl4or/ue4c/9QY9Gu7vzZ5YZE0sV82jY1qTdj1mRWhCpKBFUwpe29UdaIcll8
9Ba5uS1zlueH8b9v6I9K9QnumYlYnxIRkfvKv58n7g0YZs9U0e+9+d609+ZCHgL8fHQ47wPBYnul
NDbGvwIZOGl7YHVnSOLtr5BdA72rPpltBaQSQV9RK9BbsYq6yA7InyihgeIkgD0Nn2xpxEc9DS5D
b2WEqfcjpOjczIB17TYDPiTqtKyfkLychpCJyXID4kL/aiakjxB67DlqzH44J6YX9HwmtAnCZ0U7
s2DaZ3dUGZPcyxIW48I28NQz5fZbYhTVx/8aE3poRn55y97/bFK7NePMMyCNamRjoCADLRiDVYz5
qz4uUvFy+W11W0zcZBxwLTZO4ITKgM2NDtX4w7qOrZx8MHwVLnTN5rI8vlhN7I2JplJGchcGMK1v
tqh17QCyGW2meNZ94i8boRRkmHC8j5t/517m3D792MaJJF70rYhS2HO/NV3xH2BdPfuqoB0gWC1u
LkD5yHKPsjPjw5XAwD9U38rWH9T2AzNh93qNpZEw3UveOZXiV95sH6YFObfidctrhZonKKze7dsG
4awAB4r1rb0/DHD6sI+a+L3ihV9dL+FbNBuLYc7sxxF+93in4EP7BxvKS+zR/Wc6Ma4EkyMCbP/J
JJVQnQWTiIjL7rbx7qE4bVnDL0ONdKLEid7HIbq5vXgw130RiacFjOCu5RoumPm7HMgaJThlpTdZ
HCf/5wLeP++GGB9LyX0HfXSDVfEbSVEvno0VXEqQouQZWK1A93PHdjQlnj4CyFu5mOAzZRpL2s37
JOc+0Eix8TzkAt6MpvKWRZ6tgvgf8gG+U/0CevhvpXpNOU4Npcot2lfiLjJ1lfOSrRoUy6gNWuJ3
TGh1rwmmRsS1hXkg5iO34/txxiqrbpiXRhpxyzNcCr3WUuFf6IDYbGFk6nFRk/lPecPVrcwSi4ly
kfxTcVwgpG+9K/5sti+fA3ZJ19/mCQzIH2fEe/poii+y+O1etM6+NDB8bjGjCRvjp6zfCYx5QSMU
2EAnJ74rbPZE2GaV9plAjvhs+8TBcRx3RIA0IjFizi6CvaYWSLDzyWVRU+8eo34PZ9Ot61bSPLG3
H5KIbk1i2S7iqnWwmrHcJAAqGUb8TPWfh9QO/qa4aVymj8tDwrj+jvIAWEv5mJWY7Lto9QJ3+A/h
esip0CipWF8EyiHePcVes48kQ9VZp5Bu0QsQX92fDROFZJkn1A2wPM3z9RxFqcAnw9Mq+yC2slCK
dcyg59eVZWwWZdyKCR+Ur1ZCwa20hsB6Ax/hgWY0ZxkE2IL09ldirMVRwNm3egf7wJ4dRh+BmggI
VcA3NoL0pqyM5ulrKtXdO57E/SazUG3+Y4DfqsZu9SFz+9FiT0FSID3tkC5cQ3smevUxfFvC9TaB
mYwuiwihwDrfZUJAJK6YHlibuodZOhLF1ZgobTr4ABn04r4OiHoT1ED0n7lRefUehXmvl9O3To8z
2ab174ykx4KM3wcVCw9936hv4CaU9h6viTfFl4pK0qDsalEZXW0ybxDZMTC685Tiv4lOvN2iKRXK
dEDlb23cMbMnmLdAFZTEJFjQ753optxLIhBP84EOeUoIggtlGNCoxwaK265K80QPow8VhAkbD5GV
dP942nJxhxjjevbp5jordtPEJsbIwscCke4wtGSqfTYk7RF8hChj/opmwE/DPHrOs9iuEG7I1L1Z
q1WNEcJBEVzT4ZeY5TAxDf4vyFC3l5SW+B5rHwJSkhOgWhWYRwnemOgo5vUywgYGvEun03IMZnOv
36bWiqRNeJrl8UQWxViCmWoffinMug3ZxzNQcE3kcAkvTVY46y48OwNEWGec47V+JkBOJHIBlpeK
pHrUJFBd/7d+aZ9kE856N8skMVtE0PxzNu3kC7NeK/IzEtDtoCWPMHIAdVSgy7osri+q/3cFqrm/
lSiREwBRQv/j3tjZQi9RL0uNhlbqXblvju+Ch6sYKI4YoKZO6e2zGCnfY5lB3K/yRdKzffWkaX4c
7quDlp+eCR53otIzFbA2QkMAAC36xWGL6NmwLENMVYiwSG4TIce+wRwkN67Ef3ta998vCDgSi1rc
IrIW2QFuHjMMYydO65h6bohi6MKkyNEsPaQqcqjhdz2GtyDm+xCxuc1y+hVqQAIxVPYCyh7pitb0
kLdlINUjB5lzgjWieYs0XKDLgZmLlapf04agrPqiD9TJJobfOS+aMtJVQph9C2KjqGypg8yTvzxq
+02ftFJmv7qPt3fUgSTsOxDjyw1vx3URgYMsENeWxfcmkNcQ6KUJDgz0HOHtLDBYZkC7m/650Qhr
yijViWqyICgJyIgTOnegfWdNIBhvEzg+IMH4n9JU5R1jQyOVyJXgP/08m6C4l+zj+5aS/NETAaKw
SM9wUaymfYwoDWGEIPDIn07RE3s6LPKZPWDisPrIRlPrBcDBEA5xmdjJFmIxkHtUMq7LB9SpiJKi
78kSiG0Gwi5VGW9KPY3tMIt9xRCkzMrr4MN/+g6mo4QQxxNk/JcCkLncKIZM+U0698tINE0aeNML
78v6kvQQB5cvryu4PUMhmmSWuzJzS+Uc4aj//vZ2iJLKDpWpTQh9oDGGM8Ieelr8J2/V6JxT/x7z
Ms+1Gv6X0Aua7zS+axRrdsP61Pp5eqI8khysSHLLbcZ7wimYt0bnaHfHOA+LWhj32oXfjieR7YUh
XgouMgYvRe+XPsUod9zKMgFXTYSFVKdrQ6Wjjvl19boYvk6xxrPfD/e440KiUF3YnFyZ1LUIK06K
2ed05YXxRBUud91yszY57wvyFtPP6ksUqf3aKRwgHQzQqbUseKxihBfVzME2Ai40e6cFEyyGjPpx
sIVO1JO/wYuy9TdAhzji6qYlYDdLebpXTIVqeVeU4vs68fZVVS06II6yyTWnrfGMtBVoYmUp9nU7
mUHH5qQNwGMko55mNnIemqc7Rm2BRsQuLXYtXp5SDtzeFsYaW+2wMxWyzikXTs7xyFWlhWKPkrbQ
n9+8MRFYyr4MiJPD+udVSLE1JS+wmN748r9ws9h96uv26w7jO0/w7vHU8bQMNxQTlUDzxnn49WYQ
YwMKiTpCDdEurTTSVyF4kHI+dgZNXW8D/8t9DI+r07DGLcAeVXHYtCJ589yjM4to8/1yViojODCa
oyDoKyrrd++fBR+qc7bWRnemMOLMkbM3EwsDIJEUStOJL9cSoZPY3R46efGJx/n3mbQt4SPtiZ2z
KyjeaSDye9sMivlbsmnOw1Gyb/ga1bHXgVaJHzZs2WgZtaMmpReyOwvutA5hmXzgo9xAKF50k2OX
swJXWAhEER8CF4TNfpQLfv44Jb1KVXkStK7hCQ7UNOIPotWYbQQIyfoKktnv8YrydjZ1S9Lir++m
4CqOk/8xZJpp3wIRKRWfC2pmdGJXAG7wao0GxK+muhJjucZxLo5UTcVILTpqwM2U+VrhtaA91Hnm
/5njCb9o076I6Gl7lpx4ou/QWnlToInqvE2fP20IkXPHh4XXo222QUaV2bx4QU+ERdhI9rZGqZok
XWja6eKWDAMuwE9Zpwkc2Ym0JNAUOm8e5mDFcxnAm7+HgF71kMqydduwFZofGvPSh33jKOBcx0A5
oz/mnCQOW0jzOd9l9UQ+K4KvAM3xfya+R84IYQR16ckENxGDAHIPgoCQZQQRxadwLRro20SxC62V
TykPxgnXmkjU3snYtRA6sHFPPgH7OqdDp4lFEcdIfXkEnfpiBBKUXxpZtM2Ir7T7XpK/SEtsxIF3
+9VPx7C6KnRxhF0sOMCM2e6Om7kWY+dguMdO/ZqD9733u291/wWk//KKVEaiN2No1uzG/7tOTJhN
LWR27zvCZxTYbo1WerORvZv3we4/s8FiLvCLYyXUDmZGmTTGimd4YVD1GwEiZQwlCIZDh+HALnbO
z3weAROoo+xKc52qRBYheD6uHhVyRRPppqPAb/LflkjJH5E4a7q9ukUeF3h2j5H9Tz+5lNrDmpqR
XCgg0rVEZJLxgphoj13N1/CCZEwIsbUWIj1aof4CFAgTfdktr8zybyqeaIfFnnNlKRzvzKtuXjIN
sZkAK1gzOs+aIFIMKiA/WW/I91u4kXBIM6HMu3dvjnwFJupdEDxhSCM23thTOWawM+l2sJ3LNO9r
7hhn0by91/EEyT368tbUeS7foQ7ZBWCGSQUjLcTYz2mqMCeuHMnFNXKy3Swzl1rzyHS9hr6QY8WQ
9iK9bphpTr0Riv33Bpdvl2EvbsEGwwnDeS1GH+i84eYsCyKs3F2hT+Y2txr9rzm5QKMMkyg2MiI1
81kX+WvZmoJ21t+Tv85Wj35xihdAeD5u9CE1cHwEPUTlXkl7hAPrlueleK/MlMo22qEPfVZI8bkL
LdpWALMdvHQB2AFuRF/TbPSY55gK3a5ia8W0CVazuAPzsVW9E5E7LpG90R6Fk7Yse2AwS5/NuqQ/
Yf+RHt9lwka0cVC6uLhwwwNaezJ/ex1WSnKK25VAK1J6gTQOmSwzEERE2Z8yBq1UZca7ahPdk98b
sOiuB9Hxuq+UefmaAYHNTP/qiP1nToCF+SjoHTV4JO8Eocztt8lnhKE9mLhGnb5eikgc+y0uH4sO
YaSmjs8oG8+90JeokTd2LHScVaJQQyZUdbf6BgX920tSKeLdps3zL+woIOwC2aucRhvVbNFV/dpN
4MZAs0yQJq+6pwT5qXlJjt+dOMUMY6e32PLKC0QimTAfdSd+LV7I4gt/C2ySKGskCP2BImhYBl6g
Om5MyXxuYTD2yDD9evm8nuDZcy3q+Lz9VhRsGG2QmNTtFON08/tiI4TftFXVK5dXLx5BRiUVMmfv
Qlj18/WJ6gHme253B6x+CVMpXR5J1L0IKHNyl/b3VMiQkYDWXHFURUeHj7iadWiqMnpvLJUcCfQx
YE0xT6f4fHMCeSQQBa4bBZIz1AKZ0IEk931k4mSVuCqpwfNrsZEiBAqW+94j356fSbZc11ffnozs
6oF5/fLyIRvYgQ4a5SuFQ3CgFS3KCtCYTfnhMiXvgBCE10tfzZC6JtAXdlqb1/5+ykEdhTyEQ7b5
k+AyAtz3zp0nEdKrPEhhLcNFrpwkhR7w5sqhV4SrBbUv2nPJODoaFwRCqRKj9JtPxFZZdcRRNJt/
tSOV0nZ5fS/szBZ1EqmGnmuH2Zfth8o4CkTR5oVIXdfgXPtOKnSoJowN1tHEKR+kIWo36yWhuWXM
e54LMD6FaPLtHu2ryla1JUDJpvQwoRr51A8cQeeXnO70mEu298btIyB20ck5EU9SCIV54ciKXNy8
C4I7eYqsLV8RfNwFqo2nI2c2A/cGwc5aKUhThENfqdl+y+zDcagTTeTyIbZpncivqLHfXplIfqkU
uaefB1aW2WfvAdlZxaPedlgWMY3NO0KUHxqqfW2vQMyW/ydRraKTCVlaIh1p212ralLFnGdIgZl9
TRhTAUoHXyaup55bFR2UX2Gh1K4YJPQCEZQhWBgcd1swWhiSJ6QVV8cmjqXFEnfK+s8DTYTVJ8cc
HRF8njUzokmFhAzy2Xqrus135Kg+9b7te/CxZdhXUx/P2Qj3NW2WRtNzMP2Pc/godBpOqJ9zbWJh
6I8JvByJqFLqVIKwMBOq/TwVGslIPJgnVBLy12pxZSK4KjSHywiUgq2K0UuWKW7UD+8eqKWwnwIt
C9qgQeVXc5NTEq+3VZiUTJbL1Rv1Klzlowv1UF2UIXKgci5EWDUZWDejjacL1Dd1Jkggc7x+N94Z
ZDb69oYpU1aIg/MlhwPUonEuTWQa0Lh/qFNr2X/QHk0Lo7YMuQyO5YcawabauG4AcjlZDkMtnF+V
XI0VhNSj+kmJir3942kLMAlmdB+lyFKYxDBeqzFGJHYP6nnQgsHAb3xDbsVFoyq1nDOm7y/u7wVx
1XeJPipHbcnbr2FtQtBhbLa3SRH6/xoV0GTCvGwvOXvYOP0lR0mhjbjx4TtkQRPHMTmCSuWffIQu
7kk1jFvYfuyedoQm8tqiZlAcwZ8kLOq8lEZaqfDfZ4O4u3gc086IKz36YcUFs573oVkAPhXn2niu
qDRoP/OUZdVILAn6Cqzkb3teL2k1iyHMg3wCwAdER9UTEBKNej0NojuXTtOnaR8+1wM5UgYkYuYX
eVHWPAZLsGBEB8mFOkOsJuEPfqdSIvps6Ka6T8a8MBwWoCKsKQQ5ewpRhVbcU1xpttKqxCrQjqNj
ik6gEqBVHQspFtUlCDRSqU4PkSOMJrnejV/4pqM6kBgCrXOp6/i3Ebq/yC9sED9w+04tAl8z68Il
CP3a3c+f3AY6An1RALJ9XiI7Cja6qyirsnDboc+8jVMYRxWCWYGBIsMa2tZDD9aODRK47tGVzluX
GYdBLDKVCrqD8XtXKN+ZfX/j12FO+LK/3v56cV+8nBRtc4xBLAmZZij9H5dvdaB8yRxdwHKJfL92
lmWDYgst8a1i3+tDOBe5cQjXCsVe2Gr0fuEPQWYietQro3itD+TBK/zVGLFhdLSL65SKgG4fgJn3
fWlM/EuPucNMm0/cCROnGJka/NENO+EehOG0gjv12XlTVaKZJ80UwMxDDBVK+OWjPTqHFWC+0nbt
5D2b+/EBjn4vrKPdse6NkgTocS+Ow6G0nlZlzgbUOk9YsA+7CLOx/HaXfmKNdullavX1UembLl+K
uu1bq67hy3Mxp3XocruEE9nKxZLBfgNbyDmfmLvwikAYchOHk5CsZiWRMg2BSvNnACRMC1qXLfFn
0weOv7EG5+0KWNn856/MpP3GMyE10l3AoJJDLvOcGVxM0VfJP1R0f7B+hVremSEQX39Xcal9TRFG
AsSF1iD7tgZvqSYO0eLCRzp58449Tc7jdUVt3XAka7mS/QR8HXVfZWHOpq8WZZFkHuMK77gDJ8VT
5Gi1pn6NjeFT4tSYtzi8EwXtVRwwzC7EQNqCZ7U3J7grMZF1z/tMJnJiryDMVObMNOngXreBARJH
TZtt+LAtF/PnZch9a5d9RnkQssGvDl+n6BLK/oTN3ooETryDNQrieJJHT+NxNWdARlFpUX/N00pE
apVrewYMalc10oPHoW313w0cquVX0+h8/uXp1IfOYi+84KYhZluO5UFC3UYWAfKF3KBegNaZ824w
Bn0HZEAbEE6csNfmeTIo4Q8Db9wMsNY9J968gLJB7IsxaVPleRDIZ0kTFhJGk97pcdtG0oyLXP/j
xl5Y/TyaJV/Lz8O5wvlwYQUNOvto6OLHsxQnQ0T2uxLBWHP+x7PFhrKz2S3gP5jAHFL5x3VvioFg
kXAemFOyVNuZVCRQtWHPOwuSBTe89md4EC0stoGghuWR2gEdZ4xbMNnFLeoddF7/2YwoEScdOiDo
HYng8eA/OPfOwLfwxzSpyvLSYMOgGPccuJrbi3swwO3Zwcyx+BqHmG+uhvccRddzCOUD8vMPbzHx
0M3o8Qq5IfSGX/GasGPJh2eC/6CHKT4bTbf6KhJ6Q6Cgp+orS5aj5p3tzYEqiWsNvSkwlVEuzGRp
iMabjWVnF1e4PwyUn5tkFYGom3m8sSfsx/M93fwenIiw/7kuPEGeJ9XTtw9ddsh0oWdsOuo1g50o
Rx7qEI54bx1urEH+GLk0m1nA8KmzEhnd6Exp8AJcTbdJRp3jSVMONbhRCGFxNEybUc3T/ixkozs9
Y2beqlm+gs7RFR68gAkTMWW90fzb4yCH1xaV5OHoeLk7ofG4ENTvy+Q61lzfUb11fM1b5uFnBSgP
uDmQ9zWbRTxAsSFT/yhFn/pPWD9D2l9EY7Nm8mpFMwuuSCklpyR0cuMmCJWS6IizVqL6554v7xFG
BJDFlJOArAI/aHCA/TGiC0cXO0yVtFwg5ionoMNv+ajklCuyvxFOAI2dRI078Vjz63K1ejsjNbYe
dqeze/+iLwwLRloLeETD5cAxtUFaRWaNWnz/BF7sFzGUD7BYbKzL1BPGBj1TOIFJPWqYkqXDACOJ
WVqZvkqZUK0U6siQX0/Ogn74oxFhgoiaOCK3outz44ToUvZ8Y53pAhHYrrU24EaE33QDCoIA02nz
R9uuteugwkC2FOwsB5XUpXevn1CS2493Mx+/GtY1XSU3d24K4Qab4d2jFS3uMX3V739A+5IuycsQ
3WyYzQVHrfq1twyVQsTUU2uJIlGyK5ydiL8NzQaTPykT0wl/7ahgO6yyzU6+Ss1jh04vHxv6waL1
UTCZq+46AjVSK4kao4dn1cPaA5sDBXIDoPl8fVDKAYTxmlN0n6Y6Y8ex/ORJatjtzGooyGLdQHAI
mLUdU89oW+UA7MgiEw4KR00RtNHJX4fpga9ct+jCejlig5IxV3Alk7MGUMtsY9oakAdWVI8FjVQj
3TCg0LTmOjr0sxja44tKKG3PKQDobwEZd+o+bTmaFXoV8kytmjwv1xXWWD9cLylehJ6tyU7cqFHw
rCicpZy7cK1St4nd9pJzOc7BpFvsaBqS1VAn1IVon2aobdKKKK9h9vbJic4RLg9hs2Jq15iHyW+C
1nH3uuWtf6RY3hOxfVXu2jCOxe7CkZcavx0Kpk/UduJ2g4ki+V0KPXLVyKDBxaeyJfhgbiKVT9QY
Hwk6cqtWil1gaTHA+POYeDFwtx7IwnF0bMPVLcqs8dx+yXLayXQcnkCXAvyy2X7Tf97NDl8Zw/Rd
ZM5xmJmc5/53Q4hgoWam3qa0r8Zprt50v7IoRHtKHRopIxw7Qv4EbWGeJWM2U12K/b+f7A42t08g
Cb/6HYppSLHHtlT/jJ3azzN3PbsLvNR2hhrkGmDR7qHUz8srDNs/etfejXTTLN332zRaNzp7+ctI
Wpk1Va6dWulPQ/XiFAf7gpVZPBl1RCs71f/2hifbaGUtl2kyEZAXYdPP277E1FfJqSHWDzmdv/EB
A/nkofAAXSgrlgAgLvnasmQp89HYKxAzOELfAhjuI1ZaCDEaRUcfdx6tihVDNSOKFuGMY8fEE5i2
KCWouzdPCODAh9OniUL1f4ULckYwuraXpZJ7dqId16mTMs3a4bcNUfx6ZkucPYx3hp3q12peFpZv
dQleUn7DKwjhnls7eH7HY2lm6OAfWKXcsxTh0uYQ906KKjt2gInZ2VFwLfysKgPi/EH2WKivPtGN
LTWH5oYqusyMFpwHqMe1dyuwcbY5FddZDISoBThzzHeLwzHY+LCflJD9MAVHFIfkTmArEzNYLuEa
B6vcw9vgP0J5ZLYqVrNx53M8S4VlYEKBGYJRcYNP2TkyAS+JZwpbXat5homJAmcQjc7eFachkxm4
0RzYqxsndJKUNXnk8twA1ELpqawaJVnO54YGCq165mE9t/1BPDIRiDN2bbmTzetwO6eGYWqcO3oV
ixTaGMwYJISW3P+kstChclN01t+uZmWH/otGtvGRdkajqZnQHxgUrZkvDcrXL+HgZXoUMpCcIQQC
Gmm7wXRXcT01jq36CJKz01OnsGJyNNVzpGvbw86YnepRwM42aRTYvkgUZbQpI3eAlTtFUORD1Uri
FSPnVhL2qPkCxeXj2OlUGIwPrhrCwDwYmXyL9uJZqiaO8vbnsvHQjXIfBogRE54dXmp67NFKvJka
RzlaCIfUrWUwb8uEql8Ra+AjF15oVyaIBLan7XWw77yfV/jcvS5zucucY6I5pRzcnOpuZlACvtDj
XwTdx+VIN23x/c8aI/aPPkl8jO9qjhLGn561kwQpuQ9zRLP2KfXJTGJ70lRjexpj+04qsDURFdx5
DVimCC+xACaNeVpKSZ2fOM6pk23zZDSQyWBH1yJDMooehwnAGcuhRl4Xy3KPtsABbkbgeZSnTsYf
nfwaBJzTaLH4eidteB+eXdNnr3SkQd40D2OFtahhA8cdWXb1BzQVf18GM3khRvh7HBWuJtdmeUB3
Y6kumKOxG5RrVz1fAEhu27pIveemMVMCeZc2UkurXvRRkjCj5Wjc8PMDAdYIvASuSP7Uwx+FURdx
G5yeO2+uDQMOroTZ96WZn9luZftoLiy9WNWtRmeQA2bx+tnDInQddd+1lxfw7UGpzro5d/HBwOcA
akj2ivj4ESztRos5zrMF1xyqkclt8QseCqxc+i9UKQAYclTnN/wIo3/UxZdPRpDlnWaOHW2jnnew
d3x7hZas3PwZbeR6RFJzEMJrgZsf+S9WDiYs3NhufSAB1SAwdtSm+YKSjGmnop/cstFvWGaEcOOE
bhMcvkJuTig/d6c7YelL83XMLCahmX8+kaidBQHKxZsJx0hYvl8zn2fn5OsW+cUJA65cCRjq8OQP
5TPTIN4mOk4vIH1CPKKkK3aAh6344q8wPOqniJKsqqudt9AzmFEQa/Ht0z+madcmzUVZNsaQAUES
pJmX+SOQ4jJaJG92isNHj0mJcqyhRGiQAkbFA0MCNapvT+xnBk5BBaU93dH9xOXQwbOdrXSCE6dk
8FUZ71sWD2NC++ejsCX85VYJzPx/MuScG5puGDG+pw4FSymx2Zmlz51aubfzA0yxYt1A84DO59ky
n8p961XnKAVQhqMLBhhom/czYNRNk1ZyHnZBp5Fj4p11DUMhAPj349nzq1yaI2qhHnz2t0/mVHQd
9SSvCWdZ6MNGzZ3tWpKuPF2hAl8UulHYOXM7+XwNd30Igoe1MOYcpDpjY4zH490nLMwAp3IpUJG4
3UqCv+I9tXX9O9gJWKe+PDyJmY26sAD5hDFgzxnFRZRjALqNXIqlSCkXhIpRlPosotBci0Op/i/t
fg0d4naxJJVcw7WY91r+u05yDVVpg+fAvwArOPo5gcW8APfRscVSlceKv/M/F903MgSqUz8kRhV8
XtBnt42b08EEoZSFBhH6a0B5tgY3AcF0dZw3fxxK7cuq9AIDAqgpeRs43aLbiLzRBCMuAYtmbt6h
uVpL6crmYdhdginMvL+6NNHcm2V3D2LjG6ftZkq1kY0HW5c1Lq9M8+OYaR9rMT62V7VajQkDkEnp
pclmBPuiJhTLX+cZVkqW+tEkuwOBdzoLy7PWPqqEaFb9cvpL6CfvmsS6aXiE+LhvOrnPPCkxTOX2
3CxtA8x5dib5vj4cyDxHHYUwckgSkZKT+xKsZ7+QN0nIWF+xB4P5QIAIMDc7dzymwJ/YbciJk54I
vvnmagbMotF65uaHgZYGGNM2Q2bKWLmB3pLVLtyHOmz4ICEIXQbza5mqJc93LkegElbb2/xXpsyT
yO8HLjp0vSN1LWb36DPuhV7B2gPQTgLG6kKjvALjHCo+5EE7BG1/TKevnKC3ggpqjzB1CSM/8ZB2
vYROfRQ6qHcr83OZpCgB8QmfAebM8YelC2dAEuFjJOceySkZkBZRH35VtmYm4PVkXrlAIeO0WGJN
iROp6f6S06TF+nErQKq9yOp9ijftIHM9eggvIwbY0/2xtxQO/iO9VODsLceH2zMqf5CbwpBNfJeX
x0h0mi6nxAotRUeDJ/jpEeTgRTd2yT3RBAOQGASIw52EXekGWeu7L0lcbOGAg1PswADmosLoQ/4G
YM5a760lGiaXQ+rhSTGaqa1+zwf31X0DOS9mUoQm/zUs6dYJZ8Vbce1Nf4J3P30Pdz99AcpXLPfH
zeVs0ZQHtkVgRLqwIsVzPgGqQgKJeLIv2tBXvlG3BaaJ6LIuD/yJHipaM0TxjMPbjupQaKHR8EIb
b4WU5WcbLlpr8s7Rq5cb2o/HyodhOkow/CPonRPUhaqgOt77SOJ6l0OwArfGD5h6OWm7noec5b1C
C6vjTA7RN8cRye7CZ/lu/FVnYM8BMIghpUJKtj3hjlvhdN0Hse33/Aw747UgwgKoWthJ47XNDhu2
j403lNyfVJ/czGjjMm3YEaraXGosBaVcxaaNkPxY6q8DEuH/n2K241GLEok4q8L15/GCaZnJUDxm
xihr2UX8j4iaHRHHzb8u9VxN3q2S4KNFJSseYonHXWG4iij0q2IxXnnOSbJIkPA5OFvXmx3eJtwE
enXx/Wn1VHDZz+qEpbRY8mWuhtVLLp13S7irLhzpCKwkAgytUNx/6Bk5ziOmGp2S1n7imMLZ8/QV
7L+srqVbB6Pz/2rEUiNiE5kBDGvg3KexELcZ63DI22YM72H15Xd39ZU8PdI9oGeOty9g5UT9up1m
JspFxPFGUiyp/t9gpVbyB0dlcrrePhTIopMJpMmxpAvddBecorgn1VXff0SKNk0ARLhq6xwUWaTi
xvuy7kvxPkMWxBtoszw28/uF8Ous0RZ55iHDOBh/Pm16yk+lddISq9FvDNCTbEsrhYTDBjvl/cNQ
ItZoMgGgZvpwuy679bcOWI3lJJ/Ifq2Rlk8/7nvDcTKOB3MVq0MXbe8Jy/aAzRT4FkmmUARBLine
GAjkc1gKopJICfkJbQcOUQ4omiQqsF/4s5EIMwcpqTbY4aUqrAJyZrh2G1j3HdnDbItCafOIBASX
rezMMaGnGklIqVG4+dx7YQwwXYh6ZWzfA8xTlDoaDfMHnBhdcluX4QGCx+877ZcrOZwLmwIRpsOX
6PNjRSOWCOnhqtNR4u47RBanRNLC38K6JqYW97+fAJs1E+uxDWWEaWQiWWPhEExa/WQ7kJIGrIxG
mjlWlTAQuQVyT9myO8zONh6IDC85lTTUDt3OsoakjrycTbzt/HOe1+QMqSfT/e2Inwp7B8CnZkJ8
6i+zgw972MNWPMMi7FlMx1fevcRwYajl1cabiEaNxjc+ukZFOcoJ7CwrwdvV+qBKCkQMfMbASf6/
a6IxQAAsn9ZCzfN/oBxrrvdJFP9sMhkUJgHQ487QWNEmmUkWQNYKmHkxApYN0h/8QfYJydreSHwd
iU6MIgG038pCsB0CO/exzUH7/iNsXNq07j6n2oSYgT0BryLolkGDfVaHY0v3U8Jh9DS8MwRcspN3
DKBoordJUh6XDoLmLQ7mjNC+EFWM4TSM57rmBkdsH+AQIejFFIV3PEE+EyD85OlGzMpcvGV/TV2g
21rmBsrG8xFZdI8b8hV9p1WbX9C8twQB9Fgs1JeG+6FXT7t0nSgHMVFr7H0gUQxSBOQCj922dHh8
bjb3h4aBW4eSeOuA6oQrGPUU0fn+RzWmTE8ilWl6gSJVmCpxKR5Ms2rEjWXFoRSl/SWCyUMcx/58
85q84UWYIh77WqbFXBBVj+7HsIlcw8I1NlovTFb0Sro2S1XwiFkVfzLIKKWS3sKK46xHPOYFO2yf
uhJHUtHhY9TNRjWsMixZTKJfdAlJ3QqpC9q9jC7ZUR7ZBSs5T18L/y+FqCTgUSUzLzXHCTydCF/y
TbbY8/WEjutwmw18msz+bSgQqwYS6RqexF7mUWaQtBAumxcGZfe65GxUWLMnWY5qfzRzjR6LL6kl
q9MUfui2lqRQX1zIVoe0P+E/ryGZ6kNxS2BzAeol4c31j8zn7p4nrmCCnF1jm0Z3OhldBB+udzPT
f/gwtZ4e/HRbGHWoT4Mqshduvcmh8dPOfU2u1W5fnbvm1axfY3YIvW0dlvywODv9hrtHllgDPy9I
tHf/SIl78Sql3Pzl4xczfJ109IeA+OYhYfpnZ3ig5OrBksGSqLFQ5Qpx96ZW5G0EFHUHaFlyzOvB
x6Q8lmLJKCFrTiYMiKG03/iGbu+Evok/lcSjTS460POyxhokG9nBt6qI0J7ZhXjAnszzz3LBNI9T
Rn9woaIpb45ESxV8ywGnzk2LlmuXXdAIN+Sei4+/Pf/f39nDTBzKFliYktrbyho2WrhMe21vb4lC
MJT47UwKw6+soPcIv41N/7/oQSwQHmd8NaeQ7aoTMsCGulrfOd59JMNDyU2FGzmmYSZfapo13IPy
p3UpPi4d70Bbt4CeoQCd3moVGjbMUYnQ/AjwGrAp0cRTSzXFXKaKLM5oYYAo5ez7JOcYIOWjvvI+
gTx8QeJr6JX0wUD1zEp80X0TDE/yVD71/DKoDy3QGDa0uForMo3OGVnrY8LNVz83STKSzi6GVt3o
yzyPghREp4VZrYlRPCDZzybDKm4qK/eJ7u/TIrz6oXBc8w5xMB18lB53C5h1hD/PFtF63GaBw4t4
qtUeF0nfM0n1B7LfOFxqWvHsfm8GzZ0qp2JI0cA3VQY8uep/QeXmjrTsxIn/p4nyGkWDceZHu6pC
ho6YQVoZdub/qkx2QKsVpJO/qdn+vTPUqQNiOUmF1ghTzcma+Bxrbq+Wx82VkSADgKS4DrDYohVm
s7TF4JFMTx9XvOxVp1s8Svvhc7DYcSBOvJa13tCAX+S04vnuPwKX1XImlIsgxc13dqrfqBOxkpj7
Aj625PHJVcAPR7N8Fs3eYVPsBcjOoAUo1V4QMmPjpXrj37IoVW0K4pHgQJX8EH1InadaWUsCuAp/
e9XL4M6FvR6W9JHjGPOtNsUitx+AKPQRtwYUnZi0r2Y7PRgnWqbBmqTnbBeNBE716TvDLjEz8taO
Lm6XAsRWr0cXDBMuU5yble03yFM+Hxy4DnealMxXtwGp6r6jaq2d6vdys1pyOXWlRHit8N4m3jl8
taWai2O0gpiw3H34KnCOT27aUuNDgAHzZZ4oVhWqPjUo+6wpnVn2mqtisyXfFGjU9o5/74Cv3BDY
J4N1/4nX5pfjYV4hSl71f2unnZQoZUFKWNO7H7E56KxXAXQEA0GLRmYnC2wZeRuLSpjDpnNnGTks
ONCYrcqYFhuvjUuinSnZtq2c58jlEx+tsjE9qg3EoQPFoZ/RjlUf1cFrd0u2a3clH2YjxshG2rIM
NpzMHk+aszAu7IoKEaT8Fw1qSEIEeeDtDdonyaztSvWwWbev+/3lhaG+/cwbyI7N/UwCrbGeUU/j
/8lH0pZ4BDyGq4MncGcvt1enKQqW4eVzh8s2KFwCrZiH4TYXdJhHGshuYk7E2+l+H3r1oj2zUG5G
w+SEbZ3kDlQ+E7VsamnNtOylWEIigM3sOgzwKSjPvzftM9F/oy+gR951bKlAdy0ikItYn0FLJGd1
SzhMJmrWcx/+RUXrMYJ8Nmu78FLxFYyLadLB27ZCiJ5NvGGBSe5HNJV1XqSVxJfE3emCebs9pW6A
SGjadgOd3uXoC0/DBNReDt+IeqQb5kLscmuIi5Abc4XFQVuuIX1zcW1NDxVNbZHaxMgKMGdEnPYR
qPMTHrA7obgxQBnS3qD7EOwy8op5HRHMpE1pR/ZJqp5EShK3ogfDG5gOkCwr3W34eOBE3/G4xLDF
MrfJXRv2PSfSo4DnsMvofzZchRVGCgwPGFkeBah4CJbIgvu0CCtCH9vz7W6vxjROhyt5vASW4ZXh
QqohdbE4wUN5mkRFfi1wlpTc8Eb3iS6ClzDUBIFvoe8h8YnVvtWj/qSwQ075MXAWfKrTfoPkG4Tt
4naf8UGaa50+PsHSEenU6tCh8wHxeraXvfbGPQrZDOxCeIZtzsr8lHgLOwcAM04c4WUrqTX3xdtx
nl1H+ZPc0E1uYquXifzyilHHp89Pk9IvKyrpSryY7MmfOSGHLwiqiuj4DRN3Uac2cphwteGva+1g
U7SKpnNDlDJqWeqkYO4v/+nah3IM66mldfBPapQ5O4cfMQxgOP2GJ54TEsWgb+CXivur/rk11frL
FnLHwfT5lOw+Eokz+L8QMdCK7/jHQvhFwOJojjtO1qAz/vsCsnjdMtj1obGMtgs1FRXAsq/A3Shm
lTX9ec/DDLUf14PdPtru6ek+4CAv2CxQ7dOblc68Etrh2P4PNGu7fU3GAAfUA6BcmMjBgV5BP8US
zXcYjgLLo8pMgZOcV/+D6iMrgXHfmLKplDWrD0dqLYGoF9DHLm1tJRNnXCEb5zugCHTcVjBmE7iV
Orr4k58YS1pJRtrV9mZ1HJrI/NubvHm6m2FRkgvkOgD6XD6uJnWs7kihifiZ/OoE1kawqWsqj/vc
1j4xlYHM9aku8YbWLp1+th+TnJRGAnj8KZ/BPwyixxy5/ZPLxNVq00MV5DRJ9ZZNziucW7QdeHl1
ZOb/7mlz1L5BuaKWLZmaD9lskvVzJiYf9yEVSUYR4saiRB996z9qceFSoAoBCzXiQqDKzI//uTMl
lEd1ADCo+XKYlxLnYdtkwSD+L3j4gBohMmcfcNXUYk4Aw6+KqOHtsjROOJKacWUrXmtCT85EyS6P
CZ7Twli2CazmT0KpVQKw/V+2PUT1HYA85XLe1JxcHiesSeupktF8qwTuZ/IKaYkOQg7MUWeE+3aq
vLdBX9k8A8uBauGgVX8UQ5E1fwfzrL5fTNCmHR4Fa6DZuZ9TFHSOaQ4FX8Q+/RTSm4xWQd/uf/Fh
V9V0hRVBzUQeZ7QIUQnp5jsIBgzl9LsgwHQ6JTxOSamn/A6nr+vpypGWRcM0XjscFvpdv3m06cEV
TBhNOqT4G/pgpZrUplibao/WbICj1B44D5upTNe8lXUKfnt/5ciQtY7/WSTohm/pnoOB0knC4Lkj
pcvGEqqB+yyt6pH/dscaYj1+T89PUgr9PkFxE9GDsb0elnBXcBQo4daOeHAC50E/aW43nyRpzsqF
+VA9RzZlyftAY0zNE41Mv9SQpeCh+w2E8gtdTOAhyXqG7AmHftKjRqnNm44CQRQoR1Seb30WtFMn
ri0EvoBPZKuzwP5Zg5K9L7tLOgNvD+NdqouIqmBpciiOXYuDV/TN5rqQqq+DqAvQUZS6N3q9y/5A
6crkOn8qZxlVqi17uMPC/xsTNyjOEOwfLPZasiqMX5N0S/O0ldlt7P1es8orPuA1XfRSsvBkoD6M
+l1kdZykHEttMyD/eQkCiyviIzQAi6PufT66vlO+xdYkseBBpnaW1psCAlRc0/fwtPQk08l40xAy
OZPToBqNH2rmTg0byEs1YmOe66gcldByvXG7KFszialE/UPLgJHMJddX55wZ6eu+hisr4u1GIFA8
bjmJ9wgJOKfqh8VJVM5pAcWnvpRvZ9BJsRCngL1xc/AW5L1Qf1oXz9VIfiPQcxLaWJFid9DwlhX2
tcfs3NueAyaMggPBZqn13WbOcvipbksRUQhIeNcOb5/6X354bHCurvGZ1hJtasp+9w5IY8agUQax
Szmbx+ftnmE8uJDB1allrWoIWo1K9NwlcF+BgPIT9ozJIuKIE2mXrVb3k/5S3escDLjUEgnFKNZY
d17RHaY6+Av/spnD4ZG9gR6jSnF6Q/NmROl/rwwWUIo5gSZG/FhqV7fqm6ft4mEEtI0UoP4/N9th
ZLw3HI7W8uf7gm28gcwuIV9Sxcn0pK3p4GePikQKRBrCjjpV9FZTMEBIx26HFbdNdzBxlWytkgnx
hWF/WUxcu3jRWg4eL6IAxAATM57MuFCbD0c9gjwNuZiL9PSkQ5wOsFgifOC/lYFQYS/nIVEXZrJJ
hO7kGM7ipYzNoLB9HABihy+h55J/gyyISvy2lqQ6tdhMLSV9966odBncvJrriV8w2YTy3W3wWbuR
okcZRa4rTErslOO2qAm+9cVASCGfniNb4jhZDXdlo5P5hC9CesaWpo/bCHhZ7BoPmL9KOjQ7Svel
u7mCnwhRwh5HHteUrXpKMTqqUK2PqM/bd1fpFD2CStPQzlRxpB6sm8z5mY0T8y6Seshtd1NEuOWi
3jefpDiuO1QuSnKV+MhOr5xy6hCSv7Jr/ZRSpd9VNQq6tzQcsTvj8o20D69hQFFcT0qBuBDxHrYz
li+KQ5ahRDfWEvtQwKLAhykc93G7HQodZNPhFrJLhSLvfBUnYmEJ/XUSadcYgO47SoVF18Eo25uz
Ea9ZP9wfp+qpBe/Qoj2qU8q8RcewQwYTPvosA0COTOapxq+sBQCetZzSHEuVVmvHQKBHKqUafrwc
CzNgdqIBeRbGzwQVsSlftAPoWbi2R5DgNRg6fRaySb+JeI3H+WPTZLJqmwZ3+nb7wi3EsseCOj1/
srzv+QJyFV4pyS4MxYosix0gnztgEWVG0LPKrGNGImKZmc4LKXryXe1kvGh/OLu/cERRLJlBnyFt
HvVTgGXoGToaDSIKeG1jq9sXaBOlqxBZIikwizoXMqH5BWhMDR8aimmyc68CcxjX3oxoxSuQRArs
PGDXYySWV31hR5bmN6zW0HMJcvGEAmy5hALpVY10TK/Ok8kNBZw+gi24tKguNFxDOMWRFcbR88Ld
Ht8fsuXqhWS/OHvNA6hzlxX4n975mSjz1ueqX24NVXtho1343ETiffdBiuUCg+e8IcH3PVwtlzTW
E13sCC51MDyyOEVifWDiQgqC0JaB6cAurwMdATY1CzuyHarO+n5OH0Jaa4oUtT0nnjU4PB2oezHF
VGQ1TYbc34T40B7wWL+duN5ksGXLY3azmwTmvogXn3feVYouS7AC4hn5dRT1kSGh5TxzH6xDNpZV
2QuYgPVy48P/XAdVsnzlpKfUAnqWH+sh7e9Yzwl2uDoNj4g093qQ+35Fs6ISNKWeMA2wdoxFiy9G
ACVmuEgHX81gAFmFRZChwu0q7yx4EFijwzs23aPokXSecjGdoXtUoNJ7EtQwGjWhX4phgW5IRnCH
lCQJ9YkdJ6mEoDNzXWZp8o0D4XhOe9lxDVNNEfaZH2l3/sYcIkd6l6R/vMJOUXOJR0hbj6P2Q2TU
DzuJaLjQqN8snF7TSP9GkJkG4JpXiWyUEuynhJLog8/Zy1+7pQ0hqMof5/1MmdJTPX2ggKJmRM0G
QyDA1cKWhDujMVtxIyE2M3RSW53cdjj2DzriOTOdEdRq654/pD07gNGcbz6HngIopWGUiLz8wG+i
7nXyAUIzK8OIkj7hKkPDTVjCeTNyhKO28/oC3M+AgRm3o6YYn4FkxhR5bs3Ob/MAN6SJSC1owjse
1Qj1qAs65BIYuO7w4fth4dOKG0yzIbJUbbytyD6Nw4IZrdxu2vBvKAr07My9FXyDrpNH6huhGjdX
EG+k2+ExkvDls5fjeUTmUdOyFoLwzKLT7nmdLKGJB0mBnA9yOrjU/BNsQFPm5bTRzLaKN7sljXuD
ZTporkRhJW+iq0n+3syiwJBHt2SYB8FeUGXn/xW8CzRhVBGAguxNL9mSPiP3ckgt1PkZ5krN6IPq
Zf0NRy8URRwrNqTMF4jP6bK1O1sVlA8hMqB/EGLdGp5l2FtpRYoPPR+NbwXeIxcyIXsP7IhBHlxR
vWBcBQkGYqLXr8iFying9PS1skqqrzTztDp6Z0vTCW5o5ngc7hFt6adC8aVJoxQKTI5ZELP7uXZK
iNjjvnmb5io4uTR5sxZhRMLvQWmRcaKuGbOgURbEnB96vDXoifqvj0FkxceIoqaCcQKXYuek6dcu
GR0T63FgjvLyusH8zBBm5hkjH26o3WSMPwYlFsJnHcLQ7rdo+Rr++hYoO2SltdIKQUta9h52pUcJ
SAoSXzSsp5UWGgG8YdGqaDyYQGY0TKZ/8WGu7cuZiSha8WeoDhK/DTA1HahQ22P+WzLIRKstpoSA
i2gJJqk67Zllubbx9o5+OivCRLARJuSN+rC/Mn+Ou6d1z9A+jghfOQpFBU2vgwJho+rCgXGIXqdR
0gFeXmGiEoHio48P4WX8WMzswUWHMGZ3i4Ow/M2Od2ETEVZgmAClE2GzYDXxzpV18SVX5IfrY4b3
CBBAD4n5Y/dXI9VKUiDsxi/S798E9iTjHi8v1Hq3R6deWz78LOd9N03969o/gP5Dk+Un1B5S/IJt
t5puZjoswI8/cMnfvJL+lwCqke8h2iWeL9BSGM7l+/eO7EckRtWyeR1vsMS7ksaLo0Ghnpvnv+dm
W5epRC1rHnmFWXUdxq9kqDP7LKZ8GZWIy2b2k5ZY6RPSKVAkD1muSo7QlYEiVUcnZhsvhigZjm7x
qf80zllQay9TI24aDQKE7yp1raBkeNPy5sXz3m0HZMNjb88eIvP64O+VRnm77uiKn9YPh30Puzin
ZhqjKUFrayA2Mr/KPMnBZaPx3dJSEf8Rl937atZDT7KEvj/CuX77J3BCj8xH7l5l5a0XsNPl+SWF
o4Ow/gpBJRGZ62cGW2+LV1u/f6MIbajYrDQtxFRUYzkA9mKmk06qgS4/p2QIeJ9haZK8VefcVIzt
PYwR8/JHqSTYz/LY1rDEl1+qcNKB3f/6VaoPaZJ8WVe9f4zJN8QWzZ+9d4zGGbAmTXe1iKVLy9gG
z89120QDFmGuTvyE2q+4c20OUjd7euS1cyElFOdUKeHGNHrdx71u64gq3WMZ/xvoKL4weBRMJFYs
jULo9OHm8KUpsbjFx8f0YRn4BMdtH899yHCblqdThWLSITqHDF0Pxd3OEWcl6Ix7r5XFelM+VQnj
84Xsx58ABX3p+zgVdT5lw3V9/RR8JWssdCIxwR90fj4nfPlFh2vdpNtBGuUvi/PHOrfCGxDkSF8B
CT1sZrK+MGxQ9N/zNYbOHkXGu+rw6RXADBZziFjeyXnCsiU9ycNUN2XIzyCIj2hQn0MAhDZbY/f+
Lh2FycgW3WjK2YOTqh8TVKPLnMtOMFVjoeiw+KnulgQKqiRO/dMaq+VEDSQIYvfsxVtepD958vGh
ox7ACT14RkX+/a9aDF6F9Z7zU1p8CgLFW+bJ+3xrfsuuYDOCPMkh0TxALu4u3vppkYHPQiXAUyvF
Fv+qWvyvcgrZwEInJFzcqQtcYu2xWCC0jhBG9wZsPHMwf+X1RfDZxYktLru19NHz7kJ5a/71PMVB
u4md3k6aBgUoK+fU7bzmidAcwsZxXCs3rZwiRdyBvviqTpn6/Fc87mBWmtXRft1IdpWUe+L3Lje/
rniPN1WCRUEvHtn6b2j+FF453yCkkTy9P6axoIsH3nWPRXVRySnqDjI5Inv9AISmBp6Lu9t1tUuc
cG/kbJcyMupMJzSiS3/RkI6EHzF2kp3Fg/0PA8ehnFDs1HBcXJcju/V7n8cJqSyu9boFXseQxTTh
OVqMcBzPzk4vBFtnuOoV/S76p50vMpAAMnBq7Uz3jo9+zl3j7dKhtdsgoOavQYuKYqrPKkTreSNi
p+HldbLLcw9P/BStFUuPtf+mOghHjEPp6VBn2BUx0s5CsCT1Nfl8s/1DaC+4me506Xo9e4VME/aB
3yeF7uG1iRUn7k0zqDCRkfA4q5VbqMQUn7Nhg649NuMPZjbTMsK2hxbCgK3zHDq1BLAgtXvXsULD
qQaKn1n2iwB+WM+sjHzIwGyIvsfekHwflx+3Ki7kveh9mPn1AmBnN/Iuwa4D8125dI5tsW13k14D
f21SuRiWsj4iZR76oinD6t20XuutoNs59/XHxr2rxadMb35qOLweVQz8Ym3Ow2P8XGKTwCT4EjFR
XxpUu6khn+bRK8K8NKYWWI4P7rkopRIKVJvuBczx4jze3FP7Tnft8l/4205kKfZ0m4NgLVfpoz8f
6gvS7bCFujhjP4S6njDyqDS2Z+kk4l5Cd/06ze3lf65+YIrtQnMnmEq+fv+G8JldDpjT28KS6XYG
0QYu0uukhtyc4s51g36UmFMB6mKNOGtHZ4yC+vYGvJVoYLF0qRw5lZzJT2acwWo5Zq+yhywDlK4l
vh3deM1+YOvLPYaqlIIPyXPSAkskblVHihLfH5PYEgo+dESVmfJ4rmuNgc8RNb4aApyyU9S5PSsk
UbBsLZ7+iDmdBthiqe1xKRT0CFJuZ+YAJvm3DRGtSHJQi/36ufYwutacZb2y4LbIXgi+FKXFljpK
NVJC9qGy85yYg2dBNNcVwQfpzrad1f+4TqREFrHWhaYUOW0FMjRrtcQOEdL9jjut+mN2m9keqlFP
++a94ml/PEYjbcmLTNKr+7ypnr9XoLwCj0+N4kUwOj7jDJ6AReUuBDVtMgJsQto9LdLZe9vqit6Z
A+OrucL79Ut6BAVKhAMuJs0lxzwZLVvOsVAStt6VNCc9bEpcAmN7xlONYoMSNPQ1z6wSMH2qRH3i
ZIqoJy/MPyUBIzrCpARGzcugz05COwLuY0gNPhJt+0PzbFoEH1qYksOhtIXzHHpSJRhH1FD9lj+v
vBXvm4mViBJV1McgyxMaZ5pBAoG8ad+RILahID/sPl917nrAKRzJ2cExR5mv7GI2adJM1u/cVv6a
ze0Z7+tOBTTrVtxVKBCxsIAong5LKntpmQgClMi9aA7FSIHKRXNGxfBceIJkWwz9HhhhQNXwGByx
DwDmES/a+KQctFjG9Z4javYgbXCHbyDs3Vwment9XRpAmlwoAgQR0xm5yiutxpxxdYHrSLz3EXf6
hVJChFb7/ylm8zztccLf35ZI5h09AimkgdmbuuMXEGsUyxsEtkVfngPiZWxXJb8CfomdOhN7XjGc
SE1Qrm0HCKl6dQQ1SUEm5CWjJodkHYEs1eYuVAi3vsYWbJGsJcOzsKNKMF9xlk6ps8/x6uVtbOsp
0tIJixICW16TXLSDBgxEfPIGho/WbOmr/Z3Pvs29bz1IBcxzmg4PAEZXj7De7PnXZz3S05Qbydyk
ozAmaALTVlYK6YouPNUqBAa9e2IUuinKTH+pxnH9cxa5nXK1ZQuT8pPVV3uHpMWELETHtkz+tqm0
IJ2ydILkyidP3ukXwzyMgCOZZkcggU8Wr1LqA5AjqA/1hrYC7wVvua8x85ibHmeuKwm3G43sg540
qFmllCij7XlWQupvKkYDwhPN/RuJfguF8zrWsL9I1qrkmoWO8xj5uB9sFZkrlMhu59sDk0RqM+iY
w/mN2nUtsa9crqWcrp4bPE+44O0crudP9T1ypBDBvde+MnrpdcJFSuzzi6udmSHaKsQJXyEtJC4T
k33zWqz+f86q0UWHlWybjejCkuGPi0hSGXDKA/8nofhsLO6ebvAYFL/NSZBR6ZHzdwaPQvb8w9ZR
GN22K1ZxIRMLE/65g1+dtO+sc2dL9jKrwPBRGsdHOhV4xMzpZLOrQqfLr5AC/lgLRb78JBb9hUeB
m8H5kwLfIAttB5LsI5MfPcFJo6Zq939AcoqrcNhl0YQ5hiTm7p5LB1nwEu5uRcbIZmT2Xt2WTYNo
DnLurTjzrm6qJKV04rNUmUCP7RML1nSi4YYK9Zln9kvt1Da8Et0IRX4L6wlokPSAWhpa/ltWursH
AXKrZTROJGC22udJqz4KNP8G/QhRexojp8Th5kb1E8EebOZBFbSaRmuJKehhnt/qMg9HXc/RtyAj
VVI7O5RtZxaVbyuhcD2lAx8kcCv4MAUGwRP2wDLzFpGuBcSOgaGNN58iyU9M/x85cPAu/l7y7/7H
U0FpksUD5rx4PISp1Xj6J8FXMe1IOAKDOhEBP0ieQtk77/oKUskvXbw8RfDQ3HgIcxJ4oKWq4NHk
oYI942NrbgSuLA00ODLzbHSh7UeO22Kkl/iabjtZUU7Tb6v6ZR41a3XyIQ188uwRoUclSKIqj9GG
0uhb1zzsJGWbMvUZojHtyiZm6Ki+Ajo+J0N0AvjdIHJQ8oh7sPB8/oxXV63DrzSGF0KLXIuB5R0c
+TBONS5QBYL7AIPB2I2EsSQMepiC7t1f2EJLywr3Tb1C3+imBqV5gc78WODs8Q+E7kZI9Kcxy0so
ssQK0yDnBswH9LbhgUcR+CaRBtyyFB3dbR52V8hHuNtMP8X9cfK9GL78QjSppq76N08GoWHY8Wta
ub32o0Lo8DgWdaKoSBU2LSNScR/yQWl3uo2PyhU5qa1wOuPz4kErU5ggNGkOjGbyBLQA0GWCs388
Q9ms3GDDzzeyxmp312xcBULlydeLv6sgNd99TSx7wwoprU50FZgwDxrczG5GPEI6KoiUr+HvPTmD
s5G0aduw/FpvgxZzjTxWLpbfGxL+hcHjVKxe/+AD9OqGPMEGJ8zs3YwthV2GZA9j0nFo5U17z3DI
pXDxz+5L2e8rIDZTQx74gzSxht6RC/SyrP48q9xSwKE2jztpn6rELXFlXueKM0GQOb1lxVFxVTDp
nxVcRVE8i+9u/zh1ZvucrRSMmnvK6w1mwdMVFzHm3WTyAcZatmcJTdO9+fNHKUg3MT8NNx8YcP1J
tY1xaztcBEsgI6lFtGIXV8IGtcf9uQtd9wAY66vPCZklTnb4zTg5MgA34pVJxin5Y6fpi1d4VBSu
yribpC9xj1AiLmMchtl5sLVSMcuvF0Rp/DnSIcVa0VD6XEdDWb2sjdBlKYiMnzECfFyX1cJy/lSv
UOMExF9sLuyV8pjvsJ8rVj5rR9Qny+ihyY6DSK7L24F/OKN4IhRLemY92T7KZQTUsaz2PdxdjOsT
ZZYFMG+X+qQy9PMBbM9E0vQb9LJAplH0wmsAiV2tcjboUvGZQMSmYNTW/8SgoJe9MhJvMkNKhEUY
V1vFy58PFSg6c2Lco+VnOkJyTxVRjELb5wflc3fezefVTCmUa3Ua+odsQ80+ATMawVkhnSfY27Eb
x8SaaVsuM5aqR2n5fG6S3kDXiCVF6QCXV70+qf/N3BKkqyBeIdPdYFCswaa7E7iOGju4JLrjshEa
/Wa73mcTVKrVI8o6FONwY3YL7ntgn9MGWe4dRQUOcnx7XwFlG5m0B2B72o5c6uiWB+ROjRuGjfUL
pc5wZlpktGTXncFNIH4b+em9y1MK+7YKxSIETh73gHT8k5XawDqthhR48q2h7CH/nXp5KzGpW/Ad
NbeB2oXuknjySPkav4Enr/Z78unfXOgnYLeZSt7bv43Wpa9SUyPJKayb1rzSyTmp4EvZi9nF3LN0
Jp7M11wGvxQlQzqwpA6apo2w+nz/pD8CY13N8cc1Jvj9KoR1XOUA9Bu2L/1QSgK9JguR6JUIPcXq
4q+cOzDbrpwxwU7ttc0b3BrciQBWgKlx2zOZd5OhzpXwJxfKxW7KAzDQnesTlZxfNo8WIQYBbSd7
1XYduOUhgDjBJxMhWQo2R6FXMTOpsPo33YZ9+jYH00kf8DGCeIR6yq3S8m2/Lbonlbif5CHpbLhe
xRWgzavK4ljmAFefhi4zcLE64Kgi8tC4tI8JM8flqL7UgMMi81sEv4sFniWgdSkmcAjLQbamxi+I
MhAzHn5ZvlTAq5ce7H6eR2xFMPQEdp+uMrX673O8iwNy4xFMldIkwPFfx2Og9HdEZXd8Dy63qTu1
cSqZPrVxDZYKMhJ2Igxdp8+PHyFqUMwMCsq4sN44y38QhjYMd24SGGZpws8EPS6/KUEsyuVeZB3J
BAHtvOwSmj4TALQt2bY0CHIHZIkcYkcJe4bcEt7GaBMxYmHCN+c4Ywh8nWQfHbpeerzInE8zXEyk
x/LMYacPUeaYBtnO7YqJNPNRX9qo96qxs6+wXwbQYeRxiY5C6gBEVMUdNT+MYlf9BfV5Qs9prikM
vW1bV76InrGNGl60OyTAT2ys3ZddolbyTiorsVRVtDVkSexOfJ4NrCPGTtDbGpMUiv8N0q57npMl
UNFQ/9DeGAvrTCvohknw15SghpIiPK4qCRPiZJ8rr+y7JitYLQb6qwG2Fu7IGl6TrIEHk3QgzzU5
IG9UBVfQRXlHhaI/GlwEmVmDpRYbYGdfWSMLV62jFVDscYb5kuvVkk9j7KlGIma03unfKnQKcCsw
7exWciFxQx5QqQ/fLumUXp+MZpwJuhiaTFqFwWGDzD6jAQiIDpVsGnGcCNYFZJxaZMvdXPz9SKuT
6wlGUUZrn8+Wo4KG4a+4GjCMW0ZHdXNik2VpzdM8s75jvCGe6D0Q0rlSKt1uHzz4uHXn8V0+Q2qo
PztTFRR8ZZpUtQ/x5p4eBXtt1bBdsjudVNE7KXLUR+ME+pkr0U0HsJY3KTMKYZnJFB/mFYbuPveF
qoE/+/iZXBvmmQQX6UUn8xOHDIx+hoO8Ge1DYpMe0KHB09lr9iadmSmkMSHJdMzdTl3ZUr6iMpAG
fz0AMWhZdTzApontZxpaEDJvWJ1a3gMxP9z/1HtRADfwQrX7fkTUuwppdwPDj4ojEHXyW0urrlSI
cQmgTEmqq9ZTyRfCk0mVSD0U3IQ54npGZC8C/X3p4m8JiR8c4XCysvhH3rlORjOjG7+8tnnhMLs2
fldjOGFtSPku7LMfs90hXmTyKefhaKd6J4n4RCcbwqODX7DbRxoS9cQuuMRis2s5uqNTtrnDzwEh
TppSE8CAu9s4QJ9oJDWbS5gszBPSApgZ8Uc05eqFE3ZqvrNXbgU9g6WQ/7IRcvGOLO3Eb04Wkllj
AJH5QGC1hb1Z5Qjk3r0Q4AlbnW2IRDFXVByTnRO9NaZCw4xVA/Re8AJgoFf5BWMlgaXP2TpD+96L
d3obbif7yXblJaxqDLyPYT3ZalZfjKcrv/ROz0sPWNAoTGsOBSQBJayA0LlqaZVlul1AesNDBvlU
v+hdabkVsAwAzRiISdTQ7ymjzefoOSjYccHQkTcMGl9Nx3ssglxZaQSvc1hhKEj44sv7oixVHIPX
hcxMOAQIGJhQ1GyEHvqN2A7j7sfWxXIXXz76bhn5UBrY1AP1r/RL/XJ2ObI5bKNg/Fnewn0OsyM9
l0JMAQxiowwgdSXdtHcQ4rb28Joi3Sqfbtgzji5r9wPO5ZDQMtSTFkR3nvWGhUdhc4JvCXIvlkI1
A+5XYZfOt/T2oGDzXayNMtlaKiH7UbBPWfIyAis0ltx+8lXAQ1nYGiZcociKYFHskTrjWWpoEBk+
dX+q+qthKJlAaLrZnvh7oi32Bg4goKTB9p1vm2GUYH99IZEMKF93iVRWRIYFLcMg+rLWZdZOHNNK
3yLpfh5sXTfXtCzX4fEiAWWd7dfwsN05HQMPCCnKM1lC4H/wN/gMuR7qX4wkXlc8s0AclqAdUt6j
aMxQQoWMjFZ/CPywUH5AO0UHMQywQ4qfyKM6KXGqrlkriIOWEbFUNB14o+z4Dm8uZB8Li4rfQA/w
6qTRfxApihbq5u+MdzMJAEanAvUbbBqbonFqVIaiFzBfj2tiTQW+Jr6whLxuuGyj1mPJXiPHaBIM
m/vY3z1HXkCiFc19iK4doetUsCf/Zb6UuP/0Ndx+By82sahxtlTB8aXPczQKSNt7MP7KX6IuMjvL
vUodz37dZrgbdFcnUXGReMG5DCniPBXaZKEd4IUFBctVSz0Z7yZrOrdrWg8nCY2iOyEFN5Balacw
tWOSInCpkcv1F9ri80lCPl+HYA0S/vn5rD4+gVszTwja7JutfwVaR4oTmjJ07Fqro28v3oKgwsiT
aR2yerrL/edvZA9SsICCFzjfj5gxnRqXji7x/bEZLKwcp76M45cjiPa4Ot5NUjFYZ0f208speuky
IKvqelShappqWe/MpSWciDBJFjEme8EycZpr5aOP+j+9RlgJDZO7Mz7Q0avJ0IB4Ck2eq3Te5UXT
dq2oQmsLs1qQNb4KTQ1LSO8KnFiwSudLsXE/L2z1uLWYtk6S97IGVR06mKDYD42hu9/sPb/heYkf
MqzB68lMuwPLMaaO/oRUtzXmccMO27LKDosA12D49ySAqrSMZ7UM0ZvEJNTaVM9BIk7Gfj0Bhwkg
mEvt8Q0WckNigXzAuptX+qXgtDQr2gNX1Z1JEtbMZ5slKQodDbmVnKHWfqZW/cx4AI26YSKpiLYa
xh2nPSIUtHL2CX3gCoTJ8Ar+jzd6alnerDcxrqQ63QDeaPZxzcJ5j71FkYWLXJcACYyVpJ92JYRB
gb0/wFLj9Cow63aA8yWMW1tC2pGoCvkns9SVXcQXGRjDmB/7Uk9siYSmS8Oe9C2fdoBy/9pihPno
a0dyaRvQc6qS48/+lLEXAqF8m43iho7GQsyVSx6cCwP0POe46OSzRCEFRcYIwHgGyEDYOLdyXXJ3
i9DzWiYGW9VdRGHVc3zyhSDaOpIyiw818Yp7Pc1wPUuip6EzwGpCDuyHlJ9p5xrrenqxrbjn/Dgb
zVaCdxNpkUjX7wDQAMMIsIS+f5wLjIyqhLCRuJZJ1uMw3zQrfhib6mXMbJMDKeqSMOK5brFSTg4v
FN5T8dcqReMFQv57V6lMv7ag22+EYD8vtA31JKSg7du+fqQmpowMxk+SeXr/gDN3lBy7FSctyzid
whB2KRCwx04A3IsyCsHYPSz9bm2fuVzUciE592KE5GhbrhqHbRxQnT7POJmIQczaTQGH2dwFJYVd
P9jjPfX2yIrSx+i+xnymzGSGo9BhssnEucIS0VpnFckMAIHKztM+PVFHAexOm4PxpgkLEZiy4sCJ
2XDmPnKsj9P2s+89LO2ipda/JsnMpBq4Y2hMaStXDlrvdt6nTAsat/07QfaEKqZjyuXdmMnJXDeG
8rsc+u/rEB1ikIE2HY5dRTL8n8t0E6bT8eMnhXELxX/VtiEGN/PMGPOzB1ToQPKe/DOAnulTH/K9
5/osmVa54hwzUtmnJcwCgznIA/i5AymhmFun1ko8AMy51wquC29yF1OYHfzmAT/LlESsYopbpfHz
eLoSZ8UeN9LBNHsptc+W73Gxa4bmWelvCjH/hbBprvJIop4+ZQpMJm6XDMT6bcY+4TFtgBIo3ynp
bDKVQqQrzvCSIjxTnUuR448/cz/zBZQ6P1n4hCGWvO4gClNN2XUUUrpp3H2fkPzugZYcmr9SEV1s
auRHaQ4pPcYYCdBgtfUPNkcpfQvvM9Rh773apIkk84yqIoPVoPhceXChlRAib4D2Jfqv2LOZhcxZ
6gNf2hAKnnEv/5XCWV/0kADuPWrDPHYqEhtGmRcAx2ZIzN+IF6q53VV4TZXIkr/lvbyryqsD2YtY
96ShJk/iCEfMiNpSZJv6BG2/kVrZ0yZma0jE2cgBN1zag9Qz1BivlljTlD4SuOF95bKN3k+bVcHS
PsPzgyvBgRafzSHWjSvYowZOqLN5FPHKJp1xFFU3zEGxh36UCxrGaxIl2NbjxZgyOuEiNbiLshh1
/Xfz4x5eHWYRu2mmMvQkn7X7+w33CAxTkH3Vxqcdni9mwTj3DSdj341fM8Wk7q525w09m4ise4zJ
Zqpwd7YHGiy0cF+8eDSkTjOGU8Ih5ww9QkygFd20+m7tF9VRxVVGhRHKROwK3usIt2DVh6E549gg
tE73JRVlcPwuF+EYZJVLYj4r8xu1fWYjqntFiyvcR2hWmFbr0/p9RIRXFdCLA3gd3Mc4/1drW5uT
pZmrnK/akZoGpR9IFlN4QlZs4aH7XoqzzJ9Umx0JnYILZhQoKMXPqBSInKRbEJe1HIgv7a3SiovZ
sCwvkHZAq67tBDzMFIW44NGYsaxvX/Nr2aueANYwlo7TPZLvt18+XfM2q1JBZHQs8ffTBBmTzD9Q
mwxGDFFdpAzSgb4Vtins0296KGXKgfWndcaXid7zSIlxUwVEyLsYsiLnLIs9rv2eU9MQE1zpltCI
KcAXOhncROzlHVeYr2wzq8ZwY1bHz5zenf/UROPQVttALG6eojh3qCCU2+GQ9qRofBEgXBO+FDFy
+XCA0Nrvt6maHTonUnYC7p7wTHNIV850lsM1TpEHLuWgc6GL7Uhi5gpYRSE9JyCNX3wJEk4/nSIw
aEuL7zt1DqiIWnXbt5G32Aa0HUGW22a6mp/LiOLfjlpw4CSivyoSqaTLJ7b79ONoJsd8q2zhAX8a
DshOXwrohFJmdFy1yaV8Ps9XxeMKc8qkC0nLN2un25wN7WB6TaU4tBYHhysIjRPMRuNSnx5m/lnu
yWACQalkfukFPtA85KfGxLRI4WYTTQxuH7I/twt7mr/BS2eLn7+3kB3/XPqxbzLjTrC53DcNSNmt
UGeEbUL/b1Wuy3zBdCWmKapRAH3jyOn22RqqT5Q1EajkMo2+A1eFmHHi2I4V2Zf71CoJZFIM+w2U
IrhqbfoJDNnOEc28RToiP0u/LrcBljRu7kbY6smzp3kjquas+ElWK9WW9CStDyJx1PNb8d0gUZ4b
VpgDEMDOo+ROsjM2VaWUsD1CqnbMsIegVpvZsLuP0JG5vkyrohkSsg3RdjdY6eNuL/cFcPIxkN7p
3kXrfU99o7oxeCoHraQ9NwfFKtJj/fOjKiYi7XkySs6NwopU9BNNsLEk9b8GKUAqZQMO+5ACY7tZ
SPaMOo1jV7xDoRK4id0hHjhlbPFByPqvyKUn62pmlzD9VUKpafUUNKWexeXGnDEUy3oMkGV5zK6Q
puAwW+iFnODh+JyWzYEphl/pbTMQstadaYs081Jnj4dwzETyRuSZWht3XbmFT0Pgi7cjLjOyuM5y
FTF1DZ2sDWa735pj2q0W4Hw/MX6KiPD+tWjctvt0cX5E1Un5gOq77G8XGUHC8jrIEfWYazdhTky6
W3ahTrCuCEVIFrJscX0ghNgzSwNRSy5TKO8C6eMOY6wK1JQxldweeN0p4D5zDNW474KK3WcOrnqk
q6SngIv7R+22YO3yuIp3Kk+6SsZft8dL65IO18lEe0qjMNBxw+z/hi0WDxjbsi7Cjspcuy16trJ5
pTARv1zK8AqTmd/BBu1WZO5TqPmIeWEzQExWhnANEu7zA9EWMRG3E7MyqYzbC8LcQ8eBxwajOXuh
IZ/Uay1I4Gm5reEcMbOHLPm8oTFzydXHTywn1Ij6o8hq2z1tap24KILaIa6X6ahUS3JS2nuxPtiG
drTFt3kVrdhFQAxvbW9ejqWTzq2vkOnNfl1YyjnCB3NiRCySHpTEdaTLN417jvniQTwwF7qrqkff
lar+b7blYZLVbTwtfyvOo9HRBiSh7kfajk2MIme9oHksWqyg6tMWWtyRbO7CWMYxamkrSPZ0n+uD
2LARf1IHAG4T2Yi6PGK4rRxSBTbwVZpxHawddP737doM5sj3ZCPD3+dqHy5jJxMOWCeyiUi+D8cp
Xi6B21khd54E3KW9Np5WkSyh/4RprKjJzatIRoo/NZT8XjGj+JeMjMWJNwyv13N9zLwD51v3AUwu
wFG8NXNqTBdwFw7DbZA9gNNwicejKuSi53n4uB3cSQRywzh/3PSblyWkQLtUVub6KMerLRRO+PWh
HzhxOR37AQ6uutqwSX4eIzuzSCxRiEfr5ZdfRea/1OSnFpLybsKG9gzMZYOsBQv5bkELtsBAT6G2
M/iIJ4OhIo7feDwXw4UHg3nTQeBuji6BflucavnPSYddxtjHQFS7687I/HS03NY3VSzx4t0BuLZg
PsAkbDe9z/teFPMVei7uND7QBzoM4UYuaikYzVQFItrAbTTYvtA0NrFoSc0QZfaJjUvXxQkdfaMl
oKhXCKCRy6RoDscESWUZeGagn6vLVsG34MlfYg5c2XMqpH7tA/DaMnL9ydWGNXEpjjAYKUnMKys5
/tkaEkE8mkhAotvawIuyMYQtn5/VnS37JUmXApwsEL0ec+IIzyqPCPpnoD8TlkLhrW/adFoqjQCa
oyeOaF2ATJjOEIfAVbftBw+52/CjqaGyMhW74YVntuz8OqqAFPjAM91ZwmTP9ERQCosL8HHWFO9L
/icSdQNipCTUDFRcRQf2NHLX4CrV3Thq71/wpJY6ddq2OvWzMS1rou02KQ/FypdK6cUCvZXx/CQL
wzzlsruhU/zcWQ9l0T95wUwBDSHhCCzKazdhqD5FzNrCyYa83OZ4F8kXb0YrfbSXrkOIVArsF9uN
WvsyHj+5ZiK+WYmNsb5sC/DRSdtTHRjspHnSDWRUiJ+qsXv7i4vpRrBt9H+ffIP7M+z6O4A38yeJ
a2FNweao2QH9BB1tVdOUh5aB9/Xcsr9E3zohfApN/T6ppYsTmI1Y2DK1PavF5u8E+IYPfMqKF1TZ
mKix4hKEd0OMfY5OefISRtC9Foi9t8iWaEBXzXfj0eZrO5MJ/OvPHV2L4txQeq43CDMyTulWjRMf
6TJR6mVkN5Ow5JqQ80F8Te6gabFL9COw/zHTCHt1XuDBaKzdUlQ7r6BqBHMcOhGyQl6cGctg6V6r
OLvolR9MLIAg2pVnRGr8farWeG67Gs/IllRa8RegiC/NkCIlJ29ZTQpaz2LSmwKk4hcqeHAo923G
MNJEJTLFS7UHIeqwx8r/aVdGp4CjdsHPxu7XopCk6AtKrg0qTZPKVxKK3Rs2iM/DGejPfI0j83k9
r3xkw8y2+N5fSxjV5UcnM83PU0nj92lY3R6EujAxhn3Mk+Aid1aBejk+ZmDW/F+W6xZK7nUU2SV1
pvBSae7mykzfjafOWoVrDo3JKHWbQBWJPImPdyoO2rbbavIt8wAUFNDZGbPHHVFPBIMqjO3g4fS3
eMz+qD2S2XCgdRGaef4CShzEpF6ENrInpU8Y3R7lrgqDPeiOa5oYTxCDHg0jh5lx8I2szwoYMv1o
vfAALEET7mqK2YnV8HKG2BPhSqIvG4g54dy5RNaQtdlbOPmP51sVZn8OLHLTMet218yItxDd+7BL
/6ysYyxl4617hdFC2EORdjpdjH7tX4/9FYrSsB2hgwDheK8MiwwmN2gYkqinPHi2WLm+fJGyUkLG
eUMhSWWgnE09/ToVojR/Fk5HDcuDcVWElcWsXfOLp6RQhJsE+jS+I5aJYRDDVPuRjrAGkVN6pN+0
CSziN8GXXgjqIKazytNPJtr5RPYlPRewTWxg+Kd2SvSDoFrBXfaSK0abUgPf0v1YVU57BYfIoikf
ZO+JuYhb1mbeB8BX89j+SqqmshjXpQ7E+o1xdUxxAgwHoHkM4QDWQ2HXr24wqF8caaM4h4EV3ZmN
+l6LseYc1kJsCcOBZ0T/7A7f1agPd9M1FKcRorSYuoQ+smkygwpRvc48LAE7KB7rt66LMVZCNEhw
y/grO7KzuNWscoVtZiXCsbsnSmGr9exq/InUXl4Q+kP/8/RvkLurW8AQdeBzAuEaRPYVDzLk5ZNM
WU7QxqlmkpLb3F5X6r8gPk2bsl58fJcemyucvAjGIOJuVv1yQsn2eeHoYCosiUCikz6ete0TN0MY
PCAdqvxDeMow6y0j5gdvvMuaQn8+0LrzfGWDCc2Sswv6KN9nV9gTX4PqS3OelU2PuLiJUkY9OMRq
gK5/SugxqMXwuHxu6pleEprppqMdQRdrTw3fXUV7+nMHUbhV0/qhnK9gXOWVidVzBZge4hp35yTo
eLfZy9CINTayOZyFOWBW6oEU3ilk0lzDMTcVkjjtgYKI70NXyR5uSq0vzv0ebjdp5M2bpUl58Adg
n8FTyxEljN8BV85WMYg9rhfDfzEuTeb9/sJvM++nGRS+NDOQdf8jWFBp+/oxxdEoiWJBtwIHNHuN
F6llS1LtlnORG56zYSv3kcb4yGcuATXZu57d4alduOeUSsUy7QxzYPmX/Q7/D5YkklJmou592Bqw
E4BU82jcI1NrB6j5tKs6Oe7bsSoKE72drA+fziqx8l+T9pIVpzd3Pz0rDQ1N0aRnyIptxdC1dyeF
/HeX1C0K75b3kNqNGhoIlWLmQ2j06PJ6jMtticHeYkrYuHfEcvzNjn1+G8PDTsVhSGFz/BIB42fb
HO3Yd6gV1MZ+CHgm8JOBUcdibgjP7J2i/uB3PyTYqOmoQaA+ouPu8BPY4GtBjOeoGcboNrxpxtFP
g41ljR1qDhgMswbN1xOA6zbBEEmeonJR+2V0XeDOnb3BtHc/9tWesArnb0rwV285UNun+w6ISE5g
7j5CVFyAtTjuQ8rRBtWLVnClJ8Ok5WjdbkTps+SF1jAEU807UvrE3jYgB/gDzpcZAvz6ZJIY3Rxm
PgLjoHGsBaWni3CQd4v3IZwBAplGxBLVoJ4LB0HzvOHR1tqjlULNbfFfa6KuOOS8WdK5lUwdZHLd
ovT9/rOmamAy0aY8u/fTQG0Mguz5dPDTRyXOxgwL6ymP+d0pgSoBhnZtefPNPo2GmFKIemSmqXkj
RlbGGcL3KOql3HXaFcs4UJTDx2jk1NO6k3c9KjVxPI8p9FIarFikXZq8gfJcFqdbUd35GZu+7cRd
M/OPK8uYJO861zsQqbFnp9gVNzJ8Q5gyIRCW3kiqCQXVkMguASSf84GHtGGQDF8mWSENouQYmDvL
bhJ5tLgoelwb/UJY+SiMfBIC20Pc0U33C3lsCL8YpHAGEhFVjlw8zNE+LcRjpsFdFgqe6Xdn8f6r
KHbMf8lSAicq0Y0TE79lFNQLYBQE8ktnylFSMFaJEzqFwbIOjVB5vEhb/1EQbS+XKhVl5Z/bICa9
RKvoQUkDfUC4awgb8GrrE3lGrEZyBwcihR5WJyEk4bnKdaUhxDEsXUxCD2g4QeaWTFzB1CilPuRG
MVtXxokzebSI9hWbSHqaDpbcgFftn28SWa9mPRwIpj66IlEV+Oau1GL39kaM7Y4nSjTJVsGhblz6
16fO2n0bRwbiWFoQHNqr8n57bIfqpc146nc3Na4ZXnMUB9uZ0zn2qbbouZ2vofgTcMRa35qXva+X
0/lBPg2qchK8f7V/2x/sACTdhFYes7P58BUAVDkhsACG/8u3OU2rRKpja6qUaOa6jkNapEbzIVT9
ksluAp8smXU76OBgsAHnHwjcTe4iV2BmGc3PN6fz7cToaCs+2pnq+UIE6Vm3szMlOVY+4zAfemCO
98lQUpeMMjVP03jB5j3dSY1WdhDiJzzmYDEtpLJjEoceeacmverLWzDNYI6w0RjaQOxrM5aKnwiW
bs/rfunW/mvPD57q++PocX/ITvaAffCZ2gcii1qWX5vPePhAkQN1QsJmdy2WhUvMIkeJ4v8QdJU4
/91VnlxgtIzcFIhp6lbhCcZRU91Q55uDcjExmgighET2bnXevxTQddUaeG4VzF5EP+ofZkFPCnB7
ZYFsEAz1pOor2LjqHjOcaiDMCbsCPpvg/uCrP/HeP7lSaVRgSmfp5fC4wMNAL94aU7vyz6ATPwFO
uoepDfUtX9RSSOkz4/55wQR5Hd7jSLJiP9gn0VxVGiv8XCZxuCpLRqiPSMaqJ5464sbbutvmtSll
m/qkB2SvgtvpZiZBdIRZo8OX7Yqsf+njGBWpi68zOZvPe/ph1zlA36+z9/cKKiwWHNk2y0DhbGRx
nsHpIT3OsxZ2DK6fmyx0Z+NLKJNh0ctF8OGxP7nmfLIWeCfMROcZDvan1k5Xb2F8CMnFp8KSuNbW
vZkoTuF2p/Pij7JSj78rAEUl2E9TkidG84DOZwfSSyYV/iyS3kMk3dEVGbWaCEerrCZIa05m02Z4
RRyz/dg3oxvBFW/eTGJxNVSevOP8ydSKupJD9KLMWAhkHpDVaUl3Rst96me9cM8pmyjKSis+sh9g
PJnxAAjq9SrL39VpI/f1QSgHF4148ICR5L0tvxnP3oPd0vUDbL72ZSkLTfxEY2M9Rk0OWKmcRP8v
1igO4lMdiWKruzP65o1zvvTkbw2AWF/N5p3FvKdIPujm7KreJBkaHyq3mElqrDkX5vmIA5CvyD1y
aiZdRZzUjgsfza+UW8NRPWev8rvq/jgAapGqg5LDh2Y6+jWmwWZUNC4b6edRX/xCvzxvz8tK/yfs
f4l8ouwi13jv4rWUXd3V1OUi0vsQWkGgxL2PKvp/MzxSlGdHX3ufqR+1NGfph14/WJZNVWfjo4is
eSAxolra4MVv9UFOtRlXiUlwhVM16O/NDZ8a2yJcyIZpdQT52WCpXEB8b2uz69+0bRTeb1xnbAMK
3pDrMnHv7i3hov7U7gEf95L+v3YzQ/UEGbs4I/NsE37j9pVZtOQJwx1TWtAluWqFx6WRSp4WCVLy
Vvf32BAlFkqIZTidjraJ1ctQnERaU3RwuZhhJmHZrwQBm09EpAu7O7CkUvXB62tWumytww2XqhLJ
NtJVyinDmuncthBcA+f8hORJv5Eah55w/x6xfJnvP238Fs68LcKILttDH5pbNVUMKIQ7jYUbnh7i
77EP0zTTnUNtVFiqsrqdRBA7aMw9eU5fBpF9Vahu00x6NeXmRu9xFg5A8hE7l4TsIJHhrHLH/xsE
eHO6cVJ589o6uuPzynYtEcpCQPquaCt1Ue+n87ZG0VLBpBGyKvR0MCBLpjzlNMoY5y21txET7obF
bQ1qF/sNQsx3PR7k7iITZ+wdMtt6+Lnsefp6cp7BK9Ip4HLtQRu+hFnBzMUe5uAObqgCrkAbVh/4
sedFurOa8LhlmcMI42ZAh1gpq0Cm7bK5VjW5Nr5EUfWmldP+ejoW/02U/Zp7nU++SXkHiH0WSw4e
ZscpxvZbs4fybJb4Syqy+/8aiSmQ9TQ9KgZCVUDlCG/xFbwN/4F3oE/ZeGkam+iGA7UZKMIhHz/T
9Lbo2Yp7g/6pD96RsDPK+dEr4wY7qgamG1MstyR7XxwT41TMFl3svffLEwKYKvSxyZpZNszwlNEL
buRDwlpiyke9jkV5uBddEEMJwoR6MIfEfwjnlgiZiKLd1NMXkoQniFhtajBhy10LNY5GOaUTPQHY
WxE6ZRNC9+KIphHNIl2YBekLVney186CTp5q8hI2IWm16005g6rya3LJPHfqvdrLdMddVTB1uzd9
WQ/MWLKjHzMzwfTjoPng5mCZsBUSAujY3CxMNLPQIyDDZwVd7dD/U3vIkvKCo1hwcYL5Uktj7QZw
1Ep4/SnOZGAkZUyGa66vIANX3KR8E+Nd/jdVVR/fMUbtT/3qx4AkpeGa52Y0zshoudYPGvYw399K
w730Gb0Z6OGT5HAQMCJ2fQCJGNqYEk8eU2wF9ZYzvn6Z1rDg2DFZxm41UQzmO+QbcHDhLrlpfNxu
zrEvIZ5ySV85FAOnC1QK2Oyfbons5znFUzbl/STU0V+60bYJM2nPRaiOcBs+r9L8x+Oo3lICy3OX
rGlanmr26XMKrKesVkcOnLTdZDxKC4JmFMiPZw/jgjROYBzHh7Mgd6KNkHaPup6jhjlMSGVfm3Pt
3RxZjPYw6lTmns0iJ/VfQn5oQ/3OSahlSjDh3i6YI91Om4RmI5AgbWbmsvvcoZA3VCMNjCypWCOT
IwqPwjq4PkYSw+8AEUhszb/bjULTOWR2vNJ1WLMIGRBDzge1UzJv9uq3fha0AD1F0quFjIyNna/a
p+jT3EnCtqfxO1HdJSg8G6+hv9L/mD3tdWKud5qh6jsFNhemY1JXnff+Im64GQpnAT8ygRCR8TaI
0vWMRRqcoktMpFnHKcLgCR9sc5YJzs4M90yxBeJuqCmOTTNksyUj/rCEIdn/Qdm41eCgrCXw7i01
of7BAvyIind6Wuft4JhLWWzhYoBfxNTJsOFPAlI7Li9DwVI5pCAihw8jBFYhcDF2JNx/35H7MVmn
FUkAVv3sLFjSX0ZufU08i3lM3zVoX6gio/zIrPdAz9wATz3RKF04y+sz5ytDwXcRx8Q1v+aIJV7Z
pLj6/oiPcKtOsiMS5ROsES2Q66gzGweUw/etLoS1ftcKMEoFzEYErq5Gw4T2lBK8P2RJtDaluNH+
Z81pK432VJr51bYK/Sw3Th/ugY3wHhFMkCa+QlV3hW2OtJplrfUxNESCwMcwSyF9pvyyYPYKBmbf
Pa0PNpjKADZ0eZUMGhh9Y+avP3V60Ga5OzIx/HW+ZBM74Rzop57C4X+NxwXCtSKN9KF7hIyzyXeU
aQKBBs4rNp++W9GOM052ViZyUBDxBF0A3QmVpJZ3h4zZTU9hmD7BmHKE3RVDdCh8rd7harMgjbPq
g/TWm25D9YJ8PteAS34Eai+JBb7L5SdajIjsJctWJA6ilo7pkl75qpNmXb1EJ0Ne2b8BqflQGgLT
FP4oSjw+vo2kJ2ljZ1alfPPNPaCJpNKLZebJR5Qum0jl7MQuhzsOiouH8rd5UI0JM3QYIRRLOG7X
WtP4rR4DRVfzekxT0B8B4QcVYZEHiZ5xBWi/a8EXZiC+/23eCIO/vAVciFWQxJPjyf66z6ewSWgj
gs53JXhZopVaiNFDPOab8MCKM8yl64JYnDmV33VWCj5AS9rYVjnjKtWSlOth6aEqQonDsFRtsz6C
Ou0gkW7z/Zpf9u92opLRwbbUKwk0SivhqRE402bIh5VDA99El30bV1AeEIIPTt8Lzj8gh/t0C00O
+jo+MCYy4DzXtLD9ekYVGRHGSbMloAs2BEfBisZunuX4R3w34EOWbn7pCkGbIToL7SYN+L/jSwLy
NiriWcabuQmCuCJfh5xmZc2rY6lBfBXrjZd5x3L2bgBwRNbYGewMrkFsNqVrfCBiW6Z+aGIcFX+K
5Zl+N/rxx1J7mD3cb46kBzb7Pj+jJRd0eszJKk29at2O9lhCkwCUdKWzyy/XS27kD54gjR4UFERp
ZBnANreSeiHdptFo7JQIBt4pxAg/m2DVC7HwCvG8ok7Mu0pVJQ5umvdpSgLL3DMQ3ZcBab9Y8LL/
IXM966PwQq+f4iVNp3PSy0f2NxLL0eBoP9FiQic6BoS2zrsqPLmwExw0SB2VmMtZBnd9cQyYSGPa
Re5RvMq3kTGpwY0qiP5+YNuX+PU4Gt6VgjcC5OiWBTDiuPfW95r9iLgQA3dIIs4zGPC+63ber4g6
BhxRk4C0Zwe1sCg/jZNLCBNaGFucUeZ/tRMEXDx+VZJ2/iqEScCS5jJ57LxU4JQZgvXGNZ/WfyVj
kgshO4ho7PIDb3y+O6caVCIiuz2eaE63c6/2bt6N9p42HYuOqhCdvxjPEijgdh3DWg0NgpLDncnY
+Dl6p6WW7Q0b1O3qq+q4HEEKfFtwWkCexb4yQS/A3Fe9a+QZPH3FMnNhWzuQIOuRhjBAIpkzKvvA
1lB5MEE/8h93DBKoI2JfQXDm89QZlIfUrS58YrfMwVqFVinZYd5dAfKZZkXyYyoUf3EFMU+JhD1Q
eJdJeE3VSRQoZCKxD7Od66TDiFIivwsBduScz6BCpuI+4ifJb+xpLSVtTVw3Vj4u/I3CJQ0LFKiC
akkJi3JJMkjTxP+SSYhyGe8UHgu/eEQOw6PEtilrdVbsA5j8pzT+xMxtEeL2JJ55fW7gMX4rygIa
WhBM0FMWxfWNMiZVuxy7Vo9IPMgU7MYAA2PhUa8Sw1B9Vm6THDk1Z0n5tLBLW32TZcMFqr+tE92M
y7tV04jQE97KDEKV8ErF1UfKCrHn+mBjjy+GlTzDu3IrlVluaDpm+gNvROOeHqmlJdlDXVqTHBaB
hbVOexz+d6YJ6WroONhv38z/HshARAiYZjSCeIM8qOrLm4dJ6uKv9KvVV2ydtzg+x2iOAQqF3ivS
MeacHeI5RqKn5LZFbVs2kvUcDRr9Vnj+nbi3Nd4NDfgs+QcjOoctk2UwXokh0kRY56786NgkB137
/SStWmWZRKUrrhxutk+KyTEb0Jlfc1BnFnQEMI4ErjAbqQXgCuu+CwSeJr/Rt+zYzoO2gMRmyGgU
qv5uoIYZg5rKLpKESzGq3N1NLY/MhpUMqWulyZfl3g57Vjn2dCnVtsWZWECeoxmaUnUy2yWAEIX9
9LaaR/yuZqrR2qJ0O51iBUe7td98dvREFfjrQE8JJ6IHFfgj9zWbVqaTqZoVboflKghoazdDv976
8n5mT5G5Ze71fY1r52A5y8RbLYfWMIg+OVHtGhIDjnjICLjQxRIU01yo2BPS0zDb/Q7GIz4pIKoZ
AIYmYBxKTNUjwU1/PGLH7PlAdanj/qZRpAfswv0LgalEIrfMulIrkjdc1PvAp4HRpKt5xQxkVkno
DOqYF9ULx/Gbgb4gOvfxEQDXahFhjSO1v5AThHVGS2hmQgFgAsYA+SpphzLfthX1t1KvjmULhsS2
D5FK+YsUnZTcEuPnA3W2k5UnCv6hxfOP7o4kWgUSmHFbU4FU1Lox8jCoKjZ2d3RtmyX+WtvJcYeN
r3EbgQqH8Pgi94/n1TN/oPuPmP+7vpkQ7qvceCVKyMwK69UFXBc2EMd9tZA97sL+YkTMNq/yePg1
Q+PVGgWYnArjZ8QAZr4zHsIBXnZhI7ojjGv4rf1UBBpyxC7HMk70toUIM+BfxRmhLnVMZuz7+yUc
C3RolHezVTAoOajwWBg74t3WoVSvV3CI4MAVAT/pR+25hw3o+Dos5WTrPEL2iGR2fczvEDZECwMY
le5fZfkbssbU8ft7anpqhppEI1ymJjPkk0A/cGEoKwif8qTQuzDwkIudCAJaTHMMPw2aGmu4n6Oo
UjnB1+MTkdUrb3qsDLoa3cdvbAOoMFnc3qWEIV8nFAOR1IB0CcGDKQUmHH4dC5oz09PS62OSMs6l
WxBPfvcnlMwR1QqzLyyY7Y1jqeI3zdyls3+/KzAC6wtwo/Yp4lQzMXcNDrMWD2/rPELcI1qE4A7L
4v51EafeNIG6Ltc7ERyQVlBXCVkMdfQyNlCnFUrwVZR49DB4BkoJsGF6+jRYJfqAaG/HM0AGFZei
poTFoSgSl2eq3r2hpBPCC1pGwyU5XBp8sLkOjugNARAxD0uZQStmYSwwxpfrtdkwFqI3ps2km61T
Qtpjq0HxEi78CIrHO2UXqnKLu5C1Wxxtob+WinCHf2UZbywpSEftWVytXuqgvfbgy/ehpXosBHMa
6vczUpF7OVyhRP1plDuBpktL1xqASVmeeJajC034yIBQucS6LF/PJz6gVJeJDKISuvQREgysptI8
tP+/QQ79xc3eNL2XlZnS2QZ8HG4ayAE8YfC4XoBc9Q0oUhlxUnYnx5FcWox5P3nsYxUi+TN6YeGy
WLujNBMRTwDbrN0kNb8fG/MaSHRhvD1bU7/zRZ50ZaC5b8a3CoXsz8CtCxEh+WBXPaKCF1UUaa4W
s1WUPI0Qz56RX+Dgejjz+u/S8VAzWSpumOGWecpQKIOeVXLDkC5sY6tvCX0jzKK3/aH31sz41aJj
EpwTCZmUCDqcZF6ECH+1a3BQmTKyHyRPHhQHLvd/0QqzW6oP1N41vscTx7E4fQNXUphUHPZFrmK8
1PpOVn56psxRQXCiEYdnM18v5eTO+Mw4J3n1BSMp1s/se2+bnjz9Kj/3djqDszpySQ/iZuRW2bsR
OZylPB8ipHmxXoOiYC0lKRg1NlV5cozweLBcSW2in4p+Jm8fL2yANXnBmWPfgkg1Clig+aa24DVy
rEdFFhCBRVBVaF3B6VYiS7blce4LG+c2Jbw/jVkuLU8xR1KSfAew94lNtYc9VMa8C7cRW1yfjUL7
GCLOik5+sK8wlwmYzvkncRaLSZZpPM7jzlAwAUoMHGdpEuTA7mqEDkVfQq+/5PzMIX9S+ugCLArs
UpDjp+1L4hnr1q/dVmaJKKQw35OgT5VWR8W9XhzK9GfP7Pu6CvCO+2DALVBHbG2g5iBKVkl0JdnC
LeCR0tG5cmLshCRvNB0tJ/J69hEu0Xf14RS6ZCkodA0kk+m+72qYYu9FNWsjOxYNcpc9xue0dl5l
d1/HVkI2JwXLintTlvR6+7IBclVPuIJdb4D2c1pnRoDKQ4n1oSYiZv6w7m/8b+CrRtp9uqP+yQ9E
8jg8pGXA2mgLfn1Kt5U9bQtXZu5gpTV8JANGrh5a/QHYave4IPUTgJ8Fv6UrXbJk7ZmhjgxFk2tR
AsdfP2R6PSt6dtiJjJQssKqNkgMTmNNXhTQ5iwDZ7GWg2c/i4VOBp1i1Ik/ixYLI/X+Dk+eC2yIX
tZ99GxN38S8S5sHYMNPX+2xlzdBDGy8L68zUGwO+QmbUfAuiXwpRNx4O8I+i+mLes7kytAGg2rL9
dkMkJfwUDV11yOoh/ERaduUBhpjP+0/iKlHpWJy63jreoQRibd8FaDtfD1lFnUSJFPPOI7u89Snn
kddnaoxQ8ftFQZQlP9tI4jZp4LTlgG4CYYAEn1iJqf29xT/ZmMy1NvhC3vJIHDOr4U4Y5FEn4szh
OjJ6XJOxeZnLXALaXhnO29Vc6F4qBWbMM+H7hdcLRtmdUnEFLZeWjpHxojUhTaV0GdRtQVdszLtx
gICzRyUOqb7mnv9RXjHGQLEPVJlP1hvtlzJoE+B5avQLXNSBo+kNWKwoMyR3YlvL77YcoWV1wtI4
DHt/gwRnn3VVBs050tHSmzNVGi6tP7NhGxp1ukwOFu8+aH+zxg+TwY9plaRKdgFOqnMHG3z4qa3c
55voS7UDSplLP2VyWJ9Si7AVyJjrYgjEdHT2v+ZvbPjEgjV9aEAdzIJlM5WCEkif+M0VvmcHt/06
A244UphGybJDh7DDI7NkEnsfyLEu2MKo1KOc5XB+dSk5zzE5YY0UdIN76DYppCzO4CT8Od3nDCAa
/1nzQEgFsh/Mp7bpYaafx2d48VdNRwE1O2a7qX69K5pnDvAMhzVMs7SFOh6petVH44JqjpSprIy+
aZTQHF6h5DhQuuASw8J32yhKqtNFTyqpM0M+wM38NVzUf7czbo/H3mkJQj0y8vx9Pcq11W4LPyNl
ujIQFABunyge8s10kpPVB2X78SQa80JobwQQZ5J3+M8etjvGr/Q4j7vDV4x1dBn/GdYFfOU2Iizx
k8M06/K8IdpnWgm2lzWSsXsiQ+Qgs0I1B3+fLnmWwYL/nAXJIA6MS3Bmv+IFJk2ie6yWBC4mt4Qh
1Bo3M0dAP2su2/LXJjRWs0Ugi9hRZOzAmQAS5wos6dmAYXK6srAhxiwz2ymMONCxNNztZ+fWEimg
/Ku28Pm0O7SvXrPJWzh+huzMc+Vnb1JtljeWUQ5O1fPDYrrQavviHsKz+NAPWQgJANFg2Bpyd+I+
8JZ86jGfAsUKs5niawyPvrKbNItja8Ew+EAJcQpxeYkhZ0eugLhM3ddI26OiwQvnWRTczzejKEiN
dVJ2RPeoe3/p2E+pwKhHseTVUPoP85D4x8+kYutYkGpzFlDi9Yds1qpDNfAtd2FUn3Ot0bn3n92Z
uajWlws1VosZJ4rXjyq3G3D56YB1F3VNQKtI952xTanVIvxyy52JNelvBaANx8EoDFQhstp82OiI
W+6FcpkQbTMLtBWkAS/Fv48HjP+nsXoR727vpo2CYx9pdUNh9L7Qufzid+IS3k2AvNJi46Npxl9U
krk6pEGqGFQYAJbvprU3zZaW+zvlTiuEdsN4FL3ip/CJx6nW/iUpn3/B/beZuCv9bvjaytp4XLQK
vEAKCaNDCmGtXLT3zcEt+W9VXcYZogaUb1NGTmqXjCq4oncinu0PsYTAyzjC0mNNvnBg/6VL8K1f
P3l4Ij2ZKMmDNHofvDuOwy0e+ugQvz+D4AY5W4ujrUbRF0pCYwxlrHLPyJMy6WLDImAqcBWQNnah
5RhqA8+2O/bb6R2SjDsg6a9ewlMpAJMgQ5pt+1lBQPSuSwu6xE3TsVHHszv+MEksE8+wNWhQ5WI6
eFQIWZiQuk+xDhR09ec4uSTyAtu9j5GZ5JfkZ/M/MOIweC4UAUO4QYFFHKe75m28sbTEAb+zPLc2
Lqgi4+uCodo/kh1NTrlA1EEyQxePvWt1cyuiL620/xnyEXSfXusZhMWCFu0E65/NjC+fBk1dFL2o
wVBRYTJrD5rzeHkiv94XXFPGriu5BgRMnaKqEjg4Uqyhj/EVKaaNbJKugBv7BYHJdDlX8wvdW2E+
NhzrM10K23Y9wlz6GxxQEgDPBWB2+sWoI2hWzMV1GyJbuDu3Rd/Z4mMQrMs9dSXGTCY3lMF53qTG
Um8yh+4snD2zdbJJrsYKQkvEsivW02M7VFzIOSe/b3S+Df0YTJel0X2A6s2WZcxJ6xIMEhcYRpjR
FvQIT4XiLxlLOXUqq00fClZHAEAvF/k8W5qku3K4GDtaCqbqoc5DG93J0hJpRrYsHk160s8G1RSA
vyjc9orv88AZDpHYVlf5S0m+QWiWr077LEgkUvEyhKUCIG5HI/dQOJzHbipOKIk96OWu6eunB69h
ylYGwLuLjev5BAIPNUcGElBa4fdsovdI0tE/5Fqr0gcdbRfseoVurfDLGxfDXQz1w+IpFBU2LEwR
UdgCQd+8c2le3WSL4ucVbcpbRcKfhWBtxYnVXEDIjwZ6ucfitOJL9yprkf86JJ1iDGkivHBWKcFj
/nOXgTd3IPtfLIivNi1s7zRhgrJWVur/Mak+eVYSNdJpzj4xic4ZOuzcuPlDe+yOka+LwqH5YI5/
gBE0IDDgzkLhXjiSOBEmJwEwNawd0C0waakkBO9ipjUnp+vmpI5e3Ndsz20gAh0fRZHU+udLAOpV
HbYkwqBMBt8zEStYUgX+NpPFsIeK5Tgdo2MjcGGRw1+R1ZlBWEPYw1QHN+bslW8lrnQJJKHpsHpp
TmS7JuOh4Wiq2l5PJXLByqPG+AVrQeMSXWhlLBCXjUZ5G3+hFq2NlZ6Aq0fNMO4FrV1luu0KAhMx
oyK4vvx55i89zapKldW3AhHfzorWlHXDRRs/glzQgMyQZe0E2ATJ32UbX1VqJ68vZ8iVy++Y31A3
0cK6wfZlDjhq0pQKAbquQQnCDwTy9PBrCWA4h4pQfwjia1VuOK0tYK/b70JIO+551V2bE46It+OY
feCW1oEmbPQpnQgIinJqDXQpQUxTiRDtpijyc9WnRccA66lrbnitvTABAvKprrAyRfW6tZcQjYRd
V+GquUGqgypp0jZwGGgxAxEZ6WgN8+y70eLg7jOLqpTEU+QrOhSdPxLbVapO8ICj5tzSy8cxClid
vsVi333XWfizbNknSiDwhvJUYGhilCE3V5yMrCqvFQdKl75+UZYGCGu9YnI+4n8NgNXtZn4cyFzl
Oz5s+/5Cm3++cIUYhWrfR3EkdmOYumsHkq7xehtbEShDV+XkkEG8uuYaiMxWl8AvMgVKu1iV+h1V
0XY7ocUEwJR8Pj/yUp8eRayJJjdIXwPDaaoL2gBeQQxDlV9oDkFR/FdpbELuB93ey1NK4tciq+IZ
Af3RmIZ3yACh7nAANIxGef24pIS2cuKS3isAQIsp9SHxlbe1uHhW63sU5EEXTpHljERhTVpV4oHP
fBFimPQZpjo5yTnNRNZGg3rFe9g+1NHLkVh4XdlLqVDjMYZbCsWR9Ni+yxIWC0Gm24fKuEXi9K0M
cfifOmwzLMoZSuzC8RXlsW61SIi8V8pz6HhKefaYkcRO7bxsLClC1ODAbbzYWy4/qQhd6uav7StK
0qJIB4idnOdD57ONuLgcR3cYZyUCNr6BI0DqxId0oac99XHYuuckObotwGiGoopLlJLckO2y1ctT
talJh8eBp+2xDwqAlGm2F4r708SL6RdDq3spWwmwfo+ZZ4Ad8LiSmIdC0XUtx9Q+qxSKfly3ZrOx
4br+RHq9Afav4Q4gJ847ikYqcmxeCmdkcSp/nftofCPjrUnFImIWeVdR/r7uNnD3JfOvLVq3MVA6
yEEMwBzn4PKvhLDLunShN9FIEPEcjsiOcjGFmnl7zdrbLY4mOiWlqe19ybH5fpnYz51olMnmgMFd
2YMhL5BWZCuBzu2VjxfpDcYwEQNkMB6fEWakJOAw0vlvzTpLO+Xoc7U7XmX9043cVMCoOq1nz321
t8u78P81mzIZ9JaKWf/HV/anRKhtJbEtA+8dIIfC2wOYr/NiEkYrND+Ef9TEqlkItmocfdEnhiS5
XR7WyA6Fc6KlOS/pHQ8fnWbJqA8F8xOf9M27b/5QVtpVS0dsJu0dK0qC5m6AFBL/Lm7Q4Or6evPx
y2bhSoyoTtCJcOLO4NtZsMIkGj5MpYBI5m+8Nek1Y3poiW6mbdyArNyfTcFxfEkwQisnCkXt9Xz7
ijeFMkArmyxXE0lqgWcz4lfAVQFhjnKl6P/zzD4DGIRNG7qfbT11rOmWeNcLoZQBvO5oyTmE/Any
ViB1ZX1AYi7oHynU13eW9YTTr88j+WD+9T3AucPmT+5D69ryVk9Flk+w5d/+HRhv998bnkGXrQxr
7M5v7fNdtt7dMAz14+Iu/jp8/NU4Db5aGK/JoshAE7vOpktRPB0JRQozmw/R8ZgZH9O3O3BErfFu
jFFKDwdJCpoEUc4d+wvyoN6V8vomZoCMMp4gBPXjab+Uktusr+k/mhcf51d4nDk6LR4pFH7qRaDr
riKiRHWlyux/y9E3PKu3szxU260HqzJ3hQicvBNuvNkdI2bBkKtdRWUfXa2fGDhG1P+5wm3u+0N2
5Uagdao575N7mikM8DyaveRwGkq1GAgMdEuD+43SBvHKovM/5A0wKVc0E3jMIg66be+mSSygIxzX
7VQSWPbWrBbK9p9M7OftQzmLdneSZ6E2Ws3xi2PymgV0jFD9pp6LdDGnyTqIRQEfFu/tE2CAaot3
gmaE8t9xYWbVkiEYAhh6CUP83cm7Lz22O86xTQ0s0JTKNAev6ZBpnFdS07q+VVoS84Vk4dU0xvjQ
rQUPwd9/ZX7ZEga2/c1j8/vyjgsfC8z3UoPenVo4aVSue4jWkKOp0RWLVx4CxepsKFPgNFY2w2Hy
KvrPTy7FEnnkjbhWdWx7x92yzTzAMxVfRYuYJuiM72uqEAY9MbMI5LmyOF+5s+JPe6q5CGe0jYrF
dbKY1RPFHiyRCKv9VvgGoqaoKwjMOgfFcFCuZIHlkDOa4lb7h9DLHG00/YiomcSKnKI9jzVCI89t
aQgc+zxYl1jFxVMelBP/mG8NsHPAH8jJ2VmJnM4FqML+dmpfXDOCvpH18sGczlC7S5Kei4ooYd/c
3guzxJF/wnLAkapctPtdWxLN39HofvpwxJCb4cJ1+eQ6WnvjjZE6+B9etGSRROCfe1M3KemLKcat
oKkO7/wMAjiWreHbBfVBq2H/bpnSjJBAJ3REAeVRAYQBiKinZtWGqIz1A5JuXmHqb02DJE5x2zXf
kSrc1wm09yz6R9LvARcPcxjbjaVYnHjVsxqWSrO8K9IWuzRFaNWktbQJVSt/rIi5tQekZOs17WuP
yOJsiaP3tkSzEuabO+m+cVsBLecq9G5XxEvjxn+8pQ2TgT6+Z9dmrXuaYZUNjYJNPVd/InPbkLzx
m4HbTyJUnJp0PibJA5Xo2Aru32ku1YBNXqPfZpGCCBdqHFopidKvIYfeUzUEMGtcEVN2brp5D2/+
g8gK7O8wtudKp7pU2MWXZ16lPDSX34RpTNPOtPLELqqLLaLpWgz98RYhuh11yLHVTfwI46ic+eT6
bc80WWsiOhXh5hBYlxPeJVU2yfMqlpSXYY/ctfi9tyqqthrcg8Fmatsi4W9ybu5ehqLeqwZKulqM
wuA/6g82NKe0IxxWxSpd/bfqe/eQIbH1qrPw0uRs0TmKrNftUfpfJpf4EcgoDJGuCRD21eSB1WmQ
oOiCBmvq41qUvtCdTPARxJRknHzvVvkOUbUXr+aLDWFKOioVo4im65Pf5AOo7GrDbBMlqk9UCQX7
4oXaUcZikNwXaPpZ1rXQ6p3vbwInw808ECdaD8aDPkIXGFEyrn1GtWXZpVQDp71CxNBnRrrtfnKG
NeZO0FbzAyUqx7EK3zy7Et0x8/gt3+ctd4ELZV8xpXduKd80co+T0XctLLTuKfSeqmrBMl6IB0x0
cgJe7w9/mhFnSk0nP9zcU3L86BJrM5/kzVg+MLkYQylQCuDYQxFgJSddB6J6+ISnvX1ksT5PY3IU
2vAwMidj3wcevxA50LXuoHp/WxdIc3RUaFewSvgNmV9EsKUtAiubovLc76tJYKLuoc3tdLDPcTMs
q1ZgO+VvmdmI/4OGLAZSxaFbSPSIPmMZbWVfXOSJujW4oxdpdaFleOiG2wtjChf7zgAfLlRTi/gE
qlPB0lIfZBp75hE8CRD0T+x21d2iEcWQeGmnnPX98yOFTIo8mGOHvc4eg8H0sc/5BCh5zw7vFgAl
7/ucLGKRGcXYWzBJBesRhyaNehg41uzlJm3NFLjD7UzjPay0RMSnCJ3csbG7dSxWXVr24GBPd8cI
XFNzPasEh9SEoorMbm8wVcv+Jk4VW9JiS1nK0j1ISWcRX7CONv2FASNylMj7iT68JUmRFDOLV7Tk
AaCFlDXHy40s22Jl24Ttukbh+lAlfnyZNVvzb087c1fH7fpextmxXIz5aIKTwvX2noVGJPrpUVL9
klTizYVB3v2dE6bHI+FPpyDiCLNlZAe3WcGiqnlswlVushgZEzp2hNX+1pl1cKKtN7JYYBvsJQoq
jzc9qdd3T3CRUHr846vSDWepF9WmKGVxTLWXFCxEzSXgp2kDqcP1dUZ/Dpz7FeZlZY8ll83o3cp6
cGvClW0YXy2SnWULaQYSZfgeJ8uXxZLhs7/HR3NAdb/gn2TJBUTTLkLb2FAD/RvERApDZ2Q8SBIn
kT9U1bOg5dOjUGN7bCHJkfBtzzFVi8LS5ANTdtYOp3OSMZx3WpdZDH9h41w/Y+2nsVACBlggYOZX
1UyfutMocqHekGcNU0wMSRYWl7oTfVAt0VqbTMH6KJOdXhRSkA3ysmJWg3zG3g7ah3aaQwuDYhJL
50yl8FE0J7k2B8Er8soTW6Rg/Tzh6mw3tU5K5+5JRLQzxYHUr0oodSdpuAtDpLjc5vOK8nNGyIsF
0oCr5rN3GIeKZRmUB7JTXrQMt98lmVh6UN9O6l6oVdiA4zo56aY4T6/TzCRVil/84+JRK+x282SQ
sWy5ugmoX3QXcITe7Cgsi0EAYoZNr+hddam+I8xaHTuel2Rb73bOwLnV/kXlZplyXXQ8jcdFRQLV
EJ/thxWyvyg/7+fMvD/U3mtVouNSIe3VU68I1NZcbf9WOw9f7MpTRl1Y+MrV3+0UAjJtH3HpNTTf
l+UMBHfBJ6s45Afh+lJR/vAKwMhD5SLXLjeJ+AVm7I8vLP2HuO2qihAiO/dakyRpF0ruvCrPUZPx
Dx2sKu268/FgSf1ifznurl1XY/2mANSmFCyoXp+zd2tWABCdkaLP5jfJOoekY4iLfB8gzpS1xzLj
p4qYMgRvIvyrjrfnQpgV5LMLBF9Bu+kDlM0csWIiE8O05/6+SHCnTWhFUHpXqCEmfF/KSAaQyDCj
pGF+lZMONimuUthGFYZz6fkyR6jKNJ9+PDF3C8FWUquhxz0keT0eI1CNRJN+YtUgXwz4m5YIHX3x
9WppRqjZsch1C4njQQp07ZnkIyhM6+D8XjNGgonqwdXPTOrkhk3C9mopNITi2X9ntpmHBtPuBl78
Q7NmiAMO5f6BKIVCXfGCaaCvGAe+LWmfInQldpEkb/8NIcqGegETncFdSfF3R/UoEvaww3eS9bR1
pRSkupBlYKeu+alrGvuPknlC0z5H3JFc0BW64SGizYYXamvfmihtXl0pvNzDqOEQeDG0yd7SVJHM
pokpadpXicxtlBL6hp2MvK7JlVcr6gPXs3EcHcMopI0crw4rRl/RryFLAy69JdiTAiAb7Ec5ZBoN
lIIqbYa/JglG9YS7L/gmMjuLvIk2sL6qow+IIxRASGWF+5mjZWlf8peUtSXtpSEKKu7ifOacGulx
xUeixFtZdkV2XYvMHtqL3bP3TRfo8GSFluRXpMvWk8AIZVqzp5p0wxDNhiHnbSqc3p6gU5oducP1
So3THSNRKWPdmSI2zYsO6HAxK6IrNPn3OylBgyaE9UCCXtu1UQ1YHgnABAcJ9x6gEQ8Wb0p4+yYz
j7kg9sDpF4KWiWuHoHo587qAP9hGy0XYA/r/ucsY4ugPZH3SCbtykkPcIhzhqLhIAPeVagogqBke
RMMjgM9rGGHaKBSvBBgsFEbmDGgHSGVBp3KkT2OGUVgTXjaSz6tXvGpGW5HwbcnzUn+80RVaXxni
jYihcCBirKTXRuVW4NG6fpF0DcExsiXpePSrgUDnGAZ00E1hQcpoRhIP760yChIqNbsOA5cPX+Ar
fHE+cSI2BqXY27Jo7oRX/LSbN068saa63WkNZpfA7vE+kroARS44Ipw7bpYyZu5pVoxdMj6uah0O
odDeeYBU+dI1Kb/gKPx3wP3e7uUP0ATUI1lWfj2X9eWYCsu3RW77a9MWAPv+9ii5naLh4w3z7AKP
3hABAcWVh/+CX2i3Z6dFbBFAToZK5LZNRJi6oqrIaU7wPquS9Guz99MLRqfW6zDuQ01Uu2hH5WML
4Vwka2Rs9dKGZokMQtE5lBA2wD/jZKx0emA9FISHQiU8ybDytL8A3Xp7KXqsjR5+k7NVbmSijSos
ctFvdC8ATKoEbDO1gq+fksPpesLAaOhIZPaz5cN3dIB9io7udNoWP7kNUar+SqoPg+lD/2lPfVou
xDJ+r3LZgu+WlxTZ5jIILPILwv6Q1+cWHzVdJzzuKQc0ZaL4H8MBNuZQaZP9xKDBitaMeeEwAAGD
wuerJ6fe3n7ahN8iFwdg2c38MrzIFvnH9xDXz/UPxaPPLFG7dfs7VcihRHFjKrQAntf9AjoE0D/c
YANlvJNpKdiGyoyML0gxehK1CbnmpenPFtKc9EtB62Wl5ffS5JikrAVCUtpsY/s+e/jGfK7AnvXL
y7TqNpX8SBVKnBuxGD1mACJa3yW8rbJ1Ek6Mia0w40gRBDghNt68Fzcw/d50Gq7zrTz0I0XhzI+v
faH1EEY3EvvyOFJZ5HjExiWg6v37iRt8qINM0VGTo3Vt1DBXCBVr5D0iohkpI7yf2lj7AfovmSXs
TdtXhy5jGw7xScEGLoqtdlRccpKdr3zfaP7Fz4iSw3MRahGTyUQmAhUOTXiSRpFeQUDk2Zl0Pd6G
O1pQCkDqsZ/HPB3QE4zfcOV0kmIHZo1p/DC1EbtAXfBsia60RRpZP4GnlqJ6Z7O+aYA9czoJymav
IYe9HhJWajCpI8+uE8EFGx3wbQsIs9yL8RuIWOuQX4htSMI5zkr9Jt++1cyJxA6r0KFmOy25k3Zi
28DS9CUwyFtRjNXucBp8PpkhQZdHS3rlmFiKTe68rbJW2wlm5wzncu31CwCli2k1IONODNKwnfNS
aZl+rqe57+l5NpmFN+Sv/ZrgZwCzCMOUU/VWLT3gCpkWx7NkgmHEdmJs8UYAu8pC1ibeZR6in1r0
Vo+g5qS7fGGvoeWh/ZXGHprnCT1uf7i9za9ieMb8hBehB4y32DYEU/acXyGvEydN32SoaNh+uRBk
Z9JBdIKcQtTQwiXkVQRe5A392CKvPkIGVrGth5MU8bLxpgEac5/SyEfO8bilDRw0s4BAmnECafsQ
u6jEfiy2vWh+91vndWHg/0DbeYFElU2tDwoJTz9wqrfQ68vi66s3atRfcMB+AXCLzO+JOHy3N51K
dm6wmtMCOZbijDZnMdaR8sEctJpIbu2SoPbycKSrx9BiMmMBgQbsNg+SiSfrQSBviBneMEU4ETtu
D1VuSCLMcEZbLBdpAvGTG74RVeY9RDLH+e4etXF2rakJQjqQYwf3F1TX8Ardbwqd0voJpY7fHpfS
Ah85QPCz4noc5A59Wt3+xFJ6xW5GiO8f9Kq72Notjx5nHxReHybznhG53hNqZpuGf473TBkwvjzh
HlMwrYPRXFs0GIAraXcNcuCnvm8wS/f2uD3DMSe0uERS2gK3U9m2iKwbTDo+W7MgLNfVdNXFrwsl
FIaTKOysDmfdgjcmQe/Fo43nVAc5whuJWzRvKeMyoK+Sx2wAt62y5KKqM2wQFtDYxL2cRJq9ycdH
rHt/uf4rdE7+g2pe5CGhdlLdVR9E+l6jY2gTndw/KHe9q7KczPxF264x1JsMHicFDqlo+7fVvt6N
U4iFYgaGWhIiuHM0qdIpsXLCB2Zz9njwUES3qXbS2BwBCpUyfYhPKGW1RtGnRRMKXRZDut/ZVSJ+
SMzdfKscbhs02Hh81a7u+0lH7ez7pN689wwCWE+Ot/HAcUnO2KM2jQrPYw8op2OaeMQuNeA4cU6u
Ecg6GNV6KOIIJnVUAXRalw8CjFD2gFfQiV3Fzy/9mX86UfpmfYhy0WLhIwPEi4/9yGMlNBRen6sm
4+y42QNeoyNlwY0Obyxb5CxwQBK4W/5J7cAuR8tGjss25c7cGnhD/+8Is9SI/MPrV+pzEXqj53eR
lZhqRGj0qHFlW5rOFzJly2Ix9a4Msga5cftOgiuseUGcbpkH9Ci5PyvNP8fY57Pe79ACLNZwh+UE
+EvyLfD3pA+26gt/V9qTRcGZkTfw4aEn5/ief4IdRZc4P0/zA/bYgOKvBj/YUP9QDPOAsiinAyqE
JyW1JG68GT0GCc+QTs3+L+XZwMhTJVihIsStHnlokc4xBMYWotTqiuqMq0n8jwIHuNrk0GcESn98
UtOPyKcqm+BMKqfEBXVN8HMTnpoc5qQpLT2KsrNHNkS4rvYqVRALesjm1gfRZB99MP+RiLS/lH11
tf9iHNBjPZbdLNXK7skc2WG7/cZ3Oy7BGdsutBXluqqzY1LuZfAV8FSODuAhQhIjqyoRcd/TEoaP
c8ote1MiQrj72baQjTrRo9kyZYUMxxeORT9CD7R/N3p/AvUuyOaO8QhToREdKwhYkxLYhtTQr344
vtrM9l49/+yYiWA8H2KIbFhT1R2BziqHj+5JI4Zc02mBeiOWQm/X+zUlHntmRLrtY0GFrj277uSU
/Vvnk9jn5N7LWRuJh6G2NurdWPIXH2V9imxZKdfnjOHWS+8zCVtjG8u6M70sou0lS9gMQREdOLIE
q3mISXGEmFh6bVhWF7cWAUzGJOey7bezcoZVVUBGE3rMMSqT4ITpnp+sIEFSGOuWqj9K8tB6LwSC
gZPw9h1QbubAQQrOFEekS3LjNbjYFApRu0gNT9Kc2kCR+PLuRRNXAJG7uyA5ij+EM+4RRHhxgMee
Bgg6/bF4cLkxrbfvHqfUHGwE0IZlkG927wses5U8Y8aMVZLSe/qRks3yJ0nmbODInJzMo8TKscy3
A1cfeN871YCGiTbXRl1LYiE0rIYwcG9+Uk6jHuWc+Pw8519tZMrzoXOLVqdtVXXFcNLTogLQEYi7
SpycYU8DFHF668ZRSAADjLoBDzng9ZyCy3vFzLj9JfKyfhjJzC5VvP372I6ktF3VTsbG4qd4UZj7
0jynZOLW9Gs77rDWrECFLeR5WBYC7uWxfw6bqoxjRaQKVoUKlxnl9BLCHi0G8pFkhi3SrPUWp7uo
E83I5nm9bkQxToJv5gIL+bYXF+TVM7c3Kva8ZEjvYipv1Zc1q2dL8KsQA5n7hc0zZwKof1pnCTV2
KrW7rLFV8+fX9u00h7iO+rr1VkRZRkocOlb3/S8KqWSRdyIAOy0SM8Uoo9KPmkab5dJkKH12oRG8
ovohrKm5BVciNXOekt1YZec5yEik+cBUIaR3lxLXtMCfJEkW8GUQ04oYgHIL26WztnCHBBn/N7zX
ncRkKNUg9vN34j3vBFNa7X7r4fsLSMwNITNVBAPlDzBSNGJzfoLPGBlL4EMe7KZkeKqSn6Vn87wu
/15RmcxRwnY3nQ6paS7KEU0O8AjJGgfON5mtJDC1UWqDKQVvMd2RSwt3agkeevmVjAFsn0LQ5+fs
EWN26ua4xnJkmHihpTD8O9iXtR1608nFeXPLWU3j8JScrnwRr5vSY+JwzfeI4W6G2V0KBheoT3yn
gVu+jXqGiF4xRjrCawtWhIpSqMfyRB5e4iKt7mwci/K+bi88VrqPBJ+hQi+2iVg2IMVWEXGZkzqG
V8yyg2bKO4Xt8u1AbhrdfY4a79yCNzal5+luwMP1EpiEEm6vRzJkrYh0QZIoQ0b5/1WR6O29DiHu
JSug0+XIlKLiEousSa7QauAhtrPBtKgeMf9/PQxcDaFzcmxtvKMY3SDNowtHGWAhev7COMT2Lge5
9nwBHi6KYUwMkYCax4uaGSDRCeVkWkDt2nze09KBnpOB2zYFwyJpaUtGmEnJlGOrd3UkguJOd5Xp
mNmur1qFs5FpbqKj9FKr3GXpz71ltNigh0OTTKoM7lQLTvzoW190sju+eEH2KQitWxGRKB7y5wrb
SpmT0bcpSjMMrGpmNurt6D7sdtGhFPDVsKZXEnv+j6Ha52kGnIw40acAX2kb/vFC+acMLn95pAJC
VHH19jt1Gx/Z0O3sAlfrWenkuYQZcWSf++hchZznUFlT4gVbwnL+Qwm9DjIqrU1ukrDIL0SK6RVM
aiHpKBAlgA9wEYuTulUMcPIJj75P0rdhljvdlaQyHF8gHFlvEr7SsmvD+P73dgXFHjrUAF+pZYj+
xZYrUi3WigGaV+gHzV/zJMgGVSPkIGIexZ9ZBaxPBQ4tGiSXpvfKCP9WTlhOGAM13SObh0b4sujN
/FB5XNQGnNAEhqEZxZ31zHsPtWmPKbVKIVbd15rfhHgGrXLeZHTUgRGVUrDE/OVpS8h1384lYZi5
1hiqtzMnMqMvjbcf/MwvrxKp0Dw/YTtUGZ94Cax2E83jKnvOsDxkpuM8leqk639NWLP3R2YziHIU
c0qtYoXxiSFttGR8Xj4fW6mvgMUahWKt4Bd/ZxKVCnd2J2CWK9RIP4muoLiiRsz8ArSYbDBqsPfA
PFKN3DDXTnosf3FZuBE/zncWe6uDAIMftIrVx6VhOe+isdIBIvtfVC6wt/tvAj508afdnYgM1ZgI
GvTSroo2RwUkVs7qfV8NRy3B8BMToqJtT83V4chHZn+IuG8HDEJWtu9O5n38t8k94TM+9hPRqpa8
fiG8L5AC5/j+sziXbxPNhf8q1H6w8QhL2ri8ntLgHl64nHqz1lSQRbqsyW8FGXUPUuEKWzMnhZLk
O3QOcxDEwaxWMzf9yfIwv80yUguftrZg+++bx38J4REiyepeSzYQG4lXFKVWhxzj6C+sZJp+p7vO
g0Bm3RJRBwmAmcP2bYUtDIG3ICspCdQjEWWehVzMbL+MM/lT+SospBsia/klDNiq2cwXaqqrDVYa
fRZM+qvupyXEPtI6aIEl7qOKRSpG5EsaPQHomUSoTC0RasL4fhzqKhRksrwiSMZv60cLebpjyGJD
4QCWM5Cwtq2mJRN00OryzLnOQfAHvwxRpp3SmxmZpZ13ChNveA1i+PNlMrQX1ymkZmBh8BwliZi9
Krow8AOZzhVtxPzjQ0TmEa0Qqxe9ciUQYyx7/NCozrBEA+swEbFMrvr/+hcwB8ncPb/9d6PepXBo
9Q19iHTlK9w/rYAFL0NG4RJOa9/+R6aAOW8wHn7TvDsoa5gjWpWvR0WAr/NsxyZctbkR6yH0zrtr
nT+3eP7A8XGuRHq02qvH9e7rTgfz+2pEzKS3rvYa+bwLql1s//NB6QyPT/PUhwmx4dgaoAW3z7ro
4JMIHd+tblBQd25lK/X+AeHmMv0+cdUzOIbcgq5LXSpuqtXJcapjHvIyOWv0Nmi/yY22kzjjOxUB
6G80N58AArY53cu8qvpOyXQ5pbya5hoNIyLhnE/IjJRdd23fCJB/MN66thLYBw7C0MkwsrgPbczE
s8KY1pW9k5sZxQpmDebpnXNiqdX99d/vUS7Dd+TwFHCxNeaDDVDWYn2eOQN+Wv7FRzRCluqm3+Of
ddHkHN3GrxXiJWu/m/6iYtabxEsn50izLTszAsjAiOFfmSapZ2GIISthpzlI+6dkYwLAKXY1Yz6x
Qcrdj3c+sZegbN2p+xkdMUV+bq2CuyqyvfjMVKR+yTS4dMH/YKtlLVdjpEjPUxGUQcNhNlHf+i1C
v9b+QvgTdqspg0m5c8iGxxpM9dpX7/NtQ2XOrbrVTH3tdI03aeM5bh68JsIYlO9alQxxdOFaxXAm
Ye2xPELXmXAbdDX4Qa0RRNQPgwvb/uK5zPCyJPpd9muTDvNyR7l60EwUKexBovNq3aueS7sM3b9E
JZxrrnpqLKv3TnP0UUkt2FlT2gzWtYZcoLCC54qNIMpOc8RAe5daJVrHQVSSbdb2Cu7GaJe4/G6M
UFC+lXjBP9An25riSLKMGqW+g+Ze6HzgM8IcaI4JJXGvSxBmWHYvnVDIoeReJ4UHEXiMb5fblmjA
rwWNcXGBFmVHj6Xj8PFFaUqpYJ5RS1iqbX133lz+RgmGSm8nxsn8YQf2nrS3UMeqUEZClbjiwqTf
NM719eXlME9cUTpZ19tNAE/eZDbZzPBTqUTtrKD2Xb8wumvhFVAIPyHnj1U7XpG8FHbB7fTpwfkO
SQghjrnGm1ig1otypQ5n9oyo7rpiG9oRO/N28RMGuVQiF1JYvwMizc82GobIZ3GyjcDKc0/SmNs/
+22vU6mS9UKf3pPzZRy6Hh72auJJP1sNsujvtLoe2o/82Qdzuj2AMR0k51sLb1ZrqgHAmdlr61SR
wcgUxTackuAzYKQPTSyYylmlBwS4DvQ9r8GlxaDlli2j3QI7cmQ+AtvFeiDEJDw4iZ9nP2/G89Vy
snAyIYevNuiQPS61PoX8Sbal5Dr64gmi7+4i1yqlymd1nma/GBoair8t/lc7cZ6aSBbU9k+VlXMC
sqTGbmexiFAC6BV/rsgfg/bxpC9FwzANNU6Aee76prRZnzy8uxLJQU6XUn/tp38f7lHkQ98EhFdV
VMDD2Gv063LZ6QhWdfZayIBHBQl89gSW0QuUsGFyL9vqFRtwUjHpKRrEYys+u4wGBD3gb3TiSLvy
WE3seapj1/Gro2C2V0ukQctkuR6KL+NDbyG604xpzJTBdrlJPc0XHw33vOSiSlCsI7akjpQaemjD
4TonD6p2ZwZdIoY9RPZzg5ABssP/10G8PKrxBHLaO3z29wPedT5J3hb72G3uD4O4ALws/mqUeSDk
lKaEEo4BKoLJufVXc+jn3OTl8869soG4R1cYO+g/9UnQ6g/lzWogRHeYRpU4KuUH17LS6RYV5RWf
ei2NC/0zEzAgRpRer+Ulv3HoDWHzjkMnaOWHDTUzkAJFRiYfP2jDPO20izzfAhVz7jVj4KAF/yt/
xwDFU8MBOK30MyedVGzU046QyQ9rDlxquuk1vuuwt0D7RRiSeUXP5HGAIKPakc16Nt1nPXBbdjGB
y65fE74MXntkxvLShGrLzlPmk+6g7w/sobT6XCDxxN7f806yM1Cd7kpksxd/STQUGs3BWgJrgOIj
dRWZgaDnlfAEPdZxp9Dfw4UJxlsvKcOBs3UYuHrLqAjoo6G3NZA6jMf76J6FNcKAJeMcWJ+oZQgB
W8k3xUWRT4ybNp8YLS/+bFNQacWcAslhJASSyw85pkzNyHZsdC5/mNpyLJd6BoYGv/H5Qa4ByRlt
UjojOqcVKE7NdY5mjxmXomi6N84IjQrZTX75YLER4sz1Drk43KVn1YpATnCTeyxcU7CQQ/PTUzcF
pOA/rxcYtQF8RhAdYhLe1jGl6SNl+4/Z0R28XH/Ns5Feb0YP6GVb+h2AIJWIBz2jfkg+tpC+acWh
ObIagBlUh8pAPY0vgce0+MJ5KsWMJFnVkqGyGqyvTKp/Uln1teu2UqHYqmGg4cSql6jKutq0Sgmr
7+chjz1uG81uKG+TiHwFuzuS0H3qEt2jj8SZVjg7gIDrjY8LV9efznliUNvSWOiFSNxmdmk7PYN0
khWfHDa8VGyP9AXVDgQNKfpwArkhZGkvSKA0T8xh6+Xrk0dLa5/x4beB4VLZb+tdcPgdnSq60Yqf
1b7u4DCdYKgonwlQAfO1Q0b7toA/zZ3aajrCtQGnbgHNX3ERR5KmmITIV5CyUpwG0W6ECRfmlFER
meVTx1GTqJ0HJQW9TyMoPeAy4ZsbaGclIFt/uuwdRdQIGhoVnggJTopxGSz+f/7nrvAlbt/TUAPC
nH0atzTs/ZvMeghOOmmbMXa26XuQwnESZnlavKMOrAmb9CGO+8g5ngDQyuqhULQaMg8lfCW4ooH0
q99G59iZkzD0HmQyMVl2Bd8JJBM74dRdL4BkIsfa3rO5aFbc/45cTMaHo0+N3QIXDDXQENxuDfFu
D4nXWriNkWRTBSVNuia/cokSbYooAffrm+RJMKoWIsYFXB5aVd3UW6rHeoQzzlRkB1PvCy/UyMYr
ZVk+4SkK4rGT2aQr4jCJDTWRY8efjmAtvg2YUdmTERBb0otl4UfImkqHkB8Z1oEEevZIGrLtP5QQ
JlqlrxMpyJVMICBEQIDsr5JEz5OCddLA1jWpM+d53K3vZzYi80+uNltEUuvfD7ZhCGiEtnDLnroy
xlwTTS/igspGREwHK0Er7ntRJJ2RUBV7QLfImSpMmDRvbhtLtyx+FOeKaDARt4kEf91kteHhnFGj
9HpmHuGoRtelJYNWBli/M7IO4bQaFL2D/woMprodbggwOhYTP51IjkW7tHhd+E8z2Un/A0n3OISy
ff8XBBvr87QHU1cbHXtyZNHE6EgKdk1DVwPXaKOhtdO7AyE8v5Wy4W73hDB1UHUWkwOwahsuXSdB
bB6ALDgEGbQCd2Q0mE6vU0rMXftwy9bhTjYnHabAYOkzNv9QWHIdR8UnpweF46EYpmwp/hks42BR
M7FUwn8Q8oUrXWuZgKc6XDI+o/m9+KjKAV34/UmukFB6WptNN71uAcysTotUaN7idxEwiXi8Togg
5+3mmA8ezd4ab9CRS5n2m6BzxzK2xquqWtz80trVZuUDf8K+ZgNyiwlLzHx7k6NaZiVU8+sYlx2m
l/02uU+wDiWUefBqpNuPzdXdOUGrW0XMHZOgIJQPfMUAC0gAM3e8IOQHC1wuhbwLAXwXLSu3f4yE
Ee72MmZMGfyKrKpQQsRqXrspxqmwzv0NtmfwoObiG1ZmSWUCGuL6n4Kqaiioa4fwCFTAZn+/V1kg
nd2htzDrOMyIouZ2zeuyauI1MinFXVZzja4qhdabo+Z625CPjGe1rGMez0TA6gY8ovpBf9ANT5uO
H2oTOLQQju9pFk051XbqmRxNzKA73XjItUtEJN3Gvq8nbipU3uc3YVF92qXeeFwWPyw1oLRkD00B
6pJwdhWMRHQxtaJ5zkag4SND1YMjmUtF+WVGpQkGtpRm2rQijyC7DD2gsvL25RkWTyotks8SS/QJ
ieJmqZArtvntGVR04r423SmbDqIMOGv4ORUSPRRZdhceVevZnxZ5o6nhQvDv+ypxeIDJ/DbfnOUR
iO43TuhM1Doe+wPsl2RUukIhGb5mCScjx8Eqzl6dFjDv71N9OfnU4m4u3S0znBFxKnqJTvTMwGCi
6/IFWdhvqNAmCVAAZyYKQ32jC8DNuDDo2IaLczsrTOEUlQgFJ+gTi+T90soJcJ76FdC930KNERv8
M36FeMDaYhJYYfy2hhdIp84Cw+zwQ3OGPPRjxfLxvVRtt+d4+uddIsJAlreEsTF5Y0q5kgSusqr9
X3vuYtBg0aUgPNJbNIjlZ/FEn/9z9mY3uUUOWJHHti75gAeDF1yBVLqZ6xs5gaYimSsDQO/PzWTA
GRlYdsH5zMzwDDRQLlXMy2/MI/mF6qckCnGQLkvPPwG6YQDRYeSBavMtOBO9hCsiwuZulXg6otkL
ZMaC88TLUXOnOlGqLR1n90sNXOd2Fif+9mHyXgJgbY45NueWS7skifI+vpB/Gtoh2eWhgsZgUq06
1rP8lfLIgt7lgUSLW3PELFjpSesmNlZOA67nDVi9s67QhLeBkmYl4aj+llIztHmegX1TI/Y1RqqN
Xj31YW13HeC+YdyhbfkJvjacX3E84eOOJo2k+BZM0OmcdyK8mURWlHxUe7w6OC2bgai3xAtsVqpO
85gte/Gh9KCHgG0lOu2cirY7ItKl+ZVAJgHmqAlG6sCs8/zKlf9pPASPJbgHKgEBCUjFU1VWvR+/
M8WYlUpWvUYYUmuGDukAVzBqXrM55KYoWe3pzQZO32KhJfOY23+5IqSxCLmuw4WafjzGVKN+2cBG
/k7WIk4thrG0H0PACnoIr27XLftxRofIx7T2KtE+AskVTf1+ng0Z3Eby0ETIK61ssyDIezUf62RS
zDKSkFSmW6WbAWtuGVl22fScNQpGL4VL3KSIM3IA6Go724xrMAAzj1BgLxz54VUKWpwQGV0i4bGP
Q0DK0Z2BgnmzVHIiaGvbKU2xZxNq9X0uNeUscZ4m9R0AyqZKNwhLLFIrIF5v7e0bYPq2luZFdLor
dXKc/t/5cFuony0T+NNKJj2g7DUIf+aAymJ/HiT51q9sxkEdJ13HTsahNTO2CE8Hmr7tpbu0q+wn
hlZ/g4yHhhUNACfCqrQve5LbEzTVH8WRD2SnZFmsXrRXpzT5v5ELum9Tei7r19N1Md2VKeglcI49
lNvoL+M3UbgTEPxbD4ssh8JyNPK4xYF171rPGgu4YKjjPuujEei7v2zUIqAObTudaoBatfEujKL/
WWSoWGAoRu7FGrXoD1xx29u0I3VSAbP+jxpbxu/yawfZKHtlfEbcoIrg/2Rtxq3edPn2iHH7DmSF
ZWRABMXpRZ48SubNA2vrTDRGXgxgOiMmePCzKnlKT+jNoQTVUVGVlP9bOHFgm7oVqxqMjO7rNT3H
24C2BKTMg6WYyH76OM8aZtjyNbiU0KsYTjTv+2hLyJncXdbwx+UrQAYA4CaQSAsX5mK1Ca8gNfsz
PP7a0vlqm1u4EIb7YOZ4pNpjtslz1DimHv4GTu4+vY6H0DsrwjM8k0Y+1RgTpwP31rmsBszOPOxK
fXVuXOzkvafTmWchj4GQ+qcueuGyeU64rUeLfig9sW9cTJt1jVaMwS6PlpwzA6Cvt/xUZ78CqXuH
F0RzwfUrgTq1j1SDL2pJDYWzFlGooMpyUp2Dbn3fQiL9oMU87EPqwUHe/kCJIF/dMC1JmZc4+KrB
cCY0NUwRyoAuYIOe8jqay84WWaCWo/5FM7bh/B7oZRGO3+b1l0o/dVtQgcc0HwYg5gNC9U4QvZNG
7tUUxiKAs9KYwOSzErUbL8WpKzQj1l46rwvoLSPnds/fF+vERX/EOU06Ev8se/+xP//jj7gEjkSJ
1Wo96uM9m6/4o3Kt5j5z4I3wiHSTZ7HNJ9iNNNpbYXyr4sCFgjDKCYMueK0nmTdW+A1sI5FDUu4O
CrRnA9EzyK++KreNKAFXLktzv3CmorgYI+SDtRB7dSg0ckevwZJeDWVaoDQqxC5YOks+6iUa+Bm1
OkUJyu2P6LHU/rfdjkSHQoaI8PnjZFoZzqKYVuLCDXI7XF2x+160qVmYQ7R48boy5BgFHg1k5QLr
rTNrLBxAaPvqDlPhiIIkxw1WxnJ2o2f52iSiNn5AR8Cu3tZgrzVIJ4CAnPMc3JS+RSqosjOWS6TF
i3mSaji5FbORpJ6JAWq7gSMXKoSY3uzJxZ5mz0jbBfCsXe2F4twdmT0VAZzHALlqj9sc6UAkDfSS
jFQpKzplXNau6odt4pZyX2xYpxwQvQvKNTGIYSSoX9gnn3T9uMTri0YrdpUbHIUX8P7GETrN03Cz
Jv7xd0wZR95sDGHeXPhtbYZlatC+DYvi7ogrv5EB1uksLolZE92WZvQprqaluL+RWVeHyjiUXGDf
QkTYG5DRw03v/dC5KhExeqL0SZRIjL8oAt30fUdbgURym/OJG4220X83pawN8j+5o72S1NWL/nfp
WHAaztT8Zs6B5/hmSd3i8ByRIkt4CTdv5/qpNCZSGWBr//cBjOjkvstQ0Jy5C89RyMpvvUC3Div/
2r5BpEEzqO6pze48izdUV8HI7KJv/1B+YXhg53ee12xmJYNUCCQccmSP20cdoc5PobOfBbFMePsQ
nG+1Z47wzsdBRyG/NPxXPuykvwnWAfgWxnjEjWN95kN3S8xE0Db2UezP+z5m+yxxLOObbuUWrVi/
pdXu4FNosWPy1vVLMwMBwJhgTwDLBf/+ec5PJV+Ifi1Xg7VYWBYa1k4kgqcE8aeomXUF9XMdhetX
o1rPgaZnGj0p2Kg5zH8nFMx8hm3dd9gIONfchal9eFPXRBN0AliPyGKwa5pIgc8ZLD6BmyQEZTZk
HG1NcQude9dhOUGUANiu+NC/mOCm3VlJz5UwczRw2joKpFQ9LxBDhgbkGYZwhSHPYl7vXRB8EA+c
lRO/W3Dx608LnO8GZ8/qyQ7cpFn8Z+NtKg0typBIo222GnhD0RcwxkczeLPzE/7kkKdcOB2ePIhN
DQ69vA2gkeRompMioWl0RXMgW0RynNymMFxT667jJdXbcF44tv4qwNaSE9VWYxipg6nesQ4V9MqV
SJW3yeWtBypCRPmsNr2zARbD5fqqzb1RHDHM1WhOXR/wYKll+iMXuw0AgOTaCUaZHGiNz6QemOw3
i4rnVR2zLeyWEsCc4rSrqiWGDiAI1rEzdieeb4lWxga0dFnl+/G8KkGHJFHoJ8l0zUN2t3LgLtlQ
uixlUBefx/rhYLLPtkfTVj6TUEDmMVDFTa+eMv/ZxwgaYwJrI2hlkPEy3VVFcYGypeqcZ/m7rrNS
L+uuyl53LIyl5jiY4YqTl06JPR8skSCMKIPOv1yfmHr70zkJtXPRs4n8ApdtFLBWGph6yBrkzBd4
OGLI5sE6G158MjBNvUMfjD6V6271aHEqukOLOvcX/Mhvava/0qm3DNV+Eft3s4v2AxT6gHIcGx7O
DiHWE/rA6emt2bAhIGoX6VnDrduRcmlR5TA+MrBeoHeNx8TEZrZK2czyAtPXFX8cDqe3BYDs8t4O
F7g6PjPGZdZFeTR7y5/BcwDE6pHioLrN4fG7xNV/HaTs4moUWcM2MZQrlr434uzNms9AALRmiCBP
nVzljBgBKcoKAkjmETTQwHsqcy7UyiytLKN3DdSRfUHygajAcy9edMwz4zQMBSs/9fcrt/FlyXQR
ABxSgN94zfdDEtZMWdtHM/ibL72HYlJYwWbpEl37zLUyf2iRh/hsL8w2e84bp3/w2XI4EvOfimcv
V4MrfTMPS8OruQZeoSHnYSjSO1N0F31PCnt1yE0sLKHAF0p9c1hWSI8kzoonzSYxDCryLqcb/RDA
kJ7ngO+YDlfO2UDuWsOBeaKxufjp7jv2osgfnXhGJIU6dLTkvm5P2/ob1arB0IZBN5J2R/7lqxdx
rIaSzOPO1hYT+CT+gMP+tYm/6RSLdJ2S/PEakIMIRdpsFw5JCK2Kb03zT1E1EuFLSc+ucEMBDk5T
p4CBnUFk1JBPi+4X4YNG3tvxz1fMOyLpRHnnVB1PYmPz7qjZ5qO20QneBY3SMzfeFHjgtMPlrmUu
S6n5FnaR7T0z7c+T57ipWIQhBKa6KQVYgugTsdSAXuvl4KSKf8vEaMuUck/nHi/EG9lwdnXXlsR8
Fv/Da3HWUS4agP9ZCcMuoeynjs5BTjJwp8gO9RrnH3+mRLDahi5e4hBXMEjdhh8Iv8ZCGiuw7khc
8qexgzE8rsfhD/0ZqkZvGo80VBDior+dgxEYnXcDW2V5XEGTykfYrtwWs9MaCT8JmEz/xskPtloK
AyzsvGc32tF3vKCIJN5a6845zIco5pO9sVp6N10AsjL+8IjsJejFfSA6Xk7wo/WHw1ItXHui4sVO
ZfF7FvQUYmVNWGFo+Ufvu5gBEYIupdN1HnFkRMX6gHDFw2TYYp4p1xh8ke8f1PQi737dpPegfA20
fm/hZqAiVouagwQerzf+tr81tkhe0tU16xEy2AIdxyK3UoTjEjO16LTvvgKnY7lVDv9XeZM0YsgD
EylerHDsLyrRATRY5t83TaWxdFMGuYNxRwDZlQPcTDc/5ccC98LbTPoD2V1R/F1DUV1/DjaCRND3
zhddVAeZrslhurRjPLHLRiikhOa1anF8VLaPcO0K/l7F03D1QvBP/sJezArgcSxDAzkfix+/aE5w
de56t0eXRev5lFZkwlYno80xRfJMHMM8jk+c2/jI4NmkMeu5nKPzkIghmBt3YYxuxvJhV9LQfncg
Slhmvws8Wbd7AOMr9QuqdBHDXlcOfFvfam7Mi6Ve8dMUYJndZbmaqOC+3ACXn8YzTOkuNR5WbDga
Nop03doxSzJ78YIxYGMciS7eqzwLf25m5yqkh8D+eA79QBxuR/US4XXbce29Kxvnw2Jq12UxdX1e
vr16ikLJKBYQ40k4vSdvfhaTavDnEqJzrqPXkRVlHYBVXWPG2tis9nqeEwy+DsqvN8XjRhnefoJ2
KPTrL5I57QJzra2JfGg9Hgo18veDY4TpuTvSan2xnRr4b0/luEtgXqmNzeP25IdGi/q0gPkW02FZ
0Jvputi0izNQIpFF6cIRbYUscC1JxtuSDiOcruB1oeJDQijlFfjMBSx3IQVPKIvk0JypJAqWXe23
Se49GxJe0mdqzILykvWsObUbYN2C/kNSI6RRVi8s4gffOYCbKKMid+pJtOn1h8vO4Zp2ErMKVZlo
hviJe0KfY7Olkr0oxqXLjGUkb4FzfZVQwH7xjP9q3+IMGfNpyn8wClfRUF+LluSK6lMLLTiXC8BB
f13p/gU7rMgF87Enxo6G9P2KGLPthoLdALTd+AJzwVh3V9ZIVrtwELsykI+0qVl0ZUekeNEfh2Pi
IPZfyfMfraFMRFGXcQOmMIt8uma/4YaFT6jLahrHxmP5gxFwIwhTPyy0Rd6gPRr1xCOW7ZRkOW8O
j5NxazcGzQu6A2oH5V/MZqKUzJVsDMWfR7ICRe1yEKZHWfHmHj/3XB91j5AfVXz2n0Vdqbpy70k6
lReOMpy3cWm0xcitPxy7OSQcbEZtOMyOMCQvW021UViix22hlSStjlXN7MOUTLBT2inn0iJ4A+AV
iyqlwepBhmSurgAIpCHhoFylxL9StVzW2QjYNtBCi/b2RPbhAcWWiyRVA0i71olrH3W60BlY3IA2
Ki0OGAaTq0zNg4ppT1qAify6IecAPRujAMkEgOc7TLBnsCoyG4LHtViWyPXEZZ6udnX9ZK5QSO2V
kYi3v7axO6ZjFGiPsITuHmX7kF9lf1r3T/rDpPS3PKa8x5JrEXtfJKoQ8OTTCd3ZWTetvRq5/r56
8wgoXhmaX1QNg7vgeBpW9GdS45J1DDf4wjoe7QiuJ0Ly5rZmpIlm8JiU2kF3OGMlIV/AaUBHR5n7
JvDkMN+Cn+/le1YWN5lvClGx0S148xj9AsFINfG7DrWFDdNTQiVcLavSCsE0bLl/BRrE00tWPmzC
MkhSPDpWM+T4CtuBKTy6nbP5jhRLg8drZMQeaepPFPCksJCZWgQWGmsys2ttHFKcLRJBtT/St1V8
0vjGvpy4/DraXzEBBwlPNHD4VZgXfRGpC5ogOioQUv5OzISWpK4LgnGmyj4R7YRlLWF5B9algnKf
bgzS+SBfJATGJD7l6WFHDerQII0UXijaAYC3Ih2XEmfba8sWDVaTjlo+EH2pKjzM587MmERbAA1F
cfDD3szyHL6dnwjO9WBnyYuopmw6bnOUW1sv4YyJQwyjLGKJ1lBne5bx9j8AlNOwburS1ebkR1jU
Zxb2XotpEwErIjRGlsVVO1zvKA4wGAbIAzv2W8zz4KyP2e9oxVw8cD/TUL+9PcDGXqtfeSoOTFSp
H0ceYKuz0uP+/TuSUxhxTRY0VhANrlNKgcKB3+zNHKWGHq6Ny11vT3X4mjLf8jWKBdJaVpzFQvJ+
xF4VrCCM5oFJjn7Zt6MI/XyVN4OPGp5xkOlx2ygpDebUg0KXBhxoWU8MjQL1TK+4N2DK24klA8IA
PLL+CoU+zc8yl7tKKNBTx4xX6CVWq/dPBIFRfPz9JnwuAR7BsiqBnZtZ7epPLnbUDHcTv41qumAb
J7/Gq97s808uiO6euOYytpyUAmFPmcIzi8WfEPEaPaE8Wl4WNOv4WmM5IPdygbFyYV2I0DJqUgNb
4sh/z66xF8Fp6WmGthb1sG/+VBMt7isz6nkZnn6ftfoTLijn0fr8Owxb7GCAh1d2QsIWZACm3cXr
cJk5XluxlODd1q209vdgBiokO/RiECETTueGCOTJDHToh4SiokRUPZQMPB3eW3xwZ0bOBtKa5DHx
R+1JeMsaUIdq2Lw9sJwVFuy6QqsgVeGLFo9K7N/zPkSzUfcpoao8to3ZmW5ViqnXCs2i5RCgmg+9
FKAxrx8YqxyGDVu//z4en0gW4g0LCdguVyEdQnag9d5YDKm14QpoefvdWorqK/j02d8DvQ5QBWVE
rPi0ZoMZpEhyANGdvXU9zY7P5xprMwDUAfUJFy08yrGhyWWe2Fjz+5H7Z8PTh4fHMC55/NRb/M19
fJl2Izdmd/XdQTT7InSMsABUt4Piy/O3nTVNF6RNMfyqjpCuHMf4BBphgfNvzqOV4WayTrq81TPp
c/04k/yOrLfFGbI6Hli5C05srs/aoD/d6HZUHHyBL+xxUSpkRp3ERf5YLzD0INd5SmyWfBPJn+tv
b/nl59xScoJzvb2kGVhXqgUDf/EjPQ7/JBgpYSlbHrFf0Q/HQhMJE1YmbnTIL+DnwuvPeg9YESi0
ng1jpNknwKHwYZ5J6IV3HB7nqQxHndRLFb37ua5cTnIu+FLEcutmxR/pjUQVHwAvJkVwpgC/rAKj
hEjsGClvIvm0957/OgItYqUWlY0NfUHhZDdjsKIYT9TE7G+hzsCRl9H9qC1vuVNabgSsNT8QRDj9
FyRgZ4wRSArRB18CC48bwkeOWRxrIObVqnxvHo6OcoszQ5E163E4HQ5kPyEVINA4MgOELmXvgNvz
n+0UeJdFb3GJvy/8rMNaUAuSl5pnBQ8SBDvO0rV4HSvXxw9B6A/H4elhY0tHzS6GJ9QLDFcSiFbn
E0rDe8R21emFVbTL8vcX/IU8K8/KjmxvIzAUOB9qvzXQgz856eg0fY20y+RBbLSuTLDlyH7wRlR5
8uzYhu2w1kswwPo5XucKHqffGgjpzAZfibPG9lnrs50MzE/igEMzBzfZsIJX95v3xMurR6AZwTPL
NP0Wghf4w0WaeQ8G36cozIwFYNtzo1IRA02hkwF7I/R+hdurhdJCpH25yPNc/PcOvRRelZGyq3MB
DusrXjlAmDGacCAtETPatba709B02/9nhOEY094djGFYUmof//bmuB268faqdK6rALEOa+oQV22v
Dua0rB5Wwmj+zEyDtLccrTdRi0Y+pd7adLsh0n5Fd89tra1vhuau2XiWp6tPE7/HOJoUVqTI/rs8
TuetrabSxaNmz4F6F6bdcFA0MXwnVMvhsOmToSoperCE7JMDqluQwwnCx63qylw7ggQv2Br6Ddf4
9Njcut0ZEyVtrtB3mv+cWE59OW/wN8nrF257tKjNZCVKjXK7RqFagtu6TCiOFKXoZbFYvjHLv4IH
FtooI2iMHRgpgwM/TZcoAP354/K063WjEJtObI9BTYZvjQgprNDScPSezLPX59O4SsZeR48juAo8
0b1Pwwv+8JZ7LUdhObkWoxq8zS8MfGM553b1aiqUIwx5HK8wBJvwEds1NCIvyCi9Y7sTboy7b8zb
hm7AiKffAuF4/K3jhi3l0nQdr7FNMLTF4968ohcU7DtAPZbHacLYZWIJWgDBi7D5l/xLS1tQ875m
sxEdUK2EA4IEstB6wEnyryGO2EI4KUsQHLl6KXgcsLeEt39JQcsqYVjrFXgb7r+ze3j7C6Rce+TY
Xi6z0ZqGe9AsbFt3kw49Rw5urWcUr5TkhkOgyEjiuJ5pSCPA10ppF1e53CJK6ElcjdZ0QJcaHnox
oWcvLht21tatQCfeERGi3TsDJXUVYCokkJtA0msey0pGAextSNsp2z5MReRt2/0sEz1BG46avW2b
X3ipcWQYRScUqJiErmgTKk+L10S0kjtaG6h8s8PxFazLCSfINs7eeVuIbTyMrczDq5PUUCSuyQm9
Z0SJuMcmGKFGRpqTYdAdg1qWh7VUNH3bw+Dfi4ewVErMtaIYyp015g2YaqTF++e5NKDbE5OBeRRt
ZuAjft0Eyqy7tFICZ6hoWnCjVzONn6h2QMSjxQ232X8pyqDNujIPVNfIPpRPQgUHa6zoIw5FkTJm
YFAsLCns0wUV6SbknLJ78Ps/UpT0X4VQ/l3fpEevaYGwaZDIkIrIQJrZFDIaaqjX+av7dlpfu8+S
neDg0wEWYn/38PJphO5LcMllmgl54KmyQKW8AtpBj/bByInAaHbB++mSWhLpeMpHE3Ek1tZ5vHF+
UWl0Z7zCpCtwEs4GpcsOHUnPRyBMIUmuCGPAIVfzyVzGxZPlSujxUNTp1gCj7iVWLhzg8niJWb9/
qe5tHWTl4G4gP+eCAooYpoPPWa9uHA8syYVGva9HT+T6ry018aYr2un/fsWmwT3n3oJVPnwNb0IV
rKdXm7x7qxCb0MrfzZnALPWHAperKuWoIGIy6WcDUUyza1KfIPIvECrWHlDC7zz3muxVsWiw8tra
ReXq0ISIfzYX02tx1GerNK6IB6S6h7CVEdB8o7+dLikC9m9Tq8FsrfFWxHTGOS3Hc/pUj5lN0K5S
Mlg3Q6+/ZckLG65KygvW7qI8ZuAHoPgDYdtTYtWX5YrGN0ahWmHNjYE/RONleJvANLlEH5p4SCqT
ovFGhQZ2JDcKrZluovLgBJz1XszQ/55lGDMTPjJl6PFIGyQfo6w/SbXVjTA7tM5s5t6LB9tg/Jwn
sm14UF6ftWbcTkk6aDyKiUSJbZ/PyglB7UzgOjUnG5ERQvdcSAOBcJKLvJhQ/OGR6Kubh/U7cAVj
s1UHZIORE7hyvbL4GQDU/gW0ZdhMEJc9pOp2Rr0F+0ZECjcYWzoIgVUYaetd9lAwpSNZs6ti8WDt
djJ6xHrQF2wRSbUoNN0ANz4MVaVHjvB2a+eeSboP1nsV1tAPhGcKsXBZIGS4L38pJHMp3NkumZLE
SccXjtONvyIcg3Vxevu1Bh2U7kruC1LGn+aRC8kmKS2FG5ZC7vWu/FPdLacP8DlCgFYUlkLtevlm
roXD9dtYK9AgCjd59h3ytJvmLEG89p4HgnAhP5IlCJN46/0jRSjLxImgS+mPc230mSvKLNR0fs4Z
ockbNXK1/6KOEM6y+NdsO0shNLa9K15muOIuskqBB+dhAIMVwTEgqKqkdBqq9zrUzeC+OXoljZVs
OJ9CTf2XaPPqX4FobVK2gcTcQAtJy2fZKYNwQaXyfWY5nlZphlPvBLDPYXO8j8XmxjqHV/ZvD40t
9qBz2mehyfTKcYidDblLjBBanp/OMy2kxJXVIJeIkcrBy/yw1PguZ7D0ihn618mRLW4Bw7nbD3HV
VftVKyWL6b9Jz/UfQBc9NtcTHjJL5RS6K4kI4J80lUK88GD0+PXD5TEDrAcCpgodgQUiK8d+EelW
imWuG1+3w17du2nRf0tIot9RAJrEbK4v9/mkJWk5qLGLuzUJiOcPeUH9HDFIdiLTCZTs5oueN1G1
41onGfWj5lPQWjcstgjvjz5ifjtkC6r9M0biLbKqw621Kb3TNS9W5SSy6roKqUzREHbmcW2VDa5d
HsI0hfL6ehnGMdFyTavjt/xI6aAq0fUgI/mvnITPwjk15EFHQ+idun8J8g6riBlgFkkEUO6h6O8A
eeLCZ+rA9AsKouPzr2CEqPK3p03l/SvzJJuvh5C3rRGSlCNSwjT5opN4eE0EoDaQjZo7yAIBYaw/
IXDZpNlelhoh5Rg0FTPkFQWxIcHSPnYX5NXRpHBChldyvq5QdasDKahiUDk/KD1TF2rUhjCnwKsk
62yjNLrMVSsd6L6fTn8E8j/+C1SrD8LSQzDDl7lXHLtWt8QBR4et7a6PMv1x1osyPk6h6cV7AChi
i29Zs8uSPmDUIodF+8uhXukYDfczYuA1QeT0N3k2w9M9ggmWQdyJFgm4XAjD2bdEKhfIdJE2GJuq
m4bOUV+qNZUoJnqegsMc58doaYk48dL1CpAboMpjVkUdO5zVPyAeCYXjHXJrdAwwZuyQ3jil1uk0
JxFyScxJMtxCXwA98dmlazTnptG/GggbLNRODuC/MmwwXpJdRs+0d+d4CYOlD+PY2BUuIdsQuoL2
J5hNqMtsZQ6AkhkaY0YukJ1AIJa1jirlyDWTfW7+tZP9aTYXY99CyE+/Gjbec5gAef/YJWo7t7Yr
1SIRXPzlgjmAJiSIccQiDZ5KStSdC0wZ+HCy7zKyNCQ4d8l8nJDUGklBEQ1wcuQJty1eggs5v2R3
hjBefMCpMjOZk5GI+y+yimzVV610cJVQ4x3+RgH85iD8EdvlTsyuxOwEhqtgtW8KmUTc/qAxdKj9
sXq0Y5m+pVzE/GsYlkrt2ar04GjFGEXIeLJECckfg3hvnlvVtYOYy2jwFWn4MQWmDYDPYiENr6hm
7ZapEyJtl9pKOnIMhtzsHTBuQhSQvHA3wLchosrGDQPR2nHkoUcgEWr5dremzlmlhDLd3FRpFIRH
AZCfAUgj97bYSatfzwOUIOLLjkpxnj6zTy4O9bznETXIB5gR4Rp27Lnbsx9E8Sh09DF5IHD4RaCS
LYa9FbjKrQjl8kma/pMSa024oHO86t1Sr0kNA/KIgmuehbeIN5+cFiwlaNDYIV1osOuBJq0V03da
oB9K4FzJBDhw/A1+MaJrgvbNRRNuHhUiCJQdjhbYkDaucMUBsuiZUlG9CEJEp4jyt6Cp8tC5oWts
1dwQm2sqqJhrciVavE5npqVYL/mCeXO66Fgp2qc4apusSTsk4DE+aDGLLasSPL5atf91hXr3unju
vyUGsw3GgGJxt/bHO5vnhxtQJTgQAptTDAHrEpQCM4ASSg7D6jxhpGzFmI/GWu6mktZl98TvsMI6
bLBmexysLBFZAhF58h4rhm+e/GKOB8RH+qh6ZrcOS+WLPaOpF8W18Eexc0nFDF7R9GIXwwuA0iT5
jPLtbyxcegQgy8gIAh4NcMn11d58QHTofmlWYoa5bxo7QzAN/W9ydT08ISYEHWDz2HAT1wy5p+ro
UmRkj1OAMD2AwntqxH05Qv1tawcLU10BKpgJZdaVHPqr21jKkL+aY0KVD+Z1WVVRvAUcnUbhOcfw
9QC9lL1hsh8GoTkm8JscpqGUJ/dOf65XHOGYVdX/WSGo03eAWeh4fQxLJWvmsn8fJQa074HCcu35
BE9uQZlPNtpGONDzBu7bYC4PyAuAnXqkyepqSw+Lndono2Urjx1/XpJVulvA7XSBKtHLBxRpVENx
E3oK/aR78NNTY5bDrisY75+Nh3PdVPwcVCO4Sj9ZV7eAJ0JKC2NssYflImaHR9X+UHENL92utOBo
/J7rjqeuRTSvawRlXaNCOJRFwv0nQGiZG6nCybuS2rFjo2sYd/oIvWom8PKl/cNfl0WWIJyrVHVr
2dxznT+Jc4MN5gD2IjHw1n6WW0y9paAWFvIgXEwsJj+wmNhDof7PoOpcX7HI6ML1fPJxXTq36Juj
jnlUVubSENyyEw+1BVWFmRaCq7FEtqwJgbaOtbBwYatHLI4hOeCFPGbXHqy09gVP4laWy1Qn9X8V
eNjguaIQ0Pil4UwSe1L8B4K7753Rvp8YMKTZEHScJpt7Z9Zreef4NliRQ/4h4NHvNA6bK/elew4I
TRikvtT0e2MKeIasiThWtse2knOY6WEuPD+H8Zf4yZ4+E85v/tFqVSMqZkRPX4eIK5erqOUoOmGW
hwkuWyrvXVTUhKtkCJztnxqPCZbkWVVGAhSZfLKgDUbAeyABjTLK+hPQW2YVIuv4cqmfrFhedQ3g
kDNtFWNQf7aZzzm1xR8tdqcFnIJGEA1O6nFpRWpJzpNMg/L7l2Vvts/zjj37tsvBx0Ikm2NScfAn
BwwJVSj0ptK5zw0BtZUm7cXxtwQShvcKfqiP63zbhSqNsHj7s9D094w+z1Vrr2bVeCD0uULVQvlR
FeIUrTPzaL3v19/s2scfYhHTaElMHd7vx3bvwvAdYrQIbHd8Im1jxH8ZxRBK755lUz+usxCbfI1Q
jcRLiWvgsLXNuoW0iW028j2/mHR5ockNuqI6LhJS6vvHjf+J5xoXAfgGdfDUMygtNL6ZwcWDleE7
/f7++SURQnzfNJZSXVBABl94VvyBRuZXL5V42POUj21r5uz2EOt20h9K0XoK8A2cXnrsiuP+md4y
gIYWhe20wTcbjEWajlt7aNshblVBADFEoOdXFSMOzrx+hfLgxJGjDRn0KYfhORAY/iQ2olgzvvmp
mUr8ZKbz/HJ9FgHSuSrm6YDvXdsvX7qy5Q3L/lP8R8luy6mBSLpttAnWKc+6IRpdhSMUlkpx1yAi
Ki2TZRx4PCcRDIbe6KVrPd18HyD4ghFCYmuN6bKtGO1tPff4XNJQpH+8GeDJiTp1y7VuG2wMhDFN
YvbICkVpX2GHFrenp2584nsCunWKP7LQ1M1q2zZZubm/cVGHY5NpF6UK+UekVjzfKcoBorUgtjq6
XdnbBsuS/F0FM7G05pOvsCbocEVtWPvb+Dw5rOWKxqXoEOdxOEPzmSYaY0NH3xf7H/ow5LURi5Ek
ADMF+dG7VG2Z1Wn7fI6+dplkVKXH1YZEd23E8FtgH4NnMFBZJL0MInEAi9EKd6lOPv1j9Iehqh8g
EMLrUYsXFedHRIsEGsTwlEb1ogySJgW5pPtujO3SBuU2JZcZWDsochtgSZqbBdND493Wln5m8MZU
U0inh6MFiYvbu4j6wKkUdqsw9FhJU3w1P22NmBxlAX8afrajY9FnNcRbjYjFOWKc+Nc+VQg21G6N
4/bzjJQiBDFCM4zDUFX8lThNFIn7BDnZy55PIt5sFM+jpGkd8Xbuhr2BeL+EBEy+ktwT9xolpheW
guqqkEYj8TF0bpGjRF+bl+yolRwLx1V1pqSJg1BcyuZPecpUifGHchgij9MRrV5omDa2RYChUvTK
dzXdQ665sUv+tFjaDWHw5qHfik7yCxTGOLKEKzbQK4UFucTQUqrce7afy4OGR4vPfufCgfGJP/7b
zisS/qjgBRIKHqgyk35pwhK0iLr75dW2qqcvCEVrUjNnWq3PnO7tA4SvZofp0EynkClekgnltdBR
RaUN4LTi8lt8xn60hi9yM6Z27+hvncTvckWHj9DWU2CtCkRLiYBhTC0X7eGpms5FYHrrWcXVsfqu
45Afntw4PIHnTuocX9s6jExD54tYLX0gkceX/RCMcxH+1cBr3KvGJbmggH8FIECyfKQiMr0wvJGQ
dvHnNU/PXRt2O+mQIn4WZMO57+UUG4uClhfMtXNoFLM22qTLw6g6c0w82EhMKqmrVQKq0Rffj57d
BhNu/RxMv8ojXEYfAtKWbTBjBPX2CINK1N3HWBUCQx3q4aYjt17EDNAguaU45w6c2JT8StQoPaUV
O0isO/gBtyEBjt+yNsk7Vx4jwyTNsmJ/n1+5X9DzTfAh51JkUbANBYNcBUD8editJFb/DYJpIa4f
mApnanENm0cTgmXFcWU+EJNeZxhhOeNiH0QHJJgOBipjKBQI5EG6jZF+d9o/W/4B8JcU44+16zII
+TJUKGBK4DpLkVQ1yvsudS8iW+sJs0O3KyaoRu0r3aS2CvKoDO2SyjvDTjuQ4ewe65vLqU//goJn
1nYbMFD5FFK0ZEY3ythXbVTfwkccx/O4JQ3uA+/o3moXrNP//vdZkzob3l/Yu+j+/vIy3UalsD5D
gy/gL1ZssbPWWXtaOTe4jAQpZyvjQHldAVQHJqVlSGwPSIBiI0fmhtdXDNoIpBy8xCdODWFVhHRN
izGea1K3b2adRCds5HpZwOeKznj0vBgjEXyd0UK4+CLbPUgOvlqWjgKubITjzO836sus7vi/oSQF
NCaLu/pqpLyyUVbv889PrSg4tTFfFOonymEypEbe31q704FTLzxCleUotl2PuDR2FLiMOyHuKypj
dFuF163I9LO12DTfUFepHBO4e1ltnJ19GTdCTr+SUmbmMszmRs8CkLqO/NTCYbYA5LPe8bfeNbMS
rZzoqMAfJUPIUcQMyQTWhI1k9r++lt3T+WFtFkQr08Sp/Q+l39Kjc1dzCaOmjVI1NTjElHXyvoZ4
wxrQ4FqA/3IsjCAmEQMuivNq9RXJnvWEV0P9+KZxoNdANC9U2UwY121L5ND/mFpSYIlivlKWIWb7
Ua/Lvmj9TmNYQCfMUszYrX/xC80S2N1MWiWDSJeYXXQAt+BOQx51TSJDODM5E3abzrKuqJjN967v
u2OerQnZtEIHvqaszUif3xHQOp1P+Qn9BxiRMHJldR+oQC7QTn7QM4DpJyuFB+0GOWUC/sAFJtqP
YjRdwWx2uXOAX8eH/fa6KWz9tLSriyp+DmmrnROi867VOW1SDIMTcUeJ9yTx/+2zzdUeulLp0iRT
XLKwoFiHxZBXE1PYsF4DJXxr4fMVRS1vAKDfZmG3PrbyCarKx2uG21VUoPTALADSqYAEIhZ/AORL
cII2AoRRnVHutXS8sWAfJAVsutQ42YBJCHUZMBhDrQBatBmmcbcdW+/q3zhSi4YzfhKK1bTs47IB
O348O4BqGkMX/VIS1BygYzIQ4mR7oR2LxSAii8KEiBnLPjVtISuSn4WrC7i6al9g2yNqXvM7NRIz
Dctq0iErR5Y8PBD4NjTr5HfpxEctuoTNXexP0dsrHKEDTnB0wTSwvy2S2piEv701Q7tsZzg8pdHb
owSNe1ClW+UoPf8CGpE1XeX2hpjdMw8etIOYjVzoCtkDa7rNOmkOl42hpzaq7JTJQDEmMWVlawhW
f0ZdzKuZCVqgPIWzxUHYtt+CJeGAYXkao9Q5SrhWIbz7PLGvUN+UU+giKE0XHd5zXwbiQ/wjM0w3
XnD1qtJIEc1oW/N5wNAvZTjEfhQhp3sLFCNOYRSbcSeuLADLlPrP6n/Nhluiy7ZvkHUNmgH1Hw+X
ZFR7JPjSxgFlKCHJf3fpdfZwegLGeBLy8/tobjIr7PxxpnOU/M3IWg7XPnI06EY5IIg7U1ZVSk9L
wuC7kwOkNSChWvajjeYG6q0GlzDnXaTGsbrFjRuc8WZwNhPKifKeSK4HhVknO57ig4sGFw66qktG
2rgAREvCHEyuNOm0tZQ0j2mGsev31nMBThjPJNf47KCG63FPMgiqQnD6kjBYdg7nLCU8DqiAbZY3
SQnySOhMPJ6Dktsfxot9HtEtu2Fz9HZspPaNOaTXEDRcoVcWRduijBZoz8m7xQFFvjnc0BdizEcF
KMhayUStvYKpQzSo+lLc2a4RZHHwHklw2gqQCE6qIzQMnB3+WZ05KK/ctS8DF2N/GnqtC5RaOzKL
UMwrDdxpAt/ZyJjxOKe5tse9RQYBWnQoe1UJOaNZPitb5VisKnFdsnF1k2kmmpPs0z0VDZO+AUor
Fk4sHUXwFcei/4l8JCyVi7+ao0dA8TNiezGN3+MQ0CxQJdNgi3TmEEwxriB+3vuT3ZjZzp740Btj
x+NId/0hav/3S1t6795JrLY4Yz1THD/7fM1kCa1V8Lz+snGQWDM0SFwMzW+ckEaYrWkC4ZQ+kGLy
IwhE6UQAeBpcEVwt61PAbJEmxLpd53PArR+X4SL5tksht7W3Ga7YUq6Kcz0xsRa+YCczof8n5A3K
SYJeyCV5bNV2Y6YMY5NfB5EqQhV/d5cDhFW9TnJyjCtLVyWG2p1Vk+5kQIDJFee8cmddhNLNyzym
LFGbsjnpfQKxo2JW881DPDAM6zwDOo6Ii2mO8eCuO+WUQi6yMvsblCRHWKYDXbmCX97LDFEl9aEw
f/eR2p2yB4z+gsP1s2LzZvqkHq9e6bIE457aKAX6pIArw5+8iaXnK8CCBqBYDk/ec20RJFK1ORbh
uLAtmtHJIFmFrRPrx69GVPBFJrJhYVysd9VH1kCWU8md1LX/oXwT1A48o+clENaJCdUBHV7YsB0A
Sz8q6oR5uOYwC2IyvQY9RDxAst93e9FTmjOwZA68zehrBeAb5sJFowyPFckL4yx5YCOzu/qlM85J
TBX+gV5wNoFb61samf+E4qZnEj008W1ZER0aVmDFsA1cmjV2/oCpfK3jiSISsu9NXBST/q+0q/RC
WgyBT8rfJkeHJJ69GaHqNE9tpJwv654GXxZx11F0Cu8w7py3vK8FjzuRaDLEhhFLTTAZ0FDzWqQn
lO2wPOqXfMKYgvjlVVZ6AR/BxsYRF0rA8BKslsVx1upcZE7SSDV/PxnDlCjJq0pRnzRe3vVFYkXz
bwIrvmmtzSI+7K/DOIj7knYxW+jjClw0Up2BlNp5oFG/du2e6ZLDdCMozHAv6HyOLMPh7FuW5z9F
WOv9QtDoWZ8VsjUzK/HSka2a7StmyO3AxOKs3EsDJAOl0yyunt5x/4aJD7+psuXOH85bxohRS8vi
DoTVrfQ2Ca0r30KjNMYBXoCbLjMKUdtvcI+SzCgRHxe8QZXjvmhZzZTwcQMIkc8K/lnAuEMFmFIx
MJz+nrxQCfq4N3DAXsLOO57rk25c392g4b2Cq1iLNSwW4bs7LOQrfUtq3m6jHc0rv3/+Lp49+6BN
/Sn2H/1zZg0FGIw+UvAzPnAqWbkb4Qbx5SSTQdZWZCi9uYUO0iCKmO7fs5jMqigdf4u0w7S0s1fc
wKOZSlyWFGqU6HFfJySll+QpKurYsZGSpNARwI70qhXlfypQ0pUgBdcIJyM2Y9dGJIV2cLtQiRp9
5jazAdNRXOPaeDnhUwa5CojnOG6BYhGHpD4ZHYGlRAepTRA5vUIZyR43e/fFcO0DIM7nrZPo5AKR
dWUS7JEFJUB4pVu/7UN3iMcu1+7Re8Bt9g0/SrrK0hNmM4dxMhGkHesQxdiqE5L0H4E2B30hR8as
EZvA1iXyrYXZCJUK+h7+sKEtzct9rxmsarBcqKwvXoB6SZFoXUczuym5TxNdChqjPP6L+plc3wsB
aAn6+zTF+sUhaTE7WV0e0Jmb3NawYCI8l0AQMFjfVeV8xAtyNv5rXRL1hkTr7ggVHmG+g7Y8Aoaj
ihdX0qlU8C2f+ant2KCP5bcOQazwx9z0cQ2wrgxeshmR4OJiiuMAQUukmweCCWtnqxFJ8NE6ZCuc
rDDSxku52+syU0poV0dEqZoGtWZ70ZbQAjZBk+nB9kCEn5Bam+zgTTFnWVM4njH2HsFZomMFsRzA
4/8vqRIe6430Nr1lNTJq9Uus85YLkao7cFHvsw1wiSicsbkhhG0KZoXmvsi+ADeZQJ8GeGp2R/mE
dHbNM67FnHTdY43NaL1eav/UGDj+rEYDcURsC6QD+cnJ/KpTsv+Dizfpe8M6be2hwjqXVDE/9dks
TgBMh2LCsLKMiEai4/dBx9bIgQSNyOOAGK3xVIzfgHNe9/6KdpJpkDmPJQGWZ+vpq4J8vC4b78Zo
EAD9Z3zGy2Jviaytr0Oxg++XIjFdOIedGt/5eoH4KUATiGgKpYBSBZnlxlaZiXKxzF/+U/0mpXyw
Yj/DSA6AMfzbmTnyBLvhoprJ1q4dCRCR3pe9UG5KGU8aBaqUfx/MGzpllF8YlR15JZyMN8v8dw+e
cOkhnMDuHJcGVSTDGTLSme5RTULl7FknBC3m9Ux8runK5CJ+LHR8mPWHTsBqjAjU6WMW3hq5mkWS
jR017AhlfQuiEU8+5V4rN3fYE7EV+OMJoJbK/rjeJ5mJ11XKg5bHbegrk0ZPpezRhZngfkDOf+uQ
r9TlkluJs6i7bk6Vo8xFMKmATA38jz8HmpXhqszd/t2AJtmgAyWGO3Tin7OvAvD53JRcJtBlAdLe
7tGw9iZ8/dv/HnT6p4aDWRmq8Ay6Qb0gPwZHYZ2zPbGUH6m/4akfoktqwgQd3YQhvLxY906SpkyB
Axm5yYI1S85qP+f6QQw2yFx7UoXCjpxlQRM3lbH57RyxQhBryllq8GeruhCPknWphjCXYD15+PLV
BgHwQuNbG7bJjFeAwWUIsLK4M9C0BjYgv9fv4yaqnfFddJlCzU3Jg+UvCdAzlTEsqmXRQ5fhX10G
FE28X4kHXTVj1QWbZLHYfpR8p1bAXf/WaI0McZ91LttJq1xB8Px834d5C68fonUg0+1nXTG9Bu2o
6PZMMy9XUQ88xomCKvItRCd/8GJbURT3KhHA8onqgwgdQ40S1TOlPRx4u5cABR8R/vnd46K4oDH3
pcsgIP3agl+d+O0J3nCTqJExqc5G/J44t3+7Z4bPnIcVOSrQxlOeD482NHNokHWoUfy8ZpB2CXkm
9yeDYsPtzCk09yMcvsP1GlKbErnlBshLZNnT4XiEjVcBay4drC3ypXYFbyPGAE9yrKBCWo9+lw6f
pZl36OvhB6JzFQubwPYcMkUfsueI9t1UjmrL8u9mmvalLrHyUcxmyz0fo5zInUpslNH/fqBVpUOo
2xiOPbQHA7he1Shi4TfC0x5HFeVMBFO0OSupl4m9s8rWZJ84sLgaimm+aYbqwXgTqB9woK86Hpqx
b8CisEyWmMx0onQn397fx+wWsztFKFdVWW+8lXpZwvaJ/fqVEuY9L4ckWx3c0BG0l/82jb2pEI5W
Hbk0TVQ8+iT5m/mdSsSKNxiAuhrAyxo9kt0e7I1Re3CRfQIM1FHdJXmVdozWfOh2qXdTTW7B72p9
7mC7vtRJcdiGf4WequlmmIGSXOodZLhIoDSXu03YPo/AvJisoBgRqPnI+yEfYy+BPvOwBLz2cLn8
T74OW0tcYvBsuqrQGtS+PBqOy7076kIH+GjpDDg0Xfp+mLYxH6qZtUujtAj2xgqAasJmMlAMjgSP
Jdg23Iwl1PiITRY5AQoRVov2eCu8KLQZMSVtISEg6hk2sH9bR8D25y4740v1GJNvxLNFL4BSTF43
enjW9s7bEXM+Sd3rlqwIL0RA4ulp+S/su2qD6ykOay7KxZiGOTf0UaX6ITt80XQ9rEdLP3ZRMPpa
NQXOFyEWjvJURfvKDmx0gHtdyQhb+18papP+6ipSFnKOo8yIAC7XH0vTEEOwaWwvkROQv1JhiRYH
cj4y/QoHkuk/rqudxaffrqAc6CH/Xug+fUUKdNVg/0m9G9Z1TV6q7UgBenF1DQy3k8B1Jv/twB7K
KIGvlba2HoqH5ncqGw/eMb00/Fv1befuFfH6+Kw0Fh3JcryvTdvpZUuKg1dbzfpjfWx48TzH2UAU
TWNiLBV3S5E++m+Q2z2u5qc7OnYa9BmGiw4kmIU5o0/WZA+T71PdoEI+BgAZtim2IfZmrXyK2O7s
k9FWrJvDzLQjmEXhnaOJnubLGF99VKJ1p6EXybFehueXV1MEKQzDc6BZGYZLRBH3ksNTJo9vVb9G
NN8w8GBmi1d+w86FywpqUMB5fLj91FzfOc3ZQXzGvaZZdI44mQXOtjY9nlUtkZrKrnJv/azuV+nJ
H9zS3I4G06Z9bMx1E7BgkeHWRp5Cf/scm5RLxi1ELfIF1Gtw1DoFV3tfSY7dtlZpUw2KxNoE9LO0
WY35G2WrUH0I3pA5wkRt6/YrA2wIOSz/Z5aDfrLG7IcJ+64MZJMt7PFONtptpI01Sx8dcLaR91b+
ZFhvG0GOA2EJsnJAEa5BJBCeThIWoohGgaV118aFalLOzassxBnUXrml68zpvSexxUudl62m30sF
8Qpav3hU0maDtr9EJiIvsnyQQqfNO7nZKpApa23BQiqL5+fosPafjB8KhumGiUYVw/ckir4X5BV6
2uwzCEjmjIVd2vbQ6aA/SC8jLHaGf9yY/ItgSgXHAPknHJZvVbrzshdVaOicVH7xx9PyU7vf1WR0
ImpbYiOU4Zyb5F56WeZ9Ri2s8JQJP0q2CDUiJQfCaRaz9J9Cr9Pq9sPAeZcYjMqHcfSLS/L8s/vO
rjv1xajyh/mDna2wZOwYpKSV4IG/1+RWor4CTpXUqXw6gMXSjipdfP1MLr/9oS0apZBz8+7428Gr
srgchAQmtXMWI3MQ237MlWT11qhIXasOVKBI2gWKOfc21Slzd+tSPWPUAM9tKD9T+SJmV6nH+19Z
ErffXyNGO7cAKB2U390MHSchizTuMwAS6OmJfdfA+fL5R/m9tO8AnTr46poSdra/PbL2XxYkC9tO
96Gds5hev7CNpkiTVaB+EE/AbOoQrdJnlIvDvrNdxRjsalUN8CDCpn8QxMrj6PoXuCX7TlbfgVgd
vGA2HR+DsXx4QQojzvjyoQuZQKBcOoWfKb4HsF425QLvp8ifpyrKifIzM2IhESsIjzqXJ5FyzEGs
4UuxTD4I1ThD1cMBXirui8Dk/uLvSfTquzZ2+nIkphWpHfe/FuY/TTevwlIOHZGS93atP+i3gDSt
fX4tdzHovT5JKEhPrcHIf2ZZoB5M7VURTSrXYXUIM5yL3earQ/aYBMZqI+TqJxMmTzQCleejHe+4
+wvUX1dhJuAPlwcHOYWIYJhdkWBvotchR9dn1bhrej1+UqOellpac6qQflF2edk1KNRsGxjdxoqw
4zXshfjZrKumCMtTlJXs5fNbQuqGxaolhTf0jTVotWmb/C8sZeJd2kehdHcMxjVa3/OtQ0Ui19ER
Am5DXiDPT62QmY6yWp7FyZsAuG6xIUOOXnALpQnUBO8K6/FKtlp1LUt0G/Z/AhTN3bKVFYC91eYg
MkMnOywVjeR2lTRr1DcYD5X2f3akHrOAjmrpHgGJiYe3333jSNQFraW+17bC0LvZAUWBU2W54Rob
m7oSdnC+E1olweMpP3YXR/MJPOLTLKc8iWR46aDQEzMd3REzTSIldrDt4DGodCOOKMT8CJCXBKQ1
JoX/yJAgu/fPIJC4UVmVTgYaeyMDyQ/OFnkomyW0OwphDvaAzDnMY/qGBlnbPv4ph2m9UndzQRiw
0WQIlCtP66bBl3mVkZXwk49XJWjBIARwdFCTCPTPJWI+RmprXmjZ0yUJeRccGbFY6W/tUEJjDhdz
5XnsCKR+EbkvZ8YVgR2PBT0UM5TQ5pCVgfGiPHYgOI2GL4KLH8HLdCzqMFi70lL5l1MQ8o5ssiL8
BhQA4Gf7/mM1OVJcch19DhPMm9fY4llTv9OUPKO85sD6y3hTuv7Ed2fDepwztEXzxyHR4GP0rhvL
u5mpVNfLQGC9ZXyfRVeDPstiCfC+nfJvVRsAqdO84pmPNeTeoWvZOr41x1+28rLHlarHiPTkPRb1
CGn8ExghgZwjReAg6MwAtN3CXbadaXgYjeKdzddURD+v2NGR5LKrxlZpBGS6MfwznP6IhM99MWam
vKWDvRNJXcebwShK0E5Od8P4fwPnSb5//AEOPD3Sdmte8FAO0oXAGtYH7vd+IBBJARYmW4d3q5T+
DpYmRNYi2Bi3B6LuWxH+inojs2VNnthYRyGrp2iHfGOQSRTNkZ6wq7e0aJrFGdeG5Fvfq5n3av0R
H5WJ8/0ym+TagrmS6SCwYHU13U/E6TBI5HhwDdRLFb6KzMiA088NKDfzpYHBgt5+2dtGYMfQdAzI
eckij2xRjPgDnHQ+a+QhzkPCoeX7a+LnyPbzrrbZ+rxxhX1uyzAHsMi6pkgMuZkhmYUw19LC4OsH
rHlc1AeDLPoCvwwCRcK29lMbSQk9Wy5h+inJ4JyTan8nBb+Gtc6IFHernnSgNSl63FgnGO4YFMwJ
ofujm9V/mlLZdAWuXT/zQHBmb/wfRFmFTaE7LGMqeIOQLSyEizO9+y67yC6iRQ5ev9E+tt82Lwtv
rNCCiwO+WsyyC5bi1SEiL2sbWJcsEwqimoBCfWhuhYEi947dZtSY4W4FUztII607gTDHZ+NzNyUv
NcKefAuDWZdy8psTCNZ+pKCu4jFZEN5DEhkdBstJm2M7yVqigKUeD7qQgi8T+7ZyjOCIRrDda6Ss
sO1hV2nguLDikgxiEw4Kxm6EypX8++CbFKJHvF5KvTKDKR5coUgmlJcf1EfP1jQB54avd844bfup
pshgZUxrQolu86HCXmEglngIfpOzv3r5HqZGRXNHznpYVN97bAtVcTRbuZOjY0FOFbfZHcI5uuV+
hRoWqfCDwo+OcDOJJBMNAMymbhwpCkTr3ys800fUAR86dR93SeCNBcsDLWhIC9fjS6HVCf2kI0zY
pjmqP9NyGiiXy1lXUygqIwUDdw5QJd6UHfT1Dv7FXXmqw1LC6ohqC+w+88H/P9uEii3bCidrLiYt
bIDvs8mVRTgqYMZRKV6sf5yYJ8fyEWR9o8Rr/h2reccvHgNRRAUEzrHmTh2aJIJGnxQ+fXQMDnts
eIklhT/hcQ5+7yBVm7/im4C9BRGkh5isfu3ZmD0Vhoo85f3fNL/GgwWL/IbJtYbx0XgsqWlLDPOq
NuDH6qYY9bpoWpVRcv+zrPe3yA85d+PUwuD1P0W5/ilSS73IJmpLzQjrvKwvt12JrOvbtIn3F5Ee
UvMxvzWKOGvpSTcuwpuPgGmDiqmRgmdqRYktJP+22t7+eMdnxVmpd5TSda3QDhmLUKgEhbXcevSz
8gGLmlb0XkJtR+PrkDEic+4JOp3Tc4+cFbm0eltoFS8iSstd2lcG8Z6LKCcXoUrb/jX+xkh8RuZR
9PWJU5Ny3lQwQdsgXTWqSCqikPPZYw5PjTO3h8dD6RPHD7FFX3ewf8i7O00Rku0plO7E+SgOAeQQ
W3+dE/fezLrhQ6QwPPIHTsMugflkP8pcU1WNFXOZj/R60FbOVk513MeRUhJ5Ocnb1a7wL+qbOs1O
g/StYTte0szRSoUCSB5BHyUiFCp7dOexeHgOBIoBzL7U/Q3fn9YlWf/5D2JGLWaiUBbyqJWeBfc8
FMiFtE373TNWHcCjW9azzFAixv+7ycpO1vNhc/8bwM0gZ7yMKrbFh2c606U5qh6N3mDmaM91F+Oc
XdgbaYMwK+9N4wE/0H1sUYUEnuNcP7SZHgO2B8f9+AMRktbYENQ5i8wMqsUsZ+BmNgGvjZYcw5P0
KYBbQwv+Tn1rBe1P0UvgTFJyLz2R/zW+xvBtP0m40pkbdBOZ1H0BbD0za+nysQNHOWqBlFQPjRVv
t8WrdI8Z60JLy5H/BZWCaNzxE0SO0/ZUVmRl/iIWHTvjarFmyu9nLQeJYFRzDz4q1jePDZZlK7Eg
0H5eN0sLL97R5EFHIL6Su0N1VigaYoRC69Z5z1XtVdDBtS9SIVSUaJ7GTmu2X/Mqmc7ifNj3vxN+
mjF+wXCZzM8V4gvg8Egx/3I7xUE+QHIK9FSyBsJdz5nB+asVev96RdEhvNbdfISMhjD9lRXSCn5F
s6Lda7d8mYuYeMgCJO+wyJqi/hHxX7KEw+zt9f+xpty1laZrSMXDypWba6B2znclEfygG0wSvGei
HO8aRbbZ3bQd7ERN09PCX3L7cE7AJOoTvPT7QoW0NbeBkvc9xYrM3q6I75QNQ2jRkzrv/+/qaodW
RzteYKhAb0EIjeTeBEkzSb06agQNxq7A878+UTkjJ61PKOHHamwVMRC9qzDKranZxd8XrKw/Tl8E
MEXiEWMLeFpK0RPD9+a7c6QL+BUh3KZMA8vjuLxLOqTwjgCVI3sJf7rcbsOKxhS1fuktzVJ2cV8J
xUKswRw7VKBwlbtj7lIBqo+F/p90bhsKr5ys4ajw3jQNZCmEpCnSE1bmOUc8mxJS/JgUujOGSN5s
UmuvPLZ49m+CCVZjm6zK/y0UoaSLnGIJgQ5S7qDvT1605CNJwcS4O+90x2Zhv/HRLtnreiASOXy8
PMM0/+CZW7WIX/47dqICUywXVG9q9BVWai0U0fg8kgMZmHKvy0Nc27NwvhaDSj9ct7ERslCM8UqI
FiNex6fwjGRmfy0TokC+5q/Awhgpwsm1qH+J3JxT6nkcpfS2RDxVTGFa+eVFAcSxtGMtvaLSY6/h
EIhXav0Ej6e59qUgAotAsMfXlfPm6u2KAogTqIAHJwMBS+VpvM4Na2G0N7lqgccB8vntW51WuBhj
rcQpCk5jsQz54L0GSsI/E1NjGMqnZOmhpplH+PRlK2Pp5KMVfJZVaGuCpk/PQLiwjk5Vglj3nbP2
g9oxywpMA9cWH9Bldb+Gdu7BnzGrxiwRTUG1Vs8YNJtpz/h9PnNULgmShI4R5pIztoWy81wFTS8/
ZqYd1CrbHwg43dAzFPuvHC0yPuMwdKjiissko7dZW3Oxblw0dYZPAU/iiRbgvee5R97zEPax4W0L
JjrBf3MyT9GGQwyuapPpqyMtZWj8JedQMmFwfvBWtRaYszhzCQ8Ewbq0+K9Gy3VogSDcpS4yCmqD
NrVRsgBrvQ5mkn0hc7TViNDFm1lW7XfXDquJvem5Z+mhtX6qzVrVphM6u5nPtEblBrJsy4wYiN37
1IjAGRwDSh4GLXOfMQmW78ZSVtMJwF3m1y0Mn4T2Jys8/DYdjn/S9nXidKtkj0prIWTi3Eepi+C3
ySymg8fQVZeZ5XyAqOzyrYKQwpE+52V9ppBHUtUrFh117njqqOFYJZZXFP7GGB3yf7TNrEhJgSs9
KB77n0rPwKkzA2dQP+2k8i+zfuz/ksyAHlCcVN8XMqD7RroyYWKpvq6uBqdGHnoBgKwQ7wIynKti
xEVwVnE6EG0Z/fYk/NZutvwhc36f4bpkKakWOrITnQGFgKBY0ZgAk4rcWNAhzkDLP64ekygejNEg
sFglID0UWOwJLYrQ9JFYGswEQgsWlmyf+GFF7mRJmELTuOfyhhu9Cx3wxvS0alqnco6l6dZvFVH8
AGEFEonQny+o6i1PaBzb6lhzG5jTmfRhObhcoRFlmwEn9oNc47+WGlSbBISKVW4U1wTnBP7qu44R
peNdi+7vXKUUApDYuIB62L4iH0KxT/zciRK+s6Klou22D6qV0moiYSh64PedqS5/M5LZJHg5yN/f
GnJYT8SV6El9cUTIvwVGjOKAsVhdJ/+IlMtgU5runZyjobNNsuizgAts8N0jqcUlRWpqIEbIcSMg
k/DbPmiSOzoCCnBiQQpo+Py4hVIP0sFXOTsOZYV1KjPvIvXQyDq2EoJQm+vboZImI8xQUCCYC0Ra
hhqmTa0axNMW1deCtkJE4VkGQe2NfA41UOc+e35lC1SCdgHFKBkrl1JvIbpxuX6BHBVhOzL9ZOMn
lF1/wjFwZoR4osvWYznCU6PzysczPp07mM1VzbI0vHbF8nfYyE0fwvSO1jZFb98cdlE7cb4O/0aW
dYT6b8BtaBrMJFdbRNfuGAqj3fZ3By4vu+oyqR1Pk1LqK3jY/zrDs0+xPIpx1jojcJdyfZ7XZYPX
45IszvQxDRE5ANa/3ZbTOaQE9JmHMK3R5jRNcWdTPstdQ5Fn2lnYE+HYIk9a/I7FWtfpPSlJ84ub
7LDe8FnnP6wp1Ci+bM6SPZ1GKO3O1YUJjjrvViBKj1rnRSewpxWeYEVTiWeSsmTiAFENJ8twxANH
342Oo8/aAjVUoB7Ch8vesCeExKhmSgd0A72MLMdjlOsHqdxrDP+nwpD0N8lGm7jA1ZtyhEcc2iGa
Eojh2AX1TpIkRSsZcrWQRfQ2+9llgI8W0NLa/exV/g9LHsSypm4JCHvDahaRi9lpwph8VcPu6EpE
BUHCMQCLe2mOxVxiCjK71kUPUiM5oI1oZvDSKJTVcwq3b3a50oFBttLmTOo6M7zb7+zvRZKljQkY
chgpR55xgdPU7JTF1oDkV3c3X218AsxlWczZnNg+/nFf+ZyaczZkOAQmkM51F0T+kkRX9PJCL6BO
dNqBrmRcWI+/twxugv4AxKKB6A0LLjjmHbTyApibzdsltwbyB36yGo+IZ9PZ/3oTV1BmCMllgJhV
Jvgu8EvtWPEyDzNBv2r19vdUi2mL1kWEnd4xeW+vbLkgZtxHfS3VmAA0/su15uizV8u6ZD/iieok
oEJhFhzy/NI3+cQs4ZYUVhAPLXM3fLpsW2ITtFmHo4hCGkZhw03PVDpp9BI3OfB3foxim9IPwlLh
MX0rnjUL/JUuuKWaOVj6DHDEHeEXsrrME/R1yyJGGEit1EhzXaF19E01j6AtN/zOGL2oMOWUqdAQ
KHpa3Z68h074xiOCNUXxLQDeHfKsWDNPR8dqJ9euh545aE2/xr2Qd3g4Wsv1fpuqvNxtATUtjEH1
GM0PgiD3B4wfh5rPDcEnk18RF+cucnq0qE2aKlq7C2uM2Ed8aey+xSpmaWimZxeXrgUb5AoRMawi
Jrl1w7TjSj9p36jt/jW7x6P1Q2KeQ/hdx1/8scd2OEF07laDTd1pXtLPLWHyg47VzREm6ZRn57Ek
t7+/v1ixSBgH3Puq/kIIHptLxGcgQJGzQkS8emz8o21veITZN+YEWcgmWhjmqX5MmVFB0dZSU7R5
tluj2lVcMBoWYZgz27RYmFI/QXux9bgSLjr5EI5bftucKPDdtW7RV2f3encTt9h/JefcJD7Uhjqa
mMB3FuKuqt06SlG7DZjPcXMzqQPdUN5f+wPVcATIl+sYT556PKW8ySAR0FcZmDbZknOdyitSXy1l
CHY12SPBn/OgUWmZfKN6zytZzsI1wZ7mRRR7EZLW+HHOSG2s61hjevKwo4BhWiEmnWJPZVgqc6wF
M//X47wmycKY089uQvzXaaO3X4Lje+dGE/7jw5VpGG1VAzdhnpLkOv4KjaSpayIktxVUD20Qn0W4
szdKefyNGGdgHDM8KbCy2g8/xQKbxRyU6UIeK8ZtyBGphkBIzMSQmaPtpSMkRbsJ43hiR7CWWVgt
MmS3X5O7p33RxC5VsGYGFR1/vQRppzL0ewXwU96S08Tr7mrBn2KbBQKZyUBId3WZup2KpCYNVfJv
QiD38TF2TjLY1RnjlODICb9SZWjk/syT/pCHTGWm3oLlEzLc7/yqhOp3rpXdYGUvOTTum5TTaf4T
/2PEVpuZtQZS/+uWKuqLvk5a5BPQjlzTIlx//nod7NAJLqC6wi2UU0I9SVww8I/+0nnzLRUI/QsZ
lPIyTQdsE3E+XLNv3iG3X4Bpv6z+7kSuaSV3ck0CQyCrcud03H+2A2bOhEELygyN9GfuYjd4forW
Q6Lq0MvEPM3aRfydLERaPNIS43dEktrq4ls+KU/2XoXFC8XM91NKaiuztUj06670moSpJ/37Gr1K
DOFM0qg3p6yE+06oaM1b8vNeCYMqMOwIpch3sDlOOJdbk2tyORLbrKThpxNr7bJhKGAKcxdjMmVY
YTNnhe73TcIB4rYmBbShgz+xkU6hn7hSQxIYTC71Ds6R1iZGFCrtWb7jfEaiy0pUfenqJF0Qdrsk
cJuPXz9DNRjIBtdbl1U2i6lKyhKxWaqr/X7bV3ceQ78MTQ8j+BMmB1RSBiAaDZJ+s/z453KtTeDY
iueJkI6AQ2LhWx2j5GqKFtI5bu0X5kEChR+/u4G57qrekuR08z4udcBVNutJYdsVEZUSil2hr9mM
VJswj+3FZXOEiHM6+XeFOrWMYyWtjX0iOFdMgSgbyk/RGlsbgauxLb7lVis/9fxl8IxtJUtk0XME
TZP50uyt1SIIJk1fkmr9AdH1JOivvDZpJ+K1VFIdKr+tjT/HG1JmZBHYpt4XNioFma5mAOdaxIqy
/qAu224eWU/8oSyRl/+lheZErYV3Fqv98fLU0zfBqqfyQpJQOpLOOUGCpFdamBCUwdP3zUSGU/HR
xF+5n1OZWnXkfT+Zfs/KKcDgZMoiL4Ip+A3oh5NycYUuj/+ofl8eU5aZQ5qmb26+dIydKvblzGNO
HGLTCwm1WhL6naa/hx1Z/Ltqm178GZeqgsXiPef6WulGbyFUyT7tOVzl6IVhmwV8QpnCCFZWn3/R
uqq2p9ktSZkr8z7pfcSB/zDMviAgwNGySUNBYCjHoW3AiQNibDlkAEvKgmcPuCrx65e2jZ5s8P5n
OKhrN356Z3Ks+BP0u++dIy47nVLALC0g9c7CXgwYS6GNEcEq+kKRwKkFIMQcGEBgQr8s44+E2y0T
0/2qXW3UmD5kG+c+gAnjos7sTlpedwyG9JKr74mPMG9hkX0WlVKFcpacb2CwuMJLB2bfe9Kp/HJB
IDqMInp+DsZwLwrC8kG9mc2XDHQvQLR6CQN6OcbDCu28411s0+KanrA7pQEHRqS9Djk0w+kOcE+q
W0Ev2N6Ad8FIyCLwtDac1XBfaS6cdBREiSRcTGmwFh/Efzk9icQk11N9Oj+YDLhmg47y2mSnOjCg
D7w09Zcel4TTwSsZb92HW7e1JD5pjoi3T/CLwGQ3vjVn5PLsTYbK835UTGf7SwC3dLxngk5tH7yM
uNPagzmbJzsbm032RFiDCiPbol8PegQTiCA3JGstaivfITZk0iAVXt8/W6G61Ce4TwTCyAPhOqQ8
I5cJdyCTtvy4pEn+/+KglI0+sEgug6JmTe1/+ci+7WNIam11OQfnIazrXzSdh/arJorELDUKtGUX
rbuFFykP/2kKOT/g8rO5U9CHKFewbS8uqvJr9REVPbrdoU3SrVFJvKZlQOVgk2vTg+fWF/LYXSpU
/IyFLbJ+JVYJPEaNinjx8oYf/Vprnmu984f65uJJJz4rPRecGu9hBYARj88O1iMXA47u2RYh9s2h
sq3xzxiOPwW+Ny6mtm8BB8RQLwoE4j2mmejxbJy8BuQs6LKUvFKApF/dtzZEH1iJq4OczR8vbJnu
NRx7xhm6w9s4twq+G3m8MK4l1IHg8C3hreiha3qLeXnRxG8VYv4qFSiIYx8bONJsmeFnQy3UqM5G
wnTIREcIFqZyB1g0yQ1PkWd/KGWVqWsNQ0Zw+4xn4dyLn1jozc7hGXiw+uvOSG9AmUpCMn3dJvBm
vMOAhyN3mBosxxbvRK241C7aYyEI8UFIK8fmASQVZvYr/nCI9s9zHG0WLsT2WpeJt1IR7BHb70Hy
+A6vuiDHQaWZPYUdCoyJSbW0tbjwHw7UHbOvsH0g1YD345Vqi7N19QjhL4gj+gwGE/UYfIdaVKdc
RTbiNYxY+We9EDbmxcEdj2PDACl8GV6EjislxwzeNfcXVx4NeS378m8SH20Gm3qbsCDIq0T4RyMi
CtfwLiGpmUuATOoldrNDZOnGQzbp06km3fR4MFtzwqwWDqXPPtRIPWawSbVjRFBmUfyQxgC2c8qV
0Y9/gepEoomKOFyGCAqObOlPK8PrADyOn8iqGBs7YPOluzPxZ6HBf0Afm6+zn0OWVE6pzFpdsiZm
88kbZOD2DsC23g/8rQvCY0TfkWZAEQeE9vVvTauaasof25QRkwyFBoIwVWAWfH0bXpGuVv1XiWBq
+HQD3DRgkUt8/bPlcoEgqUUoCp1traDMfQu+F/Ie6LBFxebBgNn7ykVAmSN1rizU69RfS7fh69ZO
9+oTXFDbdcNVgzQZ19uSHl+EMHo22EZiQYRzLp5AL2y/UCvuSX2z+OZFymMYnIKgk8+WlRYSaJPq
qbwqEnnU+YKkGAZ1WVDxcDJwRQU5zwFs5naufVGN59yaAQJDx1mxwBUb0JNJx9qaip6g6dTYgPLy
k1/b5p4BG+DF7NWcDsT3C5AZZGJXPb0qIOUXS8KqY2fpxV2LHfgfEVZ8zqySiK7hghmMXz7jFu+F
MftmJVNCub5n/XBG1mvVJ/GlwnQXhOR4BsFCrYah/W+2Yzn/IDoOYXuFBLfkwOgYa0h5wBeFIyFO
C6d+CDD0J5+BSzEQDfocow0035JbXN9ju/J8zfGYLJlstWVE1LSGb11+LyG6V/wzfuL1nE5L+i78
NpOtQIziqmU3TRXV5VsXyj8K5LCE0YgWQ4qcPzLrw456TAZ3jUSojmzP9L4RlnOjzAruNPDJ6jku
flVKE8FatsjC0YuSbpULAELKPInfigJ8gTVjieA7qvTfxtaSA17qR9h0KMY5fQWbsKc3lNLhHB2H
SV1+ECUWXp6sU9v3dR2AtlER7p63672f+7VhiIYJuuqtMQ6dXE42MhgWEahUT+W98DH21S8FrEYz
9TjCLHeH5LwIVP3wXoKDgFbIV8tZb2TTKyX/ikhVEzlgCt69xxnxazszeuMYAobLVSfUTCQUoOg+
Crv1N+ssFoAz+FpDKSgK0vFEpqHArJGJPAxnojavhrSjSxeaWYe+AKb2JKg9bsYjghQ/0xA9gbSb
5F0nf+stVWuGu22bCNKdm5yJa2nOljNu27v0eP6usBAgz6MmTWdLqooIfLEmi/dstbiVLSf1efcS
zc8G/USZ5VmlBFvd9mQiRGaAFQxYGvET2x4zCDqnCEKgYXRYNIFOXSEtL/pKfm5Vbiz54/yIba7A
mExmUqCU/edJwxYYV97D6++w/iYrcaC7LdHtTd+Fj7guwUTkoNIkpLO6ucNBx5qMz3pNhJvP0Eog
OI/dZZELb2XcGOi7KfxT9dVIap4xfrvaqnDkdUFLcZJnNtTveCpy0+a3rVsTC0T3gBLVVNJZlDYI
ioeDLjseuw4pqffQJpug8Lvj/SiCvQE9fi+CxEZiMSuqXXOXdzOOLhPdfuhu2joFM4Ca+MotsbUi
3u68wmEgrty3ZLv1Q5vC7w1XlAqfn6yWxxXwZZlrnOT61+bv97Yd5RwDnXHJjyXzBGhvEJTx837t
hQo/NB6ZASNqstb4tHnQnYb2cH9tAzG/fb5HJiPz7hjQABjrNpDzftnbZfSjk7HmOiMpcjGtHC6o
YSgPehuG66T4u48K9eGDYVHiVB/Dmqpw+GuYpOSft6CPAJUkHfLB/prxLW5uNL5z1NG9E27Wq8YN
MbNFzwtSbbtUtwX3nZjfQfZo514LQIeJWUUI/ZfjwgRGoHE29NKCAfGnBqNpSRlTS3PDCr9k5jDL
FpAaiSiQOzjPvQWZyMeHWd10mGm8+5QyRtMbOTz2Kcfg/aStRowpLM4bRlwR38fjCTx61wH7gsKf
nd38P1R3z5jTErvR4ufJWjxC82xZKKyVEyF+B7TqCc5YLc20/cOo1Pg3czJgCutJ/heR97eb+Vlr
e7ggRVyxfW2WrE1gUpfIKu/sVMY+OHzDkP9HKrkwYL0I3ugDrcVT2o/EcBC3Ufs6tAX6FO3+ZEec
mTjScdoOPt+abC0juHd+3T+GxqeA0VbSR1eimchdkCa2yFhJ1bwLrxSb2xZQBCoon6kIBwmOB+Tc
LAoswaLeEsT72sgKOp0FjDAzNEm0XrHepVVmD/GlAoFNISYTSArDOYH1k7KVuPp9IZvFQDLCn9sr
XmKbRYSDKj0Hg7dLTitOoUEc83pCWKrdl96/3WCi8NSU97i6JvNS5IkpGZFMaAkmt5F0Jmv36lNU
MBdJbB7INyCsjcCyVTGbBn/VKesCp9M53SBm8nQ4QmDJYDbgDAnuzlK4JqRjWxT4O9v/VGxnD3oq
XIBGmN4IPF1FF/Tdywo0q6LynjMgJWpGjqH5Xw+JuwcCgsoOEF0nOj1FTBc1kqCEBMzZ16WKbVJX
QSMIEDEnNKNXnHoOcCgSg0kuNzXynyMPsf35RrT7onukHjbI+cvb3UQsPSS3Obd4Ur2f1z42mpBp
oDEMO6168/JnKPwxS5k9H7K9jCtvfRTxzMIRUqS2FIjfnCUGmBIr6L6Y6hUwXo23984jmqm/e8xd
fpm0qMkLWfbClRFkALrfvIcv0Vsdr3H2bXOWBHUnvb4u+EEzxzUG33r/Yrj49iIxrAc7iA6yQg9v
LaovTg2e1E2EH4jUTEFYfcstOgAb0NiTtbynOXN0PnQWMh/MJMi5ax4fYjHBTkIdNFoqdLyTSbGC
pxCoUsUuf31nBGZsQxiDO8O4ZkiIFGhxsQrzDqaWreQe7yDmH6zXUoyI2CNEMa9mZBjbWtPmrSkn
iZ8JHMmB80GzuUluB4r31c9vXvUEPxRCSV+WS4R2C3INTKUTW7J4R3A7CyKOntMQqgY3c7QWmOFG
R/VYHa43EAurgNgXIbobk/+wxqmRuakobMx4CrlR0GgeOFl6YY4AnnyuXJSSjMwrh5KtEGuN+d39
8RQbUw7ipyFBAgk5BH4bcjmssnJmUXaD0M2YHVn5Z8VRrhVQL4UsFGvvlJoodVN4oahsi4rHmU+D
o6/2gfRTbesh7+CAElX2wm8xPhJc2AU0s2/ZjrcgigwZ2HhTwnJbT+bUP3rivvXDspqJlJhi7bB/
J5RQ1/tbjo7ucGhE/U0GpRxoQ0ZvqBplybn2vuPHz2ohhAaTE0NJWqzP9JCOe9lfAKG+wthIuOXS
g7EzEYYCSHkn2XUznmNgbaxsyIVGAuJkLXimWEZOf5Tat3aZsVcZjm4YcfzTzvp8dKJYuPc2I72J
uxIcGOMODOTs2IwrQ340euSdAzQAa6KC5gAMeGdoU+5UqTZhmHGJ+xfRrHvD3m29rpHF+8rdptIg
O//DlYU8TEIX3QLae5ngTqQ/H0YC2HlvL7q8YuRFwqptz/WlFnppHnCjdZGlhoVMAlFtwhw7/G60
TqvZOmELii+xMMHJfXaUGj2qzL5+YFijJSao08N3CH31di56iNcnNMQNsKxDTFHI/uft43eXH5FU
2j1Y1uAx5wFnCjzCq5LSqzATrFnVgHcM0aU6GpU6ICGyVvHpUkputBYc2LWzQY7lKKdiRtxEZ2Pm
tUCJxxlgZmxONfOklbEnoBeGJvF19gsCWD3T5BeIASNoVpCp85l1Bq9LRcmmx3u5iVlRrvWfxaJo
h+TPbXX3EvBHaVb6kz9ujEFEYhg5EUgVtrOJ6qaw6TiisU3Q0VOn3//BkM81uTYEtKDVLHwsl+Fe
cG64feoisySKe1hEzA5TWAMAQ9NkH8MK/yBR3Ydf73kBhwyYcTYGsPJaWOYTJOFgNJBKs+zlo9i2
DbIW8NgsXuWauB11L/IkuAjQaTRuLpm+dsdSWLNuHr/DHxtJBujgtwRvvQtcFt4APuixTdnICYMa
uhsvvUwQO/cSvgpsBA70GO36G3hRKTF4wamP1bmbZGS237hDjoj3Qehs0Qaa6wCSD7aGZrnscbVX
Q9hL5o8Op0UeTiYGvoIFvoBeNOq7u5HmsyrqNJ4LKMyRWeIKWzcpB0aX8T7pb87yAxRkzLWUjTVH
AJEMRp2MuOJpnPhdMRjkCxZknoRx56T1MSos4AabLE4S0XXqPbrzB7RcisQhS7twR6vU+JylHr4I
RLP9nHNLc3jLFXKWT585D8aNy58NnmfNb+iXQCMXV/+89nfbS9m3kTJaWkLVMNy7DH+791LUuv0e
PTBRG6xRYPBxIdw4nO4qQN7l2XLOmr30Pexq5KAYt+VpUNgDxu8niACfkhSGEkP77PSf0NOiiTlf
KvajfwS6raeSmIcNpcNmNkmSqfoXSszwc4lr1YQbHcxkqF8+FZ3i/7CosMcaKqp3khtbEr4X0PUF
clwNobfv9dHIMe3iQqXaRm4Gv6Diti1OjOKXmbFefS2AVN7f+dJ2lFNk68TS6st199wjS/WmZ/7+
sS6YEjJi3HzNbSZaWEAJtqjFLYe9Vtkeis01rvEDN0eeKSk3y/d1t3T6EZ+U9pynbg2dWE+p1OkR
djQckboL0J5aCopU4GbthnXOTtgBtxlq6bBigpf5E3RcXv9Ny+NiBG7wD2iZ4HlUvCKiowNgQ94W
6c19MvMJ3ZE3HNpI/QePcp4gCFPzAmsdKBqeD5UFXAGr5P940fjLNzppjKBbI+EkOJAH+Icmn1PZ
1O6Ooac4fnwLweDTHxOU7elWN+R6HeQJEFNK2/a9bd/U3VTgES0FzlvH5OeY/3j71XR9Dn+XCNjE
XVDAPiEADITinorz5vWsUxhLbKw8vDGObH40ifGU1RGNEZQs6bOhJ0n1fBkbocHYEJi8yhZs0Nfa
IhHjhQ/8v5V4AbJ9OVJfHVh3mHF1Vxtv+LGJktbypYUs1s9fCoQ8+5+I3DGZ1uB9MUwyseELeUOt
m/sB585Vxn78/Zef1ud71925UbSo+2XPaPIPyuKFP4D1fM7WENRFLRROCb69qg1XmPqTYbSB7iUw
wf0A4at+Nz7gk0MCguoG0hVnbMY+Bl1SDDpcu59QZadDEN6S9GoLyBZIsrsIxcFhaZqdWR5k/j9N
1P2pes4BQNaeZH027+MGsmO1l0otcOjNbb57KcLg1/9pfFzdv1E9cgB/pdn0Tk4D4x+4mEu3wCzv
Ii0tN8c0OiBv17Kq8FpWud8JZLMVIz8o7KYYTOASfTdUACMKnIkZxI8q3CGsvuYPKSHbEUYcfPSE
uCqJLwBxpSlg+iEklDABMXrQYsP24WnlHRyp8oDm2fu6gltoSjf5oUu5K7jLKfOm/xqh4wxjptq5
jY5bYR51qR+m7CEHjrmuNGIKVOTR+odRbBcXe7D5Yl1SUJYNVMnzZPYAcUFT0/HKIvgd6HEFzUNA
0CQmiyWpfnCpAcUxYQICnqhwMrGWOEqn0Jqy3g/EzIZTh3ls86ELjSL5LrRHzjetJb9jbilQupqp
WwfYQYFev+JsZd1wsJS78wPV9iekbzh8heaMpS45q/UH4cd7Wbj0kJinss6liU64iqkDcmDqcpjI
b7swzbZ9w72M/xx39TvZNGuJ0ltP1KwL++ilxASu4J8Dkb66iPfTtwRJ6/UIqrONxopecoUUZpQW
DGpo7O9sxzB5KHopdXY7XQCTkmCjtnqt37vzBeGMawmNxg0U6mtLOFfXN0PmmTfwIl9FlL6e1rlH
KxuHh1NYWawbe5VYylpihc6z0KqO85/FbDXhZGtKWmqG/dGJGNK14ZtcCx1WvRD6w0cUY3TAs2Kz
meYqSNizijo0LZccAG1Q4hQuKVB3sWdhcz5TIduiTXGijBC05o2jDuc9ibGkL4B0e7t2s2CaVVRB
bau1nXbB3gLOCfT/d6FslTFPRh21BNqcPaoI5sI78QL2lrjM96oZDsd6W8KuToUZDntfCEHX1G9s
sJDJFICKb75ThNpkSTfUufuu0k40FPmLFt5mLhiWEg1P6QhbivszBzAzcRY6TX/vR9KH59Db3nWF
BBWz3YeJ7OTOvDslQNN872v+ArWpVGOwo0Jtt20zHMMIvbKZK332giQqJrpOMmitPX6ymDVnovkl
IGPy88AWi3aHIBZ1GNA0BqT2ymIE/8oeylz8JZdSSPfDeb9oayrlxMARyiApI5mjXfbUa3F7gpnN
Fh5NaZpxOtnF7t96QatU8YtdviilDtMMEkb985AXjThOzrqdJ4xX475CUQ1ofoiXXT7i+SLyzReF
PfFc8vOImaqTGyGLzxK5U9voc7RsTA+v7NC7GcH5rbewt+LHoqX4X4oafZ0yYd9yM9z19I3L0UTE
PksIvv/LDUbbEVaCJKpH2+DRQZv6G+4iwKt8UQsm3RDlEkyHn8D96gqFxxBqAP4T1YDrSfg5MlOo
CwH4bsLBKIHwIPTtjljvM587WPPsI5yXfy5eS0DOosR3w+2ZF18hI2mTH/6dv+Q/9xg64+jY1ut4
UEfphoKk9+xfTxU7rMxID2RO6YvDXuIygpQHdV2h/HYqKoseqypV5mhVJofyW2L2CgI8nO6vHL+Z
TyK/vz95XsTPixrhCSYmEx3CFB9BpDZ2cqxIJHWsNMdQ7Bpohs1a69khAj1zNGs1kfmmoEmNpbXh
2zlMQjp0bZXk91INh7N33o70PThE6sJ6IZKmAKMJWahtD3DrLdHi4ZjnYrCdC12/t1Wt3LGHSNs7
/OXRVAKVwTfb5HVfmkz3rFktdkSbzAWzY1jZ+SgzVVGeGsr/SGW+ahOpiMqa/xWZjyMhv7fTxPs1
3tHw+Xzzjb1GYLvIDiaU51yLBxjn2rOv7VcD8bep/ywzqSWygLAk4m5QvxFlxQ4qRUMsm577WEWv
Zd5NB+QBcocHt/jBDmwPySQ+TPEPfCTzZdcNUH5WK5WlcCJ6qbzwN5ml6hPqCsRVe7jonTYLkkPv
UW7dYq7nlk9PZv8c1d43aB5aOjk/GaQNTBE+PCb/yEY+YR0//Mq6EtdAa8O6o3ukAf1nYLDEkw0s
ByOS09xWXurgVxKk6MZU0rmlAg412pL+VNJkekDi9zrQQjlN9OE/nynwjK+4ePJwOKEc0JP8iuZb
NtDf9kvIjf1LRHpE/K8VtTJX8xv5Vb6X8J8Bzp//H7nFc3wT8INXhNQiUsgySUgz2q8fcykbqpIA
g3/Go3icPSCvP7KESOqSA5Gmk5BV9/NubOuC9pB8ExHwbVP2scVBb4We8BxOTK9ZxFLVoBwIMCl+
don4VF2ux3wIBm+9ufTYlNSxqZiuFfkFg09Jlm8Xz2XLokuk58TmLCJ0g4wPNyVKOD0PC1fU09My
+ngBsJMvfyFKeMaviuUXAn+FJKelFa9+5iWNnzWi5PP57EIb43uvC57OMdLy1d7q8wqM+jVz04vu
2ehGtWgCPh9fkqloWYjjSpkKmCheaBOUlFALHi2dYXBzBHdliFM79FPmEhf7AH8Q3T/r4Ot9ic9y
3zhwhgs3P2Hk2CkBfOw7uJrGLtt5LwOXr8GQJhQ/W4pAgaEKixmn5TBhNPpHTEbGb+YH2PwdBJ6W
BV/IhzvDwozQafzGHaVIjZK5KGll/krj6FcrakdB1vSXCZquyxhE7t84zCUBdyiwQ3bHWCV1cavO
p0lIWYs97bukE6pJqwWCBoqk1Y06Pt3rjg1WO/pwG6L68FmB0ROhs9pXRP7+3pZePedOnxkID0ZW
QOKSrFR/TTTXNijS9GPJTSufFFMQuQSoysjzBmVMfQk5MlSAVGKbHMnwb2m1WhbfWwo+uc6r4j2e
w6eDZiRmctrfYP41SPhUcFvSGC9+Jich2Lo3TsdOuJHUmQsc02XwVbBR1DrJYcxtqc3/EJhDY3s9
BVv78mzy8vJKppLmdG1rrDqj6hSdO4O7QpX4Z51VnHpoq1HC4oMuA6IdO6yK1NN72/tekacf7FaC
f2lvcptX/BubPF6Vf62As2RmSfSSoM3CiGwTSZuekqKWHNPOLHyD6XzsSPUu0vhus19m7zUwua+q
LvXy06MbzcVHrqS6J+7xGo0sR7TOP0hdZeFrGoSW8kUlaV9lri625C/EYTptACb45EMKWrsi9mhF
MAvrF4yLvKM5FTmbXxkallRkzNsSyNYQAfLynwfXW0kyEpL/2cxw+5kZh1yH+PaQBe2UvtZTcS5x
Ou8gQ130OwQwUrsYGExCFaxo/TmSqzTEoeH9KhVJxGxeOpLZZKh8l3DS8kaN+PpfT+Xhnn1m9RmT
EejJah9p4/QiGJ7Q6q5iagqBayet6jds9BWKL1ws4FQ0+pDCLAIF5yeCVfe8C2WglpP2rox1jpGn
hewGHp7YOFN87TfT9tJcpJhpJwpkB1+FMOZMETe5yjiZP4daFwB4Ba1vZBRnJpT3obj7CPV2+Tay
TsR0Rey4/hSYpv3jWHGR3xQQmjBIr0Wmjk1w6K6S6Dg3gKBJpUg6R5dyrluGCgT7wJac7bnWAwWM
iKBfoCYsK65JT1eP8gv5ohLi+M7sRNdfNWbx7k+LxFejNKarKUb+zQZLjAP5l8I+9yhWUmboeNaF
tKpwriT53tx6osQC6zkXDdjcChTM06gKnri1N9m+IY6NAGtA55R1JRsOtg9gnXu1k3HixG3SieVX
ugLoEaT4aEsuMwf4aZgrZGlPxym/XclKhiKG/NENLH9CJyFS9+49+K2hsngpJ7dbcKlIVY4gttcY
JXOvPTb3D6ZkyGa/G9M5m5uTh64iuelkPEAJKS4HK+2vz4UzwGypQ+tKYC0OwfN9zAiN6XWfd8Mb
Q/P10IsaYXGhb/ZdbVqWSekp5E94cFNhvB0/nhC+UoIWbA2TyGd0+aZdzwa+vFkYVJfM2oX56J/C
gNVru/AYCiSRi4gqwWEctDzxIRGLxqkC6vSUvAmEtGALLm2tliIeixz23E7y3Q2u/IcTvuGBOy+5
hZbZGk9CbGQVyfQ5Jk1/Br0pQ2y01uj8WnolM2xcb0QO5G8p9GblTAeinCmukBs3OVRPX9jF4B+J
1AUQsqc+E+AnhHTpsoEpGNDX3TpiCjdL+wNjCjKi15QKyh8Wj5Djm9Ehr5HpRTfpvu2fekT/9272
vj7gNKJ3WIqw9dE/fGAbK4zp+mYrDNkcbcT+Gv00ysMCE6bYNf/iZGsi/bhys/4pv1rJlZkF176c
5lOeiPo/80V8Xanw075iHw6X1fhOxHXLP7VIsWy/djGoJUyyYVNv1ykE7IeYgx6YH1+rodmndOFP
8YoYjuoGtKn2mYS6SbZPWQJHL8ROwwizCDfPZC0t7ZFimxspzmnsthtftUmrLHW7vr/i7hOk4uWZ
1Rt/RL6tAR6SAKraP7HMOaHKUbCShzTmYVG+/h0SES9twrldxdNxK7nwZ+xhYDc10GDnatXun2NJ
pzPEId9FsJL/0DfNZyHdqO62PU/t0v/HLIP63sQbhUVegZYGwOlBc3XO5yG8FEdxTi96DPqkJJ1K
QNuR6P1utc5r/GaaEABE1Cg80SfpIBgVSBBIwxXdEdZVE3Ynkw1QtFgP6KhjBiKyWTTL31Ap1lN5
YqL/Ug6zAEAzeSw8T/Nt2KdulJX2Fu5DNwi3Lw65aeQhaDY6OuLxle5P88cSpBo3bgyrMdl7xm1+
e3uUXiJeYVnWx69LUbY+bHt++TRSUVTQs+zREaP94iILi6rS43yIRWCyVS7a/MyCteQcxcsEWoBb
DKmWRqMkbx2xiGfAbZt2OzCyba8KBWz/ahlo+FHQMYB11cdou8JFJPYzM64zcLHAcl29M7hg+C8D
rFTTN8i0ze9QckEr0rrtJtuCKxAfkPHHYk87buGPLHcTpKPrEnGOPLEG8UtkDYnTpQaVMcjZYe0S
1y587q19wDVZFIERdT0PGEU29hxn8c0Hkt9bHyKuxNMKBMxq9crQa4gX7Mafyvz3EVwK9xnW9ZEH
2EQe/a6BRNVmbpqHzZ093Nn02RpK1e/rSQj6wDcoe5LssFeUqLiS+YAm+TEzAItwN370ISmxj16v
idJvODTcyy/uiBc6yio4tSW4NI3JDJv2PxMM/UofPTB9GB2X3EsWiPjUq7Fg8ykRch94gDqM5ccj
+W9IJ7lgkcPAVxFpMfpolKjrgjGy03wdbmbAF3uHKLLpc3OgtnSwVYyQvXUM3ejJeeRinYgSkE+h
aN44O0Cog227Uv7NtSeyIob1RHAc6AsIQfqDSt2A/Pl+jYLfCSyj5yc8aNR8SZA1H67BG1MfGzyY
CP8vtq/Of67jXS+bM6gAUztWrff34AKMB6BWBc4LX8W4atxLNxy7dNhOFK7qu+3sRzEvL08gvygE
IHf2mUxZLtP66yq/2K2wfMc2kWj1JTCSgABCYpjgiI8dAX2SQQuf85gjHlWKABse6vz3KLMdv9sm
xhETid7JQWgNUcynjzEZCGZupveem/ZwlNARDqjGPch67vTGHGgl5dTdKXQLZwwZJRvSx2Ms6tjW
/ino81AvPtrmVxrE32fZSY4PFssQ/wqmZ1to+ZT5fRwkRDuxdcX662r2YRNUW9DTz1S7o9kI+vrE
k4RGmq0phEP4tV00dZ6n/lOyo1PMeI03Tzt/R5RcW1OXKKzVs8biU/WzAtTf03naKMShFUWo8oGV
Iy2kY8aIqH+E8+XGvzlPFedrUCvV3DJ6LcseAw8E2n/f77ltFlhrNJUbaOoy0INHtizc1AAXv0JY
pESQfbfA9aDodXtaYMZqzLptW9bKWUqqWNUz5wHefFPrxX1I+GTJSeiMjhKyvDPi8zA92qIpjl5z
uHF8gHELE9blvgrYS1fYK/Ie+kfblrhy1OCaEhxtJSx0s8D0INW9rbnivRLRVtIEhBO2zsQGxv19
RI+L8FuFhPpfa+Qzn+tx8dIi9oUR60yGo369qn6UV+MvwnysowfXdeZn0tBohD99ZppV3vAhAXu2
24UypvRyPRAcf3Ji+hm1ZRnbOghNAAe112nxu39gvmaH5m1hINauZkFUPbdG9RS1eSrhsw0CXLTz
nq6vUlR/cj8zp6krXdCXQRoYQ0Eh1fLJYTChitgNcS3PsWc6U3NQhN5nRXgSSXnMtW6NCkaYOVRv
Wa77B/Jp3YTfkQNVsNJ7+5xag0dNcfgGywil85A7yPf6NLgniQg1Quod62IIegUTwd4S22v7nr98
sOcpCVKxKxKHW+VsJHnJwf2yW2yDn/KI2J3ugoDBPls7vI/tyKA+9EyXSlhUHTQ+fi8eqrRj2uiX
QwtRpvuO8TzsHCOzSp4bK77QYkaz4LdAGlh77x5VWT4qXELAmRAExrHJXXxtvv+doCUawq087tLK
bj542cTyO1RfgeDqGi4xU6iLLkEndopMNf67FmC71UG2NKLrkJXCprVd36NdBkZMGeXI+Kp2e+9Y
6htnA9P+0pDB2JsvKifYiNDp6FIy1E8lreZr6h6hKQ9g1YsxIm2urayAmM/6DcULKATSp1q1hF69
v5wRCqprx+IF6ZQUH4tAloW5e/e8oU7u41+p+zB7SgyNIjvu28mpFelxMZn8irBUp2FybzMz7F2k
A+tbnQ54UorxMi3WWODdHN/bKFcERsdN+nyuXqQbwzTgNpD7BrlbhgKo/7WyPAUXmfZu1tPd8Gsk
qL8Jnz1pm9MGiSWjxqUkzWi3fn3pzHuyz8Rh8PIiv82G89bC1oISwbX90cvISMU0zkAnSyTuJ1Mg
wpfJ/nLnXTSwUqiyZTexbBdwzyPW6ouxP0f4SuSKbLcJLa8tsKuEJXeY2bG2/iUa0FxXTA/JrD2o
ocZSkT20m+ogf5qUYSBZQsn8CkHP1Z5WyxatlZLSLLX8iZI5NSr8lAtlc6mG5Lo9/SniifgiQMC9
FBm2Y1FSBb813l7huYKSkMs9qr32HLhyI/TrdQbyKqY7xOS3kbvzlImtDNwIRYgG8Go72Plsm2Gw
ctx7atIQhVUVus58g59FXD5s+PgF4qJ9LUHauf1mrNVjsFqXCk0d2qtfyusgdW+b+ekOgOo63Mpe
ZDcXdgPngBwJ0R45HAW4S/qSUzmvelAvCEKkpi5Jhp1npHBClt3bOAon7D1lzgTFltN3nTOxLnYl
IA2v+7ecNUchK5dBfRsAK1zq7HODXmuEsL5nKawevTVnVcNsPGA/DfPcBkFoSib0Xx23Th3gpz2S
NANxh51GuztvsJvdsvxfyjPx1gbAqb7lATSCsqYa27t2NZp6fxfN7W3aAXdqDfxapYG4htmJ7x0u
3zJGrvxy8gykzSUAOXg2IfTmgAHrYNawH+5KdhqMquvuYikIg8o6TF3bScRVeysdzBVNSuzFaTAw
QiwS9bdej34TMZHU6VG45d720sgNX5arlRquGeRnExoqEwpP5yzTsVnfzR3D4wThCqrSwVJRoVAT
sXbAc5NsXQ9ed9xmRb8QMZVWRYH7jBLCgGK2gfgjBvzXyZohQXc8DSLBvLajP5/1A1dXgV8vpOlR
bkOQDNtkDP7poWuzqMTdbYIdz8SBdeSyzzp7K+gGgrvNGD37xA6xvvnaKolU6e3eBR64IDN75gv+
4xNkBRgb5cy754j4qxGMiRnyoIDbG23J4/rAplee0TKa07EW62WWEj1XWDgIwRD2pWT3cGqaBtjj
Hk30MjDmbwH5HaQudHlAH8RwokDYv16lsIBy8mfIOespUXQo3Jkq6nQyjGGDYduVE9GmccWgHDSn
zEerP4/4gdCLi6m6yA55QjI5uuBOkMC0B1Hm4G/nTX6N71tKSiDeePEZIh0s67J3DRAG1uY8gy6P
W7xb14zzBedrAxR85mLejKZEjgHj/EVPOqzTiYHH3djXKYnPCLMcmHS+/Q42YPCzAaia4Q6FMFes
dkF9HE9gk3Wz7PAWlkbzMEvTUxPgNyopCrxeHh40MOSv+rEBsO6TCFfLcDbwXphipD3Ch24o1WVA
RVwGYEivPi2Q7eSPhJJFmmIwyIWlYx4RQsqZpT1PsO6dUJlh0R0kehf1PUJUw0XDyWdd9C+ZwTre
zwZIkgJulsDjQysZhd7GymskJpmZ4Kez/hzko8cgR+RWeMC3XYj37Azo3+uDxPJTr7Joy0jSo5FT
LIsPxapXkaQmT36h3y0IFlZ2FVSvKJdKKE/KcCSU1L0ntyN6VyH6ECYRPgoCiNwS4/kKPob7R/g3
YZBtTWxG0aDthE/usi09Xbgt/INRrzcoT/Q6W5TFg0Jygc3ZT0mt7aJFKW6fj9DkBoeP7A6DVEDy
3r/mRV/N+kAvw5Q82Lxm6VGzHNIOSp8+9C1LLWFSOzazKlK2Kkhu7T/Eelrw3xXxnaVDNkuwGuyk
uJX5M4NxJftXD7Etgub1XePHNLVbYCH30pJjR6bY/pKGivaNydarqYIoXBGyuiHOjz/+xrEBoQhb
4T8zJM8nxumDysXl7Nlz1ofgv7OwHIULz5lJTar0rCNPzbFZZTaMij6PXs1GNwGfBnsXH+6zaV4g
5qQh4lSX0OFi0+q7uoRQKlPno2dfEGdq/kGOGy80jU00gKrbnHawUfpOEBebddEHibP/dPjGOfuB
XDffM6/IsAjcjcExlOjoCGs1Zur5w0UUGpGdc7cLrAL6WFPIhBSm0rCk47LUdamAkZtSOWP+F7sB
r6LRXwvvl0CUau6jGOTVngzIjPzhkMgQ8L2cPEvDA3b071N7H7uJLuOPo+krykBn5plmQsrD+aAv
+vCpEEZ7eQ8gQYLziVG/OXvEgzR4xBeLp2Z64lSQXSyMsuQl4BD1kcDMU5ww9VMZ9jQDq9lxr/a6
p0NZ7DjBL8Jb0IMUn99pGEafJtEezdztAzG6tiRigYpam2Z9oRo/1cR5iK/13Crm9bDKUNC57L8m
SkcOXpe4HT0UI5kSrtWTK5YBLdq5PO5iGZ+oBeg4RHURPiSxJiaflTLCWTtnIEI90ZKX2C/mml3U
5if2RguiXblxgtamRCZmFqXrZ24JD0MGVKz/Qrb8UuQWVG5ORO4bnMYwpEuB/O/bNN6hlMUfdAJC
7hjrkkMYT29nSABGyG22UDfFxUHEDybqCJzAlHmnyzv80ZbOn1HQTPnuNyywzJ3I9vEfCMYb+rvB
kiLoKjY9W7eN0CHDyVJkxg5U5CsqI5Iy0VTdffZc4WvqCgyvED2fU8OKycPwyTAhfnzsOu4/33bE
jHGhXB+KN1Jnoyy9Ka8X7T0isHGYL6syfLOmwfi2V+IABKGwB+iCt86NjlxiMptQMBmLuVQqfyLj
6Mu5qZNQ0HhDGjDwb8mRiuXj8nk8+M35GBc4HMdrMQa99qoM9Syf7T8qQEd+NIBNXb7TYDWvGk0r
dZyfXNR3VIo1tWpNn0Ax4+m21UVX7WTHkIPCMr3oR6wRbnWGjp2TQAZDEtK0T7kF6m+aPvOL5755
DWW4U/vxSj0qDk2V2cP7hXoqHwzX32MhpaSmwrbi2tS31xnPUFHL9F9/G5iRcVfpGkOGKHQnvgA1
uKZ7btKi3JRrVu4zfdvi5XM3M2AeMGI+gIwnwzuwQGJg5oZYiUEjDXde8gAEK9b4u+zZ8ugDkML4
LjZHll98UOHjFI9gBsrgtz0Pu9mRpsiBuT15QVn3RJYI2wA/1h7cs7+m0FRs/WDsn+ocqdZj7Au6
JyhD5PPdVw9+Cj2WvlfcWdR7XaTP72WcILr8h4z82ts3ldwyA3hm79hiIUy+ZrfW0X2B7JOFR2BL
WpLuJ65ubF7UB7nllWFkmjuSRSRKrw0wzwvu5rY9urjOq1XGeH9keUrfRsaLNT8vaNzFdNkMbbVK
tx6lXFCg+Ok31MOUWeQg/nIemijLcaMJBWwqidaMDGJJU/lsSshYWUcSwaJV2M9XgKqLUSuieMqd
e3Zge9ZVqc3xifuiTOBpZMiJULzoQe0p75JEcRnGqFqmHCT/KSCZhzNOJM6oQ9UimAcRM3F5mX0I
9HMFtIt3ARKvw6IPvXpyeBhAOS00LuZC7bstDxbJlZLoD3Pphp+JZxdeg8hZklmhVfnQ3nzBBXqP
lqKwhaUNnPKULpFPIkOgnMJsM7/OAIGbKjeq8mNVk2woqsTMLr+pFPq2+tR6i1Gavlrq3WBWtd0u
Lj3PvhwGMfsFPb1ah5jV/RlGMJFWiHRI312b9kC2YkR73x+DLf4BOsUAfOzmRIPCn4q6D8HDkPIh
GqVmuiqLAeQOiAkBHv/ZBNe0TOwQu922B+/qmN4gW4d6kRcz4lk0iV3wiAHwsB8CXQZn7f9kHGIm
HK0q8eJm+BkOSjg0Y09CKJrwPWawNT1zjxQq0btZapu1AjeFqN73y/rnUiK2nprTZiQUSgYEmXbA
gEtYpAoB9b82UockUVk1UDLRrlnUYNbg1aoHKnb77Zx9k+RtT5YLuEAzlbNW+oB6E6aZgxU3nxys
sXmUhY+y0hAwpe/XHiYHN1+PkuOMdpcWMG69hY9ORho7ywLQ5WVkuA21EZu/tUZ+8tTfgXz5ZBvG
272xkHBK4rJ75KES2+944Sqf3ZNOkR9euPNAlTKO0ErEGe3KIx+rEI2T4oDL5Aa/sqmnolQU2bzU
LR3P5rvxU2A11EFyo7EDrGrR9gLMGx41uMEaZaciaHkvBYSt/hKXQqC0DGl9kFbJOBuIkTFSgNBz
ys7hvrDSzFP2q4yOD3kMPn4tGYlCi1VHAKDlJ93gJGrgP/wwAJRgscnA86pC/iZRk8qBIRoIOiHV
xsJvvzpVbgIBEuAhkH4YwV8OhtpL0zUJRl+yKUfOg96Hb9/3tMCNDLkvc4JP2TwCYp2FcIliqTVN
hMBmZze7JZyNMFeu0iLpl46bCYgZO3wKuzNFayNme7UKV7djFFxgc/sDaQJI5nR9Y6JEHp0mrp4i
/n1oZGkAD315EjmvXcokey1YwHgWUsJVmUugDBnbMVdjWMK0iluxCHa4Jia0ce6GT4yj/tHh/4R8
LW59rwMC87DtDqqAhcxRyvUatKfznL8AwA9oqVC1BZ3voIi7fc/3omHiw4P/4xkGrM1SSlRB/l76
LlW7/Xot295nQ6LK42txnT6KCi5YGqr4uQhyoy9sQrRNHmL2g8SBI3xMQ0HsiG25avuzDiGdaRJD
54QB0p3LJqgtbfuGLjJC+qRJ+muJsQLY2KqTrtRycHoDH7ghYUKg9TEfBNaMT4cekMEGntke8fFw
vcbl9iyafmJDjiuhYppRElBUCArZBGzL2aOv5/nNMJyLWETQ+2lkjASAsms4F1JziLV6X5oT0HWR
Tm/un+9tQmCENzgj+Xif0bo3vnqBaL0Hor0sKQBiHFdzQ9nox5l0N243hLZyUONnz84uvt/B2I/U
bIiCPndPP8dFkIgI632NTmazg4F+oxw55y0sFizgYbNswCg18DTXU55Qbe5DoKvaqKdmLYMt+WPN
XeP8SnIGiAyLURPYUWrla1aJHgBFo2EV4CO2SEjphyx0xGKxj1ZtsMRwlDYSbAU9UHmgx8Yh6VOe
u4TS02vjWhWW3nAflav8dPj2yIFV2cKmPNaVGROJ1TsD9UzterYsVZz4sBYk+HimDpXmLmIwmx6y
mQDYF9M0Fn4kWI6EJ9x1xQ+vrx+zVUYnCSDnaMTUVgy0K2tbXgEUAHZQv77hXHpAvVlvA+n2CPUV
tbgB+d6by+H5j8isBFPIA1eeMhnChsQEbuAKOboCk+GWxW4QEVP00J2vanR6HBf6CqBtLQkQr3YM
Z1pCgmFhTtvHnkuL18PPQHU396VVMD/w8A3AWS/qpV5Oyqxvj+HA7b9kb/fYcUzo4J38E71pxcdO
2iOe1bHyuZpQwClaZr/xxjIa0k36+y5yejbbXC1CcqOoDVvOwF84GbtlyTbIrwNdQJCI2XFuYPlS
Z17zLIMf+DFAa6+HkrgfkvlMfMU/yyuoIK/IkVhTc0opxI+6AUdkIWA92W6wIf66yP0HgTxRujE1
Jwe7kTwV60KpUvRrFjGTPCV//ZcsyBdAMTQ0h5fhAW39bdjHgDxAR0uX0Y9sE+cfsNFFMDE25aI5
vySB4feG7xXvgVV7qTcc2ClNvzcyNogkn1KcEYWdaLHfgQIFsfeO8mrn4Ja/frpGq6FXnxgv9y01
BVz2i5kvQC+dn36w/Ab21Ny33zchA5/KgrH97f8w0GsRiCJPS7C+c274zdFQt99V//5Y56rPKsOv
ip5Yr0cZw45pRPPxPt1XRYXMk5x6uTaW27Ug52Y1w+nFDCeOIfD3Zv5MjenuG5oQWYobuVzL6EVs
1VmwDY8o6KlwCNCRwo1zjOWkonHsoXx3DsU13BTqlWIDbWqY719O4H8sCtb0iDkNh1P6MndU6CcY
yRXsWk0ZrTfkWVhGPJkjq7jCcHbGHbyyJF7mYBhPih7BUhbjwUyJj5nkVpFIdrwjKgH/tvMk9qNw
BCS4wKyJxNFFZXP2R1JvRIZsiSyuPC/LGlxSCpreeix0PFEi+ssRoApxD+GcIBDjV2GW5NRYL49p
cJa9J1yhyO4c2WuEN7fAKgegoZnm2jMQ026nYh+QHWy6V/X9l0mPfiVwXcN37XrEo1ry9ZO0XB3z
bdVB30QkRbydexuIceKro20Jg4BPQINvZG4ifNvKvHM4F8yJ9V2Aa7nULN/8Z7JUJF6Mu+FVnt6w
heXS/9f7cGM+G+5tRXci9SO/b8rNumL2PRHjnU9CNqK+8/qrSiIIhzEwNAehXcL+DjgtbIMf529C
lRkWTbV9xjbgPP1l3sA9vDqxRhuwTie5PQHDndKA7ln9HFW4jRf6ffHjThwT8qRZVhkPtzD0gXAi
a3YjxYxvdwM3spk27QiqbYZ+F2lcNkUs8CDOad3W5TGklR3/ezD49bnw3JWJU8FwqvJ+cvWYqzWM
IdGkc7pVUKX+A1E200xQpybUSF+ZvOPQ7aoNNGJ2fnIpia5mK3W9287rBz9K5tO4W8QQ8jGUTCHO
wy6yFM7vjOpy/ePhING+pR+0HtZOyW1R3mdqg2wAwehj9dXYf8HzfPd9qsYE50w0Td3AHtAcO3fo
g8LaJg3X/luI/e0HEYqdJHqaRflif8O9ZbRtj4V7GRuL4Jv4xpgFAdxjY9Jo30DNBtLXW7cJj8t0
cwlEmI+1GZJum1nMtZVDjlG7GDysNi2GM3mxNxAiE6EGTVHZG9v9Ew2usNbmmRp9ZQvS2Hg6+5VK
1QYy2+aG/yQx7YM9E5qha5TizqlwOi2ijSrGirn+ColZreXxVDtfLkqnxu3SYyqtAMg0mMpFNuN5
9FQxCKb8wl/O1xFwK0UCtLPIMv+LDhz9tO5XepbupVxQ4iLLXpjCuDRqN8l8mKWWtnBwZfP0s7vf
zgnCGrLFCkNHPFCkIBvTgVJpT+MNv97+SeVjUDpYWnSIM0qbLPc22s/0f/KULc8Os/LREbBPWKU5
IOdbehzvFLSD0cnT2sW2MjeTg7aZKi7SGI9TB7lvMFJsNmOc4hq4i5QRZTQZo/78OXPWkELvQ45u
DelRB7wAB8FNKw7fq0n9o5Us/6czxyXkSXamu1L3/UmwFDGOtVthe5oZZX0DE6Na3boyPPFRlUde
VzEWQyy9WoYL9G1lpWU3EUs3sTbi9bDrX+ITXfLZMaa72jRoCf0xYfOKqGQwv5G9MgRqfYW+hDpM
xKbox8jNHSTqoKZZvUeazbqwzfnbeuGzsQP1jJMrP37nUUUmvK/NAYsfZH8Z8oBCwQ3CD3Vl9omw
cvD9xPT0KMqAGA7rGKHY0bwl2roPuIhFKYE8Cp3glVmRl10z/gQ5udLdKuYxIiUpDhx70SKuw/y1
dHJXEIxizvovgSwfMuECu8Kd0cnHBjXxbf0nKulY9q6F+4jVrQlWhNR8MrA1Ll5ntP4eUqwEuOIL
zaIeg/nsLlTXX02JUmLefzZQ1G+b1jxc9n500dhj8ThDFaA98JyD0zmHFRwTCJLcXT+ShexGQhXC
95EdkQP8WvdiMkx0TJVCPH54GiNQlwJzsRxM8qoTvdmmoZYxF5BYqHLdOKFPTAgA6iHcvPkEdZaH
8h9TO6iI7RWQXkT47mgnkik8s+9CS5nVISZz6QTFmkxacqm5vjusZZzDt9Cp7hJOFFXMBWRjftZ1
2wka/SVeNgq6K//dKRK1fD3mwEkWNdeFdH/1z/YP3VBnGRpzYy6ewTH523U1NhWDNKo+DVmXTos1
0XTsJ2olxd52qyhXSwhLMYDU6J/n6A2DpbQr+QCgGMszve7xv/b5n9RqaLAI63IaA2ByD+QEAfIL
neshB1QGMMRZO0Pm9Ssvb7lEvtV35CZjDDN0X7XZ/q5dsFDrA6AXrdvRYO72NJJobTjc/7SjRSOY
lx8CQGfE5rBuURf7mazMGHozxZmBS9yhJGAx/73KuTi/AIC16XJryAw4JDZep2VkNQMBk/Qd6aED
nHEO5icIjFDQHZ46w5dOIT4pZQv3f9WqI70c6KluX2v7+Ed2WnAE4pydxKxqoTc5G/16DYr9zDOn
IMp0WeWePYT42drN/ox1iymSEZ2JFEj7pmMtHrgNd5cOs3Xbuy/+VB4CTBy5NxsxfGGDz7Op9YRb
kszMa22+uCVz4tAumk0Thj0+a9XlOAtYyOFWI8TrTN8ZvdKVF/TlITQ6ZNlv/u7kwhve7LjA2veL
8if3gOWIpnAyqkZPAknt9sWBuHKDA+X6ah1DnNTte2oShs8hIHErKEh4UP4c+0t3RbbuXGUT3r3x
W1bBz5Kj1Zkkkxl+iq5LwGAWl0z2RfmpRxk9Sv+kw73VkF6fV2h0uUuFymwhS5s949P+sEsclqHm
vL1iR+lLt95P8OXXT33nMJSgz/FVPnMVs5BajgcT6v2Eh/+/VyNB28Xs4UtWwJ9n6VBkbjtyATYt
250120jHHKchRwczPDwCDwgB3LcscNduuEA2BZI/Su/Qk7nsmEqujKMocFC7hPLVB7E67FNtVsz2
zfLnc7ZavJWMwQImEqw8bU5IJ7nLB4l/QkP5bk8JH/PNMQ25u+vseJ02bU7RMpykJRyWnXGau/dV
5pK4oMVu9zQLmzB3LR6WlAx26uuIMp7hTkLqiJggetnN9Q4IzZNrsBV+aiLblurNifR+Ct/A2VDE
2uKVSruVZBKa2JhPz6lNK+rzxGuODOZW02cej3Zt34K+Sn1+gbxMGiIXNeLRk0Xaj1Uq8ck/0BkO
C2BVLQ8K7j/GaywXPM9XeLG+0XMjrTIvL5iYsHF7Yiie3o5Adh7pWIKj8mnCBtfUDw0w1nN8Jpc3
voj8mTsrycaKraWTMrvaxEx4D1ccqC9YITIYYy34GZmZWsJLVkFoddCsZBIMYh4EBmGVcP8co/JI
q+q/uDxsfJXgmfFzVYdBEHa2z3AKZpO8JXO5LKxuWfa62Nehxa5KC2Go93yd3fNtbpmQpTyeRruk
dOilX4Pvlx649EZC72ioSBaCtGJIkrurPfnaPGHeDkZCq6ctMCTRO1RfIwzeuJWJTKAInCYpJVfq
1ywqsqq6JhbmWZZK2aBmS7TWmZAFCmZJ1uZmmwQF9IrrRPQ3xGMQjcbCrO09Qp1F9+H74fMiJcGC
cVp6430zFZ8NzT+WtysKWEFjUprynhO+a1HZk+uCaXNy6N1ErtqZyVt0wF6+Csl59T6k+BQwAIpZ
wHWdpEZEmkSErOMQSfDH5KxVXNHWABOUPoHWbpksNCsGBMyoRtxROVqxt+EHBqkYtwgR2ubTpoUK
Ke+35k9oEeioa/MydonR2HAPm6MzMj0Psp1FClJsGaP2x9zQkU8uCDfuvsl6sdWyStQGkQTczo62
8NHYootBdMxp7VL+qkZ8SOUICUnQspYNVAhEqGsGjiRyjmdtb9GoMWWq6VdfPtwBGkbkTXVI/wg+
+0vF70qLymcZV28pffhv0Eulfrp7hnNj66vHndaqUXpLCEknktcsWEznR7Fy0GLB4OqnOJ6cHk/7
TZ21seC2yZ1ZGGYgiU4JRwLcTB/amz24TDzL/SIDlurgcvMVMqBuxEX4iPca8HtMQtTFzgbLmzhw
wT/lCDwNRyryZTI4nBe68RjL+YOy85G35SM6N9WLd+NiZP+N+hV47O0c9UYXy3pcfHVNo8XBrLQk
THGTvNlIV3tw3phRLyRIUb2EeK4HgC8t6qxVnjdpqfat3OQACGk50lONxHC6N8s2M/ZM7XiWeQJf
DMO3iAVud5ko0V5bNZOZ+/lt801VIxGRJI9yknTW9ikNhy7jSM/4Y6leq+WUwzljoCGykVnWiL/I
D+BudZBXJHkyrmaazQHFWr9r9tUNZMf0suA3ILo+bQXdWaEV9L9asJrQHNdnBqwbx/pYdx6PbsSi
JFi1bQRWmhdojOkAZyv+8493TnRFlU5Gn/MdiL6EzhPuR3kfpzp5qKt1JQsmLjgc1WxOWgmmWlZ4
uPcJPkoqKK7lx6kEpBeaxDGP8cAjtLuk0v+myzRoWW08BBuH8HOpS8QDSVggr/Cxzn6tkSn5sUZ6
OjQ3aO5WnYPdFgcBVnVY6zaNWyMVh/Dnpe1J+z7yzHvqB3wqiY0A3Lk+3Z8HMIf7H39vaL0fESky
11JdXZDbdGLZG+UcI1rmu2IkuN6ca8rndqjqWujzmcUtunnM6E1T8eXNudjiU+VqU3MVhMRuza24
r/drVbxZdc34TD2h8o/9NOdxgfr927UrIDUI9l4yoFuaAbrrequ41QqsF7C5PZItWuc+XIvxjFUn
c7S9v9RQ/Qg3UEd+ewPcJnkQiXggqA9vjVuhbU7TYbvcbJV+fIRovlAadz/vEuldSJqFzBLfK2Gu
VSxR07ubeeKzqx6eO3PqLgSrf279+CrXpBoVVckE3d5Za3+Eom5RzCMKDHvwpTOTQ114dA7FOX1w
kDP0eG2QO+HK16v6V6uiJveOOMWkkrgIeobj6T2bSf/5KADwveUpHTeeRCmLxYL6BEcVrErfWcQz
D8Nwsh7UTaDXP+GoSyTtYi2tgtKXdljUGmRzDi3s/NOMvbCtJHxN/awiZH849N5bG33FHRjPeZGj
Y2tCP+I0VH09HyJRhKp5v2Y3Fn9yWcyNVfHmtIusROLnBfCqz+YYJdBo+rumPzUSI6qkJlXlvtD2
A00LxI4bEKbcmUC+5zGoDUh/U6Z+zVyLRJvC96is40ePla3xRxu3ZW0JuHrnYYQOg2YsRHtUQBZy
SwqpyV7zd+7K8Xi4d6T1yWd9ULIgtiIctczJcGaEwlby35gks3mKEcUmzwhwGRreLWWooGd+HE70
pmOwhJb/5bqWhteHEv4XnhU92Rm5qubQkj5fE7jB1/OCu7hYpArUIjL21GQ1gkB000oJnTJll55f
DbSsPuzDx+e8AlKkd9D/2o7eTP6fQgT7Q7Bc/G5m9JG8wG6RT8gU/D6EdN24BbgALoAUFn4RlG7v
smj01ec8sFfJMLJaAp9o0onJ49nM9zTtgnkneLeuqKxDgo4SiYI22gIGkfLrp6TPpPhvD2Z9IiuS
m9i0HdVoBqKZy3M+29/9SN1OaHggURD6KIVRedcMLLasxly6uSPSKGZ5/5QWyYZPgreiLcqG7tXg
ZHQTOyVChdkgGLs8N9nLW54toGFolw903lV6NucqqaM/cTv8rxloo6y9CNZnJkkNDfUWCgkFlPNa
9YOXgYKu1WYR5LTw/bP9T+10WnmhMpBHqWjPZr4Dg2q5aDeGKlRCwX2ZEhPmEuKoa0p43pTELhN9
RwfrnklrTEYUhqsniuiztxP4A/GS4g5bEbpDTmQybYDxyZIq+7f9I6KXP4sx2DG6RQrYnTcL47Aj
IZ5X+iSlOuSs+Usap0fQEAm2DtTUUIxSki+eF4v2Wvz+On+q4xpLbGqMqqe9wwkgSymSmHAjrRFZ
AQIugv1Nxmok7hV/4amtOY+p6Luxf7Jvo/6uSIQtOSay2XkCH3t35UiOO96zH7RYJh1jgQ3QddLZ
dgz62o99EwjRsAJvn3INuWhfpZfpvfaajGLVgNVpEKVUF5ydxbEV5h1BNS1aOfQ5Ekz2Tkea4xjB
4SAXrDKVMFdhWn+KToGdRy8X3D3u1ecLWe/FMuhGEh9CKBYqN3MBb89swQ9uL+pIHTl9NSNhuOhy
95ZhmlJX5j5tft3uZEuEg6F/cROzY/Z6aZnXr7u//zAKiTVzmtDHAMwhQm3Qb7xs896zA7ONWALG
edWvcYzIEIE2Z0up+txm15vfx9dceGlPQRH2BbCH0nQCtL4G3sLlnR345w31aZAt7aybedF7uS6C
KEK+gZBiDF7BouiZP51Olds740E/11dJZiBzH9n03tY7r1bHvFDYD1XjyGqdidCjiE1RqWYXoL3h
B3SnSlAX720dm4W/BPsFq208BdBcGzs2K2c3vQlcAHJMuhldt+IRbGIB00Q6ASJwNDhzVRNRUOd9
C2O8Yr+Ndf6xRXT4kVAJspikpD95frNEZrRnIUwbuxgnrEK6nrSKuBOMtdLkmm6juQ6ZV7fT9Rwn
ufatARQl2hUMYv9Ec/wjuawb+aFPvWa6oEwJXl9g1WyELN/GxvD1ZBwL/F88pTuOezI1ZcvS3YOm
Xy/ArHNNJt5Y8pGaS5iQsp552SdMCgSBVp/IB6DmsFSxBBLz0k4NU0nZLTQDD8t8FynIrPli7Sn7
anngpYv0iwwTJSCSTXm71Y+DW6aPTp0NETIy/gw0RqSfVhjQfnH8sW5PI7wXyGFox6FX1L3WLJdh
h8x1jzret1gU7pSOGrgAqQrFHf6JvLE5nmh1NIcWdgfvBrHM0uzJ3S6ltQ6QaVmgUSlDUv3b7gbe
OKQRt97czyDDAdfIsCBgrNc4fYFADIDGdLEwL2BrAEN/XmuezwmPZPS1Mk6B0MtuqEwlszgkxF+9
SNjQXsTsL+3VbBewdC/EnXB0Q3rW5HPWpMbY+2Hc6w7jOC7q38Xw8WTeTOwKsbo4QDAq/Qoqc2LJ
21ND0bc5TsUNdEZ5iGS7S1mEAaPPIyPglV+3Ay2HGvtBAqybhPy2j9EbhlHOkh86QIBzR3mjnl/p
ZDu4lrTZnLdGnAfr3Dz32X9iLp8xHFmT6i8OxE+jy2mBIoIsMCe/syL1z26Aw+hOh1FtHOWKjUcK
zAPwuWpVM1pf7YmTqTVwnDhvpm9ynTMeAkf/+YHwdMCxdIB9Pzdny+6aXRy8JPtxbaOIjgds3lKn
kDHeA9IdqZgs2Slu9uvCURHxQaaVrK3F+cipDVqQm1UBipNGqF1qDZD42Q92MpDlEuJ6PgGj/HQu
cjxbdia4PmxrWTbDQ1iehDZSjc31ERuSi426eKQADFOH1iTuTHtOc8mrx5tNCQdS/FIC/WFhZ2fx
24HmHc9E+FCGbJKIt8GDyiZMOpkqG82WIGBS0Stxxevxkx4a1nICeJZHUfGDg2k9G+k0yqMEq/tI
sy0d9xIpTwW3F6Wj3dG4/XysmXxa+9IB+JNXzL5+t6hneGVb00ZY092P3jH+xBoW0SFNtXQpYLrM
DXy2wwhqr7VZ98bybq1mXHvffJ/vRSDiv4WsMz4PMjO/JG3GFKBR6ckxHXKbXNpDIXdWhabyaf4d
c2M4xXSCWILRhVzO7u2lS+SztJUcdvX239kKjb5lc6wnD4ojWfYNDDiRusYPazNnDV5JCOk167X9
Uscao9nz71rwCciZAIq/ueH/X9/Jh6z8WSTULWta7SC0pribXwQEpd8+cb1iJLh3RWMPJ7fGTnfg
aXVwRVX8phkIGbu94HySGvdsVsAVmN0zcnnRc3GAo/ryEqqTB4H0hBYlIh9+19xr67Q3t0Poq7VZ
Jff+Rcn1VRNUhbnvMw7UaSn25rhBQ4CmC/Q8dIPI3EI1etMGEOOmImcf64P1Vr7YzZ2YhHCq79QO
BloxLvPv+oL7pDRZiS9syOQhtPgCCKMjKINNoZ0/Rwlhh6pQCHOAh90v4oPykdb4v5XmkQRi/jUT
nAUFeLxVgAauD+o0xM2RWLYnNi7lbsKS1haD3x7xIohp9XiX5qLVDwkwrTSOCR/hAYnFPSY2ydBd
Imb/hxMq77fyvCInLUgxSsuxV63R9rcVnjsb1+QkFpjQ/+43/CxvUde/254W+Y0AMlnWzw1eS7dE
pptNQ/gK9Toph1/+YIJQ3lxwOZK7swiqWzNLsw/5izIh4qUp7QoPtpLZFIYB8hd1+PYuQklv8u1J
Dlc240q3V/hY/P3lfIjgyOdi5hQRpb5TvwIYvurY06krbPNa/VG7Kri2BORkaniwSO6bFRkqTBcI
l0352zessjYr89sWtyUFbHyePaSeCGZG3fZUXLLHdp+ZSeEmK+EkwwV6Wz/dmTt+S3tR5eEqz9lL
ySaRTQp4arqsFEXT2z07nuQx8EJUArlqKzTOX0S0q/5vjWYwxYn+XH7utfGfCcA9Zhxb/sVxM4N9
QdKIqeBXnQ+qsjAmgqRDvekmGsLysxDXGHddS4TApiX0/SaUjqZJRr4LqvwmZwz8Dk37txvxGbi+
82u81kf8eV9r9Dnts/1Slt4zSnehrCnjNNQhiw+ogGDlYfWPdR2q76hQ3AUzt7QJOXBBpc3DvxBP
xw6i2/YFsmRtA4thzIfoeIovxVXLkASaF+D4VjYPhjPd0Fsap1uMDkT1Gx0BwKQhoWGzy7uI9KIl
NTZY30I1sozr+UvAm5b8QVWYCnjE6wimqTrhgzSThECFOTYzRTwg+Dc2me7x+D+FlrX6yaYb+Gp1
2RlkaeYlS/UK1Fmeio2lw9vym28v4FF6QydUk43GvnRA08sDHslWq1wwJSmqR1EglpmkxUiSD4lj
Jj7RWE3FbJDFLaWUpmnZEYAN4LEcjTx422yJWaIyhXRSGRaIhSgBmgGQVMs+OC/oDv55qPLh/1Ja
DdzdmSbeeElzsgh2Izvdi4lNCz4bxZaX9AFslLtI6mSULurQpTAWDUFRWhoYJZsucD4u9yjMJrxW
dEh4WM77kcYWP3KscLCGaFKYhr1CKrNA86fEh7z0tLrntqJEfWJxJbD7x484u5fyC5P0hnIlLa1L
OfdYHLzXiEcsI3lDKzVe6jw2AvRruswUtR5KCLLa/Zqd5hTEAt9gFFegelt0RD7PZfZvlxnlAwqh
6dv4Mm7vPr7s0g621LxvJFv/d9jG3H9XsbPdj51b8JrEOPPnUTu2nwriWPZ2tjjSZtIjP5/Zz2q/
HqHMmvhAowon0mK1Ybn8GdPTisMlkNKHmi9KSh4gha+Id3xBcQn24f2GwwSSh2Z78N1BTZMrYVLU
4Mt8ETxxN25FIwiSU7kAz7eaQzJylakKeVe097QAmRYwyXdfC+UtBPXmgrQhwFeiOv2KvEx/WI1r
RumXp3+YQGpNkAbXSKBUB2IhSRBOC9x/Tnt5Ezgkd1ABuePb8Q6/srE06WhlBzMDDbmpOn69pJhZ
jhx7NBB4eWXNGnMw5hT5FoqdZByawjB7286XJMo/6RcIDhYn+58Lqca3IGuKVsy5mF5chW+GhGwk
galgyuRhYp2h1POeOmkNJ8XkxbHWO5x/Q9kMZNfjDcJ2lqK2kPK5ojKIqEhuTq8ov1vtHJ+b0ldf
bcdZ4niuoPSTBhAdc0XaSjs2euAlLhtcpp1y+1cIUD3nN4xpmYEoiph7Hr9yLXbLbaaKotNE0vjf
F5LMID5az9yEorIS2oEGgkByWlMZ6+kWf0QEcZ9TuwEuBbWmhJa+NFG4kAzHnTlutRALLtdFm+Mr
JmYlqWaGMDIxyKRRR31ZcMnNfaeuuLMfKMROk4gDKJ7fEcT9EK5CN+s3M7O5/nAXbPfv9NobR7hf
XQ4vTfafw36BJ+E1PX4EijHbi/oxRgRYhTWEypxcnRsd2iJY+iOa2ELmYttLjtq8bUIcnsajpcgw
JZkc0zL1OgL6GPGN1RcEgEYJt7hez/Hf8D8zrQcKTQHMSiU3sdSeskpG0ryN3KSUy59sochd73dW
qRbqJa5cEz72iiip9257HJbATK9G80I49Z1PRS3tPCRBE3VHiQccQq0F3ug495uR11+Acpte+AE5
1WDYfCSgMhcEArSc8rjlf0I1ZNSaZnKszepnqM9uTdj3RhB1SD6F6IXXcPQlcaQfUlPWry6cS/Em
EueHeSMqawael25avPKNcBPVSx9U7Ni/7jwqybY+Su0pgmK/LeEMsbq/juiB2xKf6Z260UeSm8vW
yuaxtkPI+b+z9XRYBT9V0ZldcpY4SgNn65LE4ba5mIVhifrFwlANXQbZ3o1CJ26Td5FXIB+DhUEH
K5lyBI/5Rv0NJfqp7u1iTPtvyDSprQyx6wdNC8No7TI/i4iL33fV0qeHlHBbfHo1Y9qlAzUDvWir
9LFvkju3wehI61i9auAPfGPz+Swkzhvi9b/M+2swH1wmnm0LBf3e57oqpYRnnoczvdK1GTlz2g3i
Sq6CQIOdNken963/h4dyIgT/ng4QNel7/ajfXIn1EaShh6AFzMRzIJSMw2uz5Vf1JtfhyEr+tSpH
HWvzgABkUEc06hu5pqBKVLyHBCdLiPgQg39Z4i4vyH2rX6qaq6WbJR1D7bq7Vl9MO4cVYeDyiuT0
KWSQM/eOOgptJCZ4I5Zu1JkFOsW9q6wlEYjCYgk1hSRfc/zareyxvGdRUoOTVtlyhLv+j5VuJ0YD
p1kFFR/txHxHHcJa4sjKUzIQpZ0SGq/QDI8+GhnA/eqS5ctWgooTIyWK08TlH/82Rwo5/B+D1sra
RblZExEOmqSLIgh7CPc6DwiY/+TEHSpVCF4I7VPi080zEtGI2EhzD3/l/hhFjrR0RYAXAT9aqaYR
Pcp3b9Cgr5pI9x1UZZGyo1XKsr0eAbHj1cgdHqaTFf7TIVOhW1pkAVBkXNLMzHeuP5fgCMUknrYd
dxhZf2DzPUfSX8wKBNHkdlIUxNy88uvX/ltweje/IKFNaOpa8qOvLYXQtxEiNKaEFZ21QP0np9Fw
mhW2hjOGtBjZxznSi+N6Ll1q81qprw4M+BZekpftP07nPEwyM5I3eK7FhgKDmJlICONw0VjFAOrU
VfFrQoPmHxjVhBTNzvikiRL6Lz6enAaG5/2+ROaQbNhrYmPduTpFzxyLvfhaoiJuNpvBpKQg8jjj
5NGV6r5dWZ+T17BwXRlgcBndHR3kq5tZ+g9LX4cZWt9tVeZ5chYRm5CQKkSdpkfrk3JYnax5cEDG
lp76lt9qINkb0gZ6D7tmF+/RRG6Iz5E0Mu8wmgeHkcew6ra1G7+mQPealv3U7J4ihZEmB6iI9KcN
K1XjQEfuPUfVRrRjTqiWDKts3Mfu2XXUjiMvqlxYB8EDmqvoKsYd6VdNvXDPu+jSUsTQmVEw3Jvp
+qRtgkKlGo95a6EQT2gys5VbrTjIeJ8a8jIVBk0gW9dnUTLGblVJ5RA/Kms59vjG40Ysj3v2XXUc
/7AA1w+kH436J8pLUOZQ9XM8JIvY9GXbTaqERPt5LQt5WqpgO0SwSbbFT0rpbE/YgDbjjrL86gST
/jXjpvkhqJD9iE8tRRmFI/YWZTUcB5SuXxYyg09yfCvNPhwjIkIebuNTZzZIWguQ9Fmr7HemAI6M
S6VPrP5iesgDRZgQd6qBrViWVdyic1dhIskmdpeLp88gACqUDgAEf54XPLgpvAzm44VodI90canD
67JW92n8RO0GWnUsuwpaNBy6pB//8FGYvb3fbbonr6XS0f4z5HY4Jb3L7he8SdWKDEYk1gWy4HI8
sxWfuOAgoQCIFKUkOq7TmktlR20SaVHsvtU3yBIotXHjUV1l1AeXh7AyGjm6Wn/nP8FMzwYS9bla
74soVc7jhYipXK0rOo98vnHfQZIB9ZZIE6ftiacB5mALX2ch4+j/72BUhDiUGMPVuc+ntoIlpgmY
3vQ9HDke/TJB77t1Ev0CP8vpBPMoz/kcFcONqhT0EdCRc7mOVKPTAtCXvkBQrE3blUOWUwusspLt
N58iDlocEDRMVR6RRc8Bb6vFJGpcO9j4NZqBUX0uT5mfYt6UowbByIjHypR/BUCmt2Obgi0niDyX
yieqMjHTtUP6/723tP0NsWaFwvB4sUGgngmvYEymx2JL9ktT9OhxJS1ZH1oZes+WeBvJgP1Vrw6T
XYcqJupzPAasB09hJtp20OX4xS1rEm94HYwfvK0snJq5YQOrzxfOcZ9d1dNOuPDJJS4/l6JAKcYV
BFSTtSC6EDcJE/g5MKPShhDUyTyJUawNIUZnEw7yZyrH8JAQkg7z2sP0Lv0Obe+5PqDTCVrt7Rwe
fVVPr6y7HBkqWYXudvQDaMa3NS4KtrABR9mZm+m6mzwLbb4XECxGINhlLc/2J34tOtzUgcRTeV16
n94e1x+ySZNstE+HpaLPVvH/p/GKQImoGF2a6LfEWwUc4qRcgosQDeHHUQBZlhs05eKYqN/Lw7yC
vYBmXGGbmIVJ5O6w+IqrvdMs6Wz/10xoEoqn7maL3A3NuiYaKBdqPQqonujfBXx1ZqTKGBxAhZl7
IRnYKIt6yciPC5mfRQdzlZn3biYWpWihBhT0WrimU5wKYbE6F0OldEzlzeGE/3wae4MhGYGuKIhc
ociEvt/loXHlQQW9Wag2JcYvFI9COwX90AytVytHLdgj2LDRivP+ba/0LIxSrO+PlLFbY+erpx/Q
hcPtLiJBBK28EeBd6yAMbB+9RuXRbd7IJO58R0Uzz+Iw3G7vfW62A0P8nZCdr0vK8PNoLmYfPGK+
1dOTi7Q6w+c1yHZEwcLvoI8uuywURZZFbcOaknlQYQ7VvWrui7Ez8YHGO189QknkF+XBB6ETRyDV
lc14nRo4tSmpQPDf7PbQX1C2HHoDxnNlvaCrtPGaxTAGvphSJjMdrGcHoHSr3q+ktO7DGeb08uHK
9lgl8QQgBBdRE+szCuoeuJXHiXf3QOMg8xJ34QkQwf672zk+4GjJNTWmUwV+f05fSzw4zLflft6+
8EolariRlei/J1NkxutNdLrddMlnyVyiX+nMN8085vAza3GFvrNkLtQDOpuCa4aIt41rYmO9pSAx
8TOxfQPZrTxTEdAMLo3WFFBrdjcJaIWHBr9URXA9yMKQN/63++rtzgORvxXjFNDJeP5TwhzwBL0H
s35adO7PxRlrlUOIjReJUBq67iokMF83n9IRbVhldFpqnBUSAkBPImaijFbAgGYqCV+6ZuBB18fH
PrUlcXxBp7jrzFZ8vWJ/gAazti/cY0vaA6vt6GvVup8j4JdQIE5mi9eDLJ77UhobcLJSkWX60fkx
PpwNzvzi6UKen35gHrIgqdF5nDvAdYZbIEDsu39bapniVQ+sqs2G2Bc03B2N3Z1RzhJwwA7fVnsc
pCTVQAcTGqo6wTfz923E+ysbkluxnvA772QSklMH6WxkkTyieaBsCteN0tkOLqTrd9W6Vt61Yj+t
2b2i8LT58VJFJNXs6tO/+GACWKU4a6UeJjx7s4naOpwdW2Cvii+5Ov0IAnT7Vgoj/Q6A9rezs7kX
g0iv8r2lwK2yJ64K63E4WpjT+FkGIchPinx4HVpjui8wStaHbnaRNx8x3qreF8kToPZ4UTz5d+WS
KZ0hUuIYEoAeXIyuL8IT/Z3HIX64neDVTHSx+j5CZXbrKLOCZPiowm68CdVBEaC7TxpSKa4LpFWs
X/Xcs3HHf+24QRqXPyFbgASx8I8nV9+sMol9o0w5/sHUFZC2STIMjE6eZWR7RaKIHet4jGVZaihz
BSBUrz7bjF12My+MBHIOka4kpwEANQauiBP6pJY2dro6y8D61+TJytOrplznqMqt8W7w5x+/Ju6z
fXrRfGL9wJusaKAMc5jDsfO6DZA5kJmwQrmrEWrNQZnIuGmgc3o6eaiNA4DI1OzBTL1Fk3OV/sXt
ZCklRftIDa2PE8zL5AMbdJkUsbHbv6HRMMZ71V9KlTNcNYobPqtbuJCUYfKkolHfdFWao6ImE683
8pnQjO3N5hCHq2dsRO8dvpudq8iqWrkuxxDZiqodkTwG4d0mSzGgs3KORSBfvZFG8MvbIYXJz8Np
IhoGSpvkPubvryJ7n7BIXxc5kAj/oknTPY+osAO+Cp01hcev2lvpqdkrSvmQ1zSr+WvlXRQFoZqR
WYuvwqb2tr/F9s1wuFmwiocCNMQ6DuCzEamPVsv6EzDRjS8WVJFoLL+W5TJtJu3D7GZXMj7Q1lTz
bxio41r8yvDL6SQRRxCVQQE5AMkGAf86/Pao9subdV9rAQgpi7tTSy0ZmesnhyscjOdJ+0aXBNnu
1kj7VgiJUYwCZhBP7qjZbxPdhspUiTrzwMA0qG7Tr6S35P1X+eCvZZGXSjlktLzft2QP7lxjO+D+
EhiJ0LNbj5sK1aO1DtCR1zQe73SbHHLECS34epqSfXwaURW130mdhdUFyYvfFZCPTtt7f8QzAIuh
PTZogu8umnU43eoA0j6alCSu4pY0cKjF6Wk1qFlHEHp9kmrJAJYrbVTQed9L4YIq5XAbpKdy6rsV
/P91shgR21D8hVEMqWerNcJVi2z+RxuN62V5F1ONmJDJCm6W5ty0QAdet2EBRIU516HxTNTH5SIh
zggrPm/DRTLBdYJhaUD7JDmcTTkXhAWpBNcRXUIuvYDwmtIqAgPy/JoTzHj2B2o2cbn51b1x61yu
htM0uRhCoiHkbCsMrs8u6ogphSO59OcRumDeVHQfVHrt/Y4lSvm6B80yiodlGegvsC6VADecpdy1
H4Rl5AusVIwv+sFb2ktCxl8qAlOPOVRFL5BR5EQXcVxYy8y5hn4bEeaI4yP6+cwi8CU+ZU6fkTfJ
i7zjqUZKqjiXbcQ7uWDqgN0TaOy9nQSMnebslcgtBPbTz5F7CRn2LDQZWYPJNGy/mQ1R39DHc3qd
VHpUdLNbRHAnC39NgIxT+ZSAy6dhOsjCID+AAvAULKRC4N1/ZRGOMLEFoQg6T+ak5GwcwRB5FjSx
y2XNS/g/3Q/AbWRxoa2FwBAuqj/11w0k+v3Mi3sLXcnTn7kXmHgPlXJjji/8wWfl7P/wUzxa8H9D
RvopnzLfdJrdyl8CjX3rHX/Ii1iS5Z444cynmHUSgH4xoFbG8p5WWSBPIlEWqQyX+OioKFL9R3xx
osMQYNfGqZ7pZlOzbKdct0iR8iBTwTvVwXIOKVq4LREZqoBOWmt0WQpyMWoovB3xGQCVkqu2qz0v
8MkmvbfC+2Vpb9iwd7B3RnY0z5yNeAQ5GQass2wjs/5imS5c/Txio+S09/Ifsrt5SDyq7lvA2/td
kpSaJ5hdhkz8u5JOnWsxbgP92XWlkYZo6ux/gV0YQKFC+i5sg5VNNDdYNc+DT52VWztLhCSZSWgv
/qj4O3beJTuNOxL4PTnWx645r8XKaDYEuSZ5lUUpHlILCskj6axMEzpM1zvTEL59PuxotpIGFC7U
Mnvqn2shAzrFEY+q2FHFYsjBVYVHdL95GzVhS2kTxBcAFnGYnLqntolAOOrz07lOgvedmzxjb+hI
ZROI8t9EU2meVuyet0wvzEKDkVoWTmREGOCNKukUeNoglRSfkQLacxRmON3f+3WKoYdwepw3V+5v
mtlfjPKV5ai8PFFq3ghGh+V7VyUfYLO0vyFf4f3Byy+YUfN72SH7vvROuF19OxpokGgf7P6t6jte
o5QjSjSjdngQndSUFmwocanua+YaZd570MOtp+Tz4ZKg5DwAYqE7IlJ1M4o7gHk4tTE40itVCmUj
f7tLVjJJrDa+wnWYy1O7sCt/BldnW0B1dGUIs1Vd49OKQ0rK1ErD1DiCL6IY4Ixpt++LyGGeZpka
YKELjEJGG1qyp+SHkkeOB1Ul9tez+4+mMhAsS0K/5UV/C4p1jQayG65TRxOenXti4q8vfhYSoWjQ
dYdHiKk2UX/nMKex2X2xWE/Jfuh/YbyUwFwzCklGxkOklVPMT8aDOLXFVxWBGOUK/nax/gMa13Sn
sT7V5QDlvo2VJqp7GnLyx5TltStevjTDJBOVgO9KTOFg+IOuyvc7b+XMeaKR3r4P6VG8dy2DhJxS
ks/bGANa39VFd5MRZqobmGkpQSEgcDEPrDdNgPiK/i/PB+Mcr7s+r5h6beaOoFZevshrlQpKtwdb
JXZ0MaAjJQqYPZCuC6Q1uKS89HwUJpEI2DYDehcWYVVerqIvOMkGzof2OkgSE/5RJiGQvgsqyu+V
TGPMAdh9/ji4RKghIOi1JsMRAJvYb1cEDwvlPllL8ALu+eU6XJYYXG8eP6AFBriuaS+K2GQjH7qP
r4IKAom5ObE1TJZVnvzqHgfyjMv7pOEWhFyxTcU54T5KrW8/uSWfxiJC41DIlIknCw2LmwcYITNx
tPF0+pJwClWsDuhgN6Ywbw5VshQRcfJBRGHR+DaFSYU8cQoHawg2MIZoAvw/mbpzZi8OiyeFPo4j
SVEdz1hfg/Md+i60h1Xbm63d0oLeHlChlfHtI/xWLXM3zJfE1uZa2NKDUBgGpkndaDp82es8gfIb
cTxfpVIktN0A0BAOelRr64PUx5E5/3tuKUXpsPxtRrN/jbUe2LQtXNr5bHAoa+xKF+FVhGmH+//Y
i1aLuTSvJEhZgejyUmwNJAibDSeJSuJ/TwszailBS5zdS6XBL6ryGTMLjB8gMMoMnMLzZQUgHnkL
8ffpEhi469XVPJT+rytRh8f2NEDKDzQlMIgmOAjugmglIIJxyB3NLFbxnuzRYs+vC1Rc9Orm44do
TymIVonCCETNMjGsnvP40lH4rvMuFQKTzPsAcA9kGQgcWfJd/Ol7V7G1OtKVI+dn1sw3xAwCuMAq
ETIr4hXmoJ+MdfvqX9wt27L0ii4NMO4GyW2vG1bZTVJI1L8IdD5MnysMKnvjRzq06+vUk3tQnsD1
pQfpzjvTXYtNsggCq2DdydPuXj1swKzpsPFSi0wVwbWPM249IEJwxvzT8c/KcL99cOt31o9EB906
RczKfkj0Eb7kRY8Kbf7i8Z+5P6MnuY2imJtffwHXbiEZvqZQZ4WiaBp6f4KAcaZ1bQSuDHLsnlax
A1Z3gNqA4IWCw1fjw4mWMKkeYq4zx0axOrCqRSuGYjZo3wVaCZNJNQqhpnkhczz1DAYxutna+YT6
Zy+YtYQ6STr5bYkcWGJV3p6ClIxMHGIENwmVY1RGX6go4vuDUkiGRU2sbL+yrMK6g0Q2Yf+5p3l4
Tty3rJAa7VEjc+wFzR2KhKg8HIhZA2suLAxXCiVys4oJPwUeLzh/9Q2f8KtCcFtvdZyeRNwBT3dH
DftHKhROIAK2rpOIkas2rf/Lj4dWFKHUsA+16L1KS3+YCPoUEtbKIclwzshAr15oLuNKJKMuPZ8r
MD8zxe6QKAJII0JyB0g4kP/PIdzuCs3PbBkravEOCX2IQW+elx4lBFXnOScgWW3iiqbt21gAIbXz
qTZ7MTxTUo/aCM88SSJJNTj7tGW90rOIXJwlWgDSD809Q8hNe0Yhsl5PrQyx4/LnBrSz5rVjrm1R
HyYpY0VSg08uF49em+UiHOpECOtMUuyhnSfLPMkL9/0Rl3qQ8PmnR6DWpBJSoTVhUG0GeADGIMdo
xZ54zOdt6mCazCVCkxbTKtr7C61fgZ1JzI5K5AGJ9D9mJ3EWrddYjnyGrI52Q02CdYs/UNfIEC8N
RW0vYVBLBho96U6oZkLVUA0hvd9cc1qaJf+ruStt0GPlRce9om2WpgereVndu971m45vpsrT4nCi
lVhFPhNFwdxncuwyyv0bGtsqsD2ZzsTAXsrM4OFvFvGLah2xY56kDvfk3zwvJQq2NPwAFGwUZEBP
R92ESpAjW8b4YYMbnFAxfkD5qazmT7GxnuWOFzjSo5O0dbzaiM2MqtyH/rXKZCMW4GrJKM+yGst6
Sc+mZrGZV8jrTVmGvCTgyfrhhKqxbhNQjG6kMw1on3QUbgWyzlxNzzT2VqL09hyVAiuE2SIO2Tcs
mBB6H1vAMYxNIY0Fy2zC+fXeO6GLLlYwOQucOyeC7qDjURr7RfH90OT38YKJZJDxBjd3Lx1TFOzf
FZDJ9xE+5QlLDhvaNFWCSph5mwryb7av4yKZH3OAwPNW7oZEkEeOpeb62qCJnZah/b2NKPECV3pW
CLgJKw2EWG3f2rzi325moVjehkG9VO1hEkNLEMlEw0zT1aYJyqxkiGlMoYPNK4V0BUJ7wfl9kYI6
SUWk1kXg2WN/14rYXCoSKC3BjDK6E357iFF4YCgaInBhirBnzZd+y0PGY/Uv3A4XxqH9AyAo2B89
lMpEUTkszO4O2/AhCsBnNKL3JeDfEUwn4eL/ToDnddUhQSQLO0LFw5VihPc995RsCLUA/GnZDTBe
Mf9oi6qvLQCIc3PWo1r3tPMIhZR3XfaGUYCIoirdpSsPOO8mdOzQKxkbRbN3BpVft72rPXGSs3ML
mCVrsVSzAJ9BhHo9FtUAg+RVEW7jkTSukKQEhx8WF7edLXJQ0ACifsc8DoU0APE8+qk1NSIKGb49
vVzHaljiwSufoSaPNNIHarE0l9qLZEJ8VAj1m5nzJAF5y2FULgcGdyDIf5TauDGztBt2hgV7tAcT
1CYxgetOvzFYWOZjX/th96fIFxKD/LI1Caj+XRtVk2QMhUKkCuFtmYrVrn3ebyHoAcuNqZGh4J39
YmUucZWqRrZKf+PvgDxg7cm6t28gEJ1cV5/wID+zU2SH5ZB7lNlYTATSfIGTm5SSyCSZ7tmygwru
7PS7+ZzlQNy8JCzQPH4VRbOuFHqBrliXDZXL0MJyeat2bOltilQ+o++JVzZn1CGkkdKnwZtwtgEY
GV2BqG3EKDNEokH5CmH+NCjiqncaZibHlldnzi1JPLr4gAJneMrTkiout5+JeVxPLQr7b5eqQs3C
1MMqecyrp562Ty9CaOAo2xkfWaEpBb2gR6ORwRHTqkh5cw9yV0tpwVXrnGcuheHWZfAkBAaTi6hQ
eSTpmo6UWMhQ+yq2bLBqAbSe+2AS0iJZE/yVc4Q4oIQB4rW6lQlpbZpzY8uEV6A3i1pkwcSL/7UY
ZgIERJuFvFZEQ3qIqaQPSh7mwbag9yW0FImqcoZOVWsOvuv7/xuMaBRuiG7w/VaTCRLzMNimcVXj
/zZUN5n+9LXatgUqkOAdChgJn5K7brSkP5AN+AGrCVN6bmfxWrS+zGddMCLnyAHRjD7Nyx2YT+Tq
gDtDem2dwBqeCvIFs6m7e3evnTt1cEv/AhLhUXASb7OBnHeyoUMlGp/NEf9jv7P+dUVuG0+XfLaW
SfqM4dyG9jRIdBtUaNfWba0xb/d/sR0/KS5Ch2ZtmRlAfz3L50s3u1+hT5H66wkgnDru6eqnul5x
01+iLxersaItdx7XxY/ZfG216s2b9ndQuD5TpJ8o/CebFMqkYmOw11PskJATzIojLkNL7UmUT/ou
tWWKk6W7ucZYsObOu3ngOvfmrDChEpO8S0VhoyOLi8VlgdZM2vJurYkD7ZWqiqHqWwTO/EObNCIX
JTF3ZNndqrjF6zWzWVdqa8M6hvAcDBI+5Qh68UeM1NyCriDnD4Dqm24HtIsRE+XiQlheaB4+qav6
e37eA2eYHUrnAJcICF1PuKtQpGhYKmrFLKVRbKTBypOnAp4zN9o7bd6L194sfkNU4QEIIu3bTDzM
qizkwThDS7LtKwvD3gXQ31L9s3cfX/iQlppYxNFcEJjI+kLQDi6ToUsXCskeGE9f29FNLhGyZLdY
1uiZHnvhXG2rjqmEuXL6yZwca9W4s6et8KzomUWbqmDy1fHkFABbIBdosPJ74y6riaiWPxPzJCjb
YruNZRuJ3AuEdbqVOgbCLPS6EWs8idmFekIXAOx1WXWgiMBucojGvwmvXzXS7xOCKu5VGa4MgOKX
AhUBEXG4qYCCTdZiCQD6Z99LVSCQ+wmjeCTr1Fdm++UQMiC0Mm+jmDTAUmu0LTADb2KwygaqhD7W
NvsmvR7sZo/0w0XYFQJ4j3GQWqkY96KSL2kRlQu2zs+0Z6SqhjS/PNqWKCeTCwoNp5+9kCtfXtdq
wFxEJbGVqv9XFdHZs957PtLuE8qlbnf2+Ts4QpxgOKRLj/M/PkSy/roP7l2nB7WQsN46T3xaBiuD
/fbN+P4V8cyK3dTPgHoQLDj0FG4f0CkpW/ea6O9k4LFH44pM/za1fY5Qx+gV5GWRc425cg6A1M9n
SZLhk8yUYfyEHjvcdJD5XeYU+TQ9wrRUnTcs7C6ae6Ls5velQSaOZUZ467dPQp6lVPVNm2dvEW6v
9n35fFSDBYcVSZUxGp6zanWDtCkVHqQvWycoh/8VuLrMB1DwZAnL+Y7A3pF5Qe7nKcT66/EH3U+9
ObOAyY0u5Se9CaYMiWWZJwg3P4o1G/jRw/Pxtu9NdNPC3D6a6HZLcGiPkGmSbWMles1r2i4jK0rC
8EY44yxkSlcA8nEoEdayTeKUJclyB+2XFzM3bYq0iycjk/TYKxHsHR4VdRWYuPs+rmGAK2TnDX3h
Y2teRuTZ3Mg4ulELvEyy8z4Zoga6/4Swz2UiASEFcJhxv5sxa3pPdw7+CIBt+zgT0+GMtKHuMBXC
mzj/kl9jkpvRIzKN75G44OmkwD8ODz2SGbmziMiicWGKEgWtC7M2uL1AFJ9jEooRLOsB3uQ19irj
68PiW28oSwyGdmd0Kd7uDjH5nO/6tODLwo6ceUmS5lCvzKMyQOmi1mhepdIP02kNJwvosyRXpgHo
UgQthIjBsGcHiWn45xLsLdPxfb3WqvPbRD9U8v/08KwvLx57O6ytya8K+fsAgqwT+OKqoAbUhigE
RKH7pAEmtVcDy0j9ZxPnVs2ln+wvX0VtUpyQc6n9mWfpZEd5NGUVtsQFPIJHPESNIKp/Vl7k1xfJ
2AEgcDVrVgyd5l6/wUP8U5xk6ceJ5mvX/cyOSJNmuXh/Ge/4y2BXMaTfqbfZ18rCldEaYZpeOhXH
fgCwQy/XX+jkQaZUDjC/kSx1KqWUe8RfJ0jIjwjsvw51WktI3TImOQPa0P+R3yBnE81jFCutd/5i
6Gqap9kf7Kzw4zCRBKMjMbuqoFbgG1GOWXEp3Q+28TkPtz4qqFnFbFys8OSuENtbl+zEFCsa9inQ
4GVftY744voy07YL4xJxBxyTH9g0NFuvQor8pmxCjTapb/7vN2kwcWWb3Za5BgM7VqbD0pMG0zdm
ayKe0is/xqu/NoAIQOBIOeMmjV+T4A2Sjzlmgm5yjCYhAaxIdRxn/SjtcX66QZuQtbEX93Db/6Nh
FC6LazIA67DgDHJkTpDiVh0hlOpqYp981TOAIdGWKc0E1d2O7r90v/SaizHDyaD7x8stJOscJ48M
rrMWou3sjW0B3s61xZ66ln8c1TgyePxVT+EhIN27bliYk7Y4kX0AlhIw0wVphsi448C87221TYxz
fajhuppZm06DclQpxMsWntbdrBZV4mCTsv4usSKDvpHy0uRp6jw0VIfeucpPByhPdSazNlelwdZS
SULvq4HdCf5bqB2VXCrRugsOCvljESW7InEOwz89BqCQnElUHis8AGp1XyIb2t0c+rEfqPup/LHO
3TZaJwo4B9SQX7h5s5hQl0vqckgK+QjIHpbSbV7I/YmL+/Q9GF6bKA7Rik18iAXbFztq6GJWH5mz
lgX09S924RON4uM6Zqesa3gAIzdYVlXSL8xzhOhRJ1Q4gkAKN1qAznPUG6AkumM9JC6TLTZS5Odk
31lhtDnkpG2S1yOLEBwAwV8RQgLkUxShZG1KTPUoWHaZq6Cl7F9lcEBxcRGc1Wq79NDTl1pRLPTG
feYuP3G4GX8jHqC5B+YILrEB1ph3zmgf8Rf0yVFNyB2ttG4WZGERLHCSmSdsvFuZZuU9wyEvaBbu
ETrKd6JQL7GFXURH3BaNd+R12WOtQ7zUFRzmYuUmU13CrBCEZE/k/BSftdCLQJyJDkB3abv9JwJR
D+TVVS85e89RTRZtcGlGSL8huSoT7oBmHPkP6vzbVUTCQowTfehujMk8T17Om82Vc+VrC/VyZtPP
1GCuWSMIhBQ+wzXQ5N3e8oCb8oICSgTZX6JX56le1C03f54FL4ANSApdPoIuLXP+AXc8XLu+vlFB
8s+5as6By97xaJIcOg3Ape7ZxrdNdJ4W9mN5cLNXSoMjFWinLwif+p//YVF0qe3RnOJKevlmlw73
F2PJNL3D2C8BW19ANwE7NtmQSzv28sfsWH+wW6yCM0LWb0Cmo6K2E4QHQve3RTI7FAwPp1iYrpC2
vHHSmQnF5mDcwGpzRnMCCHy/usQ7dswwEDkYRsxjgyyTrokmnq/FSyCSBOwSiRpJhA8JddV1D+2Q
NR90oLfiNW90t7JSb4TQmY15DVuCfziDBoBli7AfHipNZsSIRLxZoIw1QCNmuwS9kgp6NmjQcQA6
k0ek7LOiE+bJjCNdNmD9/WJMnoSpeYbjLIV56XWmEUDLZYyMxJVLjQDwdS8IGiKQKBVnhqF0jcS5
zevfurjOMAIr4bQiEuhpR/hSdWRmwn4nZol4TElUSoXxpO9WDfiNLdAfGUAJCQIBTOVXsrNNY1IQ
NoKDky6ujVTD4tU1EUpsFsbFgFAFPDk68ColPIJW13XYwqCNM5OPt7mbcaD+VIT/cSlVGZribwLn
2/1zIGVgGs1TohD7KxOOETvATeuI5/Tq+ONHzRoMU62Y96dTBlA64HSa4z+PdNHVjO4XAkFVpi8B
Hve/IGz03/5Oj6gLyJ1QXK8eLTdZLyj7WbZ+yR1Wnk/GHCihK3DqBzxrzsMuimYL5jCAzkuNk/2Z
InSkf0j8uQuxlLP+b6jqXvLawTTsQKp4BZn8G841SWqYH/LltIJed4m0UxWvMgBL4r9QbOvYZVC6
dLYxiaws79BBei6LE23ooNG41xZJy+BNPUkE/jKO5mrnxeamhpJ4Aw9UbPnN5bKlRqLyYWySqgg4
QrSE17M5yMo5f6GMp2CqCWoIar8wC0nbhMWIbvMvxdBWj61neOufOPFgA8bXh7osI9Pv4vlO01YR
8bR+l2WU+KGg27ZV+Jb9GmcZSA8BWrVsrVu6nPUtSaz9qfoeObyKgvwCQH/Hv9pH3o3tJiiRui6u
V9yZXGI050CodXwJb8sLTJei4TVDU9V+rVq0tO9xqk2OT+0FenuT0U11LA/lErj7nBmMeegZXZu3
5LO1GpHLee1W455CGIddx8W4yjsEXczgpHTZD3KpmItVSvddZgsA7pze1y/WBSZikEuVdhnxbExI
VDhX3DCjiFmuXK8nttuuNh68+dKI5nHil/PT67asZ+Li4EUtRvqkciTK03i/IuqqILhZs6Aa3Sl+
8EYYhX1LcYeYv6pivVZeoxYWu/08j5MMZ5/Rt6jSCSBGJdKjwKbLE2/ojVxxlmUmfxmDUGNPPzR5
UtgqtQfcs6opE7D5lrHIdsQPS4buyavuCLuAFDFhQMSM2zhJH/mkerp21Mufrdp494OdYNx205xr
gRDICPO7dcHSApv4EiulcZnc9gC8bzhBKdhAUSrDk4vjXM7slCcWuA/x1fpAl7DGURhOZcqfgall
97GqqtuGJpqSPhXz/VWJbgh1Md/8F+5x50P4suCTXbd7iPCXjO4wH9e32U39JxrFnkRMnLTjtduw
nWI1PX/q6iqIHydMvX7mWM49VKIP6YWugzlvDjCJrCNPapAvnU6ZtLWq9l3V9tV4WAK3anhNETr7
qhVY1951KrzqgR7GISwJC4TPvPRJ0WQWQg6ghl8qFkjxC7RO2bV+wcYSfyGJT84nNjddWWU7AXN+
uDwGUAJrlJF9y7tdPlkZPyEOEGOFDO9yOEiK4xByD0KB4ilQj2/Qd5WAC1oFZUdpxHD/f3fmTRzT
1P1zmdUp+e72vyJefz6Sp8mDfSJEq4AXSX3y8LrzoC8RLxEEyAJ6lnYCiTvIkxGnfUPer33R7f1g
bmMofWo/Gu7BrQZFZwazm27Hq9IMcEaVb2rXnTngroHzno8BDGrKs/b+A6OVAQm0of3bPqhEJbxb
zLFn2GxTJ5YNNof5nhv0Mh3GcRz7dOLseTMFGJKls1VTvhl4fX+tIJoS/eEeb1JENnBsEVGrTlhh
nZH4gUFL5FyCt12cta++c8Q/G0Y9yuAEAoeaLapSBZGYibo1W+gQCeADdNCwDMQEvKOnefuYZ4eO
V2Tv+Z9YWG5cy16qa8OqRBCwq9AN0SvioHzMiJps7ATCCwkW/VF+uNHCQLsgpnrMGb9eKF7XtneC
t6kC3qI+l5ClJZRNmsBpgQdWV4QqaA6kAEu4FbHkr+ZBDgaxJdvLNUuZ67IyrZpbmbU79wB7NZHd
cJ2b2s++tNHGqL7tm8yPPWgbTUyDfqqDaAIugvN0NrL6x+tIkK/kiU0rqsrGCSFvKVC0m9cLbQj6
99A4URH9NSakBhL0DDvHzUxGAqXAZbz6z4rJt+hhN6KKolvUKS+1zZnv2NZXiqQO9F17kzz2N+TK
BRE6fXounGhXhgE15+JlU0YKz96bCNP31m6Curqt3FfPcaSeqUJj4KcOR6dxvkCRx5L14IWmwUBE
+nF1RnE8CB4bfkrp66Lh/WHlD5cxWfUyqUPatEGCAsvl1n5TS6u1hbByVFen2apohRUWRDjuXgVb
jk7/z8w6R85FTz0VkYpZobmE9eXlBzlYCrcp0cbg4M1wk4RrHOwYGo2TKq4Odhn+HEOQM3eXFJY6
FEsILi1pBrLl/na20/fVBRecvHxN1Yw5gJiHMfnhQr3K3MhlcKk+xiEh6qcBw9KmgH81eNTOWQru
xs8P42ldmnJKwULnT6YDGESxqUaKvgFHBbnF/u0LBX6vzt8Wb5g8SMALPak7VhJK3Br63vsEcr/X
NbcZuZNKmYCdi7wiSjHnae8pOh6aiH9B3Ai5Me6CqdV6/9O4sSKz35PZSxk0W0Y+VerQiT1zgMl5
9rYeKV6zNTB9UfUsWQUBaDD/sesWdnO0pCwBZg30WLqsnuSCIS5hjyzLvxp19GGlCmkSXEN2WbZ7
kTJE12QpDHHNvpjEhqk8cCZQukvjrlqKglhJJY/6ABdL3sNhMSQ8/0RMJEtSC7ixVn0l5xnmlXA3
UWRE+v0we0kwFN+FDiLB0lZ3rGpkQ5vsIGVQISFTtbS6+Cb4twHnl7HZJL/0jo6fS9tUemD2SPef
vXZMqtskFlGlDNBq5BbT5I7h+PWWXIDIFTv3QZvDWPtif3fhi+MstCnaXttE3Lw2x8cCgbq5/bbF
kuy3/1dFGrgh0klcswvq2J70ArrBCXnxcGomIlpLuAn3FTr71IGuUnl+E1H7neAcm1L3lRJeVTHG
YUkH0uUIBWwCIFmJoicmVkMqC5aRQbsuwjkB4wC/AfdPCyqqkAAudVKdLqyD7wiF0toBn34+zotj
/tBtjvBrGw/4pgPHD+ToxI10foOdJtOPk4zf9gGNTYz7etJ3Xqaiyp80/7oEgPuQcqy7egyAwBKD
f3HT3jturTKxdul8pVhCYgkdk8WdyP0+0TKh3SrzCQkt4EzTsGe6G2u6rzu5TEG0dsKMVHT8sL/v
v/aZOclXOCJwqPD6RTDw6S/lDtOqB87dq+QlwxrZdECXf2mQImUuRwPNB2ilRvCdW220SEtB1L1m
l5YbXRwXdG2Axa7n2jhM/ioTd24QWv3rBGRlnaDNYN1s82Qo0DANUKPSaz5vFZpF1KtFxTAMeOKf
dWWo4vccA+kkngfvMmvYs9Sk+3dn1De5JSfWeSvGmZWc68EfLfJk/ILBQNGXYb4qEhrkAvto3E34
1IPtfiX17VUXqwoq30gxRN3vvUYppfnnLYi9GIB8n3KgNfkvAfWZL+So2dWNZeZC+V00ta1KxlPo
bE03cE+j32hPGqiG+BzjXOsi/KQWaznj/1ftIBE9JNClFt8WcMz0hdCrafVoBuyesPzpkg/Qd5Mh
vfNYljP5oPAnNErtNuFIdhfWlk6XuPVZLF3tFurbHRECAWUlpzszR9118tCcUFPg8a/VcB6eVBAd
b5y4MTQh27N0SHB82FEu88Ff0ohoHsKHjD5dSanKtO2Y7Is3Vmv1mY7xNuqi+jqkA5zznegj5ooV
cz1dePnzCWFLf9c22H98SaM/q0aSZxWM65mI4I0lbJbt0dEdPdNqiG+f93eThvyyeHWbnK0OZJMG
UJOYh/T8bRRmirwpdMV7a6zo9fulfb1dN/yZljKxClvuRalWU6vuVHCIqgh9xfc6XwxxD/3+bfUP
jCVM14k5g1nxdswI68TKStynUFT3GTbrsFBkjHCS5AHCDkB6taDfM8dHeMIFiTJCQqwkM2lKK6tB
sAG8z5jjR8VJD5Oj05RL1P/QTXtNjaKRRhI1iPm8sQ+P2914iNt0Zm9C2ME14OyQQOtrnoBYbWuE
tVou5aTdyniyR5rmpLA5f9EoMd6yaNMjaVBVSHI9+tUWvFx0hsOaU58P6X2ZgOQhyCf2ZWJGfpDz
maMo9KlNK7OIZrZg6eSTseXiNadRfn59NqUH3g5yUtE8WM7xahVRtju3yD/LTnZLDpkrWnU/DFDs
tNF8D1rqnLnpoBH+9TwGmWMqqM0paJuks8JBXsCXcezn9o+99kF1twmHNWGHGNMF78/qXi3NAIXJ
gihEDwKMfnOXk7QwwHEcahEYWRAM/CkTMPhaGLm7LDHOgRCvm2l+tKHUCHjXCSKzfeNwEFpkW8Lv
Wt9VpwWPT6Z0spE7yaeaxA05SIdOZ+huwkbOAlfx1TV+aHKd0MUGFryDPdj0MizUXzV+CjCFsmpr
ji7OfwtTfB4x8XjsltPKNlK6xzPAcgd7ig6V94U1DG0BPCdWwJuUV0OGkTMoX99bli6owxaHfvww
V+J6qUE1L6hbot5oK+UygW12Ztfq/tm+/8Ed+2f+L1VA39FWmW2DGly/t3La4TBuinEoXs/yMU+S
mHuVXZKjgHX9bQQWFA+BQ88AEQAOiVvi0CrTxoVuvv+xFc4/nRdpXnY/kYMImgwKKzk/fVdViecN
FagZbl3biiQfiozMl7lutSdBLhIrvCtw1oQIBCCmCCBOpCJQtKDY9F8tI43kVjegP3j48kNJfvgD
EvLqCBA/fuA4jOg9knYLz6/j8cAHCdIwGYU5g5b4klwu1S35sxbn/kp/7kn+n/ol8ClVFko5Dnir
n1v8zcfGs2bbUh6iwC8H57Ya2g+Qk8Y9fNULJGyjFbjuDKyh8KXOM2nZaiWZkf9UU/ILclARZUtF
4uWJUEF2X7Tw5Xp+6/GVe55LnWW7YUW0SsLPdpCxxV9Ft0VWYhgMVjZYeAP2qmVUho0ijErTqKTk
561LRNgRcLkBzWiRoGXgxuAuQ3cRWoWvkkAFsGrrH1ZvMc5wQp45ZWDWbSTbVsQl2JuHsWTGeOMv
44RBga6gOCOYeLEbgLnA/5iKhTG/mYz6X7TYn98TbL/FZH803Uob8c/xOTA9DpXJGQefd2s8WGSS
hb0nDHOZPrMvtPQzaf7tKrXt2B54MXVRFnKgVozDtdD2CzA7sOuaPQYjuYA5doscjxz+25hvt6a2
8jrSWBq3GeqUdlPk6q1mGKogPsSpl42u180tXBkIHbJsUZXZjo11hD7t9kiNNhqfu11OsGtdTtZz
3PMc54eIX9raJhYAtOk6eMa5epsx0i/N69C5dcz/g/Re+SgWvsaAaOui1NJj+Ro1935CTpNb4iEk
DL5s75Pclj+nYGLzuD9iHlEVJxuQeRx3xi/4yTMsVaYBskBjbOueMaskD/nBg2Js6y1KV96vCYgO
zzbyF/56aqlObyBFbtAaRzHaT0V/bjJr2vN+DnwwuHtkYF4sveCWdysW4by071ZyDEloZQwPMDvd
PR861N48e2AExTMRvTiRzbT5I86sF7C8PMVmLmITsmQLIxEIMF5Cb5inf3fsq+0Jknqbc9/IQvqi
+4UQAhCK6znLrITSU42A8h55sAiIUJvPOu5IVh7wLB7UKlk+5bUJbBbtUIb+jhEDl9gFm0fvVaeq
nA3acR32UmVWRATNk8qoYCHhDBhbfE3QAZQgCl4wmnZcyYsjxqnCBv9ed9sg6g9vQMTdNVtG01qy
2zXPiH23xu+kT9kzvbAiV2x+Ev2v+MGDnEGOfMPUb/6kfwFCC9w5c8eQoCX9OB6ZrTh79/QxIWEM
wBKXizGnMLE7J+wYgiVJXFVvZF787wLmFtqIBS6Dzh3caoDmsDPZAKLnaU/dMQkMtRz14E8qzzxG
q1O34d558QS786qK47APAGOdMgu1O+jilanqshGGMzaasLb0cr876fQyB4nAetHKr/1Wi2KWS4Jo
A+hdcSxw9KM674rWAaGbq8Tz3babDYhDXDZB9+5jte09ywrS+c7ihSdoSP+39ka5S5I4iPP5eZEN
ODUy12INBe/HS2ASNh29elgknPx27zCOavsv9YZhp5xqFR95dugME8CvLDN0z0JApSTV+OOs7EFJ
csD9GeCqzPO3faSxQ8dxrD+y99TVgEdfEf+dwdzcUzZOIg4swY8R5Z03qHVDeWi+JeMU3hoFRSgt
+HvVSnar44emtLqODmiZqAcHqK+4ABwMCLLEodPDb7fQr1OwJGIwsG71YBCpl/MzAIsinnfrjPKE
uHLH4QV1zSRikFjDlr60d4x8s/M2j0TUus9s+opn7gcl8ULzfHxBKAHj56rUdipWZt9zhFrCryNL
lBZLbY5W7BEtD4ucZRSCxoz2JG0YnYXZV9AQjmVaqRPy0uz18CaYmcvpZLFwKxY7RZuOjA3ln5An
KYWauXza5n9fgnjovWnXntyeeKPi5Fsre12V+f66HgEqC37tX2zN5y6+APkLJ5TpolgVba7jbAdS
8G54rn2pUTk40Fwv6Nn8hhe3bn6tLqL4JooGbIlJtdetw7CzqAsznsXKuVqrv0+aeyQxOv06bFpv
qV5fBJl7aQdSgjcDjkxRNZKVgrSLrpr3o/YbmNfixwqHnqalTMjWfo0eqr+aU0okdbGnpF5cN9NB
+f5mnjmbz/d1LyB9WDesx8JxilF38xitQ05OKvnLl1ToEGjdFO03NIWLvkYzV/NmLkatDdKauv1W
jN0VSGDAPzOrV9JXBJYz+HQjcvJplTPUSbmYLfu/+4/FvGrTxOO1IWkIPcbwHMxNJeat1560fr/2
T62QXucaPvoO3aO/cjxgGQXeNy3ufoFUaf2GGoKR5J1STWxzhgp6WTJIyNobGXKhF6CKrSH8qjb6
8F9CNnvOskU0xzHKabp19gmUTfYfySOQv4wHxKZw5VXhwl7fUNmhBtBzwy+p9BBUlTRTj7uIl/8h
NCT6GBbap9Ti6EhuZhZHB8C1+LVAqoruif0xDKhPXw0NfbHcs8BT4grxo0n+FvqXMjBtDQ2gH+Z/
gFxQD8T+TSiw5amLSMhZLFicAlZggENNe1qd3h2nQXoeu1NbSXS0ky9I9IYv/EXluTOh65EYxhp2
atrK8+8m2HQMg5piY2NbqS9u9/I44gxFYosp6ACRDEy3+0yJX/VwiDO2/FFAqVl1vhyUnoNAQrvc
cPwyIXFZ/GyTgMqtExEZ+lr5ruso7biRfHC45gq7tkOzn/QwqDL90Fogqsfo/0U+l7Mbv1qDhgLm
4pTPA7AbGJvAqHAtc6s7WPyo1ioAhrG3AGap1nGQXxT+AGNSTjMxMashHzlTivNo1TVVK5ll9Oeq
TKAf38aSOV0mbOQ+iUakjELtAll08qmHN9jSoA83d95LsqWcLabxxTrNITgEm2hG6ej5Pl5wpFzB
lcpMf52/rRU8fJticdiM1/JoS1sUWr9hKn8j4iY8O9mqlL3xwJ3ayt+c7PtBi6/Rz/lnpdIilMS+
DsxdO+PtsnylmZqvl4A4InP8bEelVwnVSg+gRodfEHjqR79ZGl/av5p5YsJASnrf9ySfqwuRCtCO
EKnX7dOlTqVomhA5Rs7WCc93B8tmTrxZahGwKiSGSSZYQz3gcgzWqzFN/Fg7jNwf9owyUfQMRUlz
ty6WiqlnK9whBTxb2EGfNgN7eye0OmuZTjuNlnKo/fprX1976AgTdvoRNVu8tZZhaeA1zlh/HDfe
kHF8jnRPIkQ+rNqshc3LOaY+6iiXRpyur1eyhbTzKpc6CQHLYVr8/5Vi71DNC3VLst8V1u3x3wDx
z4iUEZECTdeOcZJvpflffk0+M0d6tQz/M6rE+OBaexMZMACvZpBZdL5J8W9OdboCw2NL9Z451m1P
mwDDpaMbi9L4VeLZSdEGlnwpS/8bkspxr7JgM8KPo1f0bF6spnofcJsbust5bbIDbHjfPInewng7
7JGeTeEs8MIIIjxcrgB0Yvg05PbVPA+N1qe12G47tly692bwrrFRPYos8O6Xy3jhtcy73yV6BXG1
OGHN1bbpJ2scTIqGrn6otdzsDjdhZ/BOMec9DUcruzjaYJ6pSAYSnOxMRE69yPEH8nxU2+aLauGp
Yv5ZVTOusoG0WjWcXk8y+XRoo2XVAc+y11Sz/cUM3P4Umo56/yixjIbbAgfO8+7sal1EVmiiglOD
K8cFN1G9KBXtOOPA1ufSZAsc7zdidK+Bwhk6F7a7M6PM9uFuzagiAzJe93FlZzyPsb5bZOO/WUFV
23tFylEr4rXFYEpfPVjYTm8aFDFEPgantLn8kns6oa9B8nzim0rNKsZkwt7nXXyj8e0XpyuwwWk9
gyyvFBEPYYl9wuuwDIhW2uYRd61eF1c646PvPvxikpJ/LZaDEzMsMuE4LYWuGhoEdO1UQJaQwyFK
PYPpOcIdFG+HhpUHimPvTFtFMvxqxLlRj7TQDlZU0lbh7UnWgtHiW0STzWHJJ11pJx2GLhnAYdFm
QPHKtJRv4+23kMfftsJWALXGR2L4NzmRahu3+5rd4vUGjDHPkjdD729JGwpsLbFJIz2kqsRYXmC1
TEYVY0XPopwkhU/hRtwiOILu3FuZ6X18BEZxKJja6Nea+OGBanL4EN3U9qPTMt2rG+u005nRfHW8
784PQ93SLleG21zE5UNBn4cwhIaoHL37Ow9+Sog0Y4yCgRJkNZUIA6h6s3YhYJClvTSidsYN80s/
OcuG6rIYNmwECdLvkiWAN96ZbQV7lFvs8SK+NesN0OGrFj7yeD4cKJjHsK8yeinYwHjzoZW+1acp
eeQpnowtjkuBgA1xpuen3oapJheTZzQAlLwHEgRMjSQg7/WvkdWCXEls3q5PaIHicmPhSZa9J22m
q2GhnZqwAlJ7VYojy/Aidxn32KBsQeBftKt6HHwG+Rxjr1W0+RbjjSwvB/JmBeWFx0gKXp1FgZHI
xoINuJlk0lXZ+zvB9rMAdis6N59NJDUbcxOc0nt1/ZrP3+EXSTw3N9+2/gaMSWXaHjn79qFvKc/e
d6gXgZyy8R3R0fvhMhmCX3w/6VvNNHCq914mnqNOuq2hfKIeIucthM28mwqs77uREc86Gjn04eOv
llxdBsMLKEu5kgD9x2Y1bSdwXFsF4PV2wCoqA9JKLKul1zyU5dt1Oks8sJfcQqODjfYlUeKfy/M+
ZaQsrtnafOMSD97NCGhoDdtTPJ0Rvpj3gmqQQcjnUCbP/2DqepBZ4eVpqkCMDSL0kLLmSy6DFOou
nze+5JacZifLuymjtnsY9C14V+fDkAXUI7IuRnECn5RUX7Yh6x0DkJZvDo7OS/KUP16ngqYFKf5d
K8eDZI2q+yCPmtJpqIUYEYxHw0ZEF4eTaMJ86RqHFJU6Hy6OQU7GRGnShTDtHE8iph6n5WMGhOYh
aMxdHi89B67N3ZYFpYp6Y0oka0NbwNCANHTk7spZo2GrvY1e9aEANt3Od8iUh3UjMeyFbZmnQOkx
F1gKC+Jl1ANlm6w5lv66ZHxyHc0NLgP8s5jFRfRz9j8fUmlGEpn+KnQFYgUb8rwwovUQhJn8U0AX
1UhP/0uHUPDHyR2H/XltE4ALtsI7sxE8LsOsXd4luK6MNVuUafh8MPn1npnvsQh0FwDWdYoLEXyE
m8sUul+E3VRj2XJ4tWkvfHIMs8E9yqRvZL+k3hH5RAPLERqkAJFSfxLg3VJUm73GO8/krz9nnxsX
ChRQcwvMJSaAJOmDCR46+mf7xfkyMEchgBzKVCnl766JTRnUp09zUACuM58gBQDM42t3cdwRj3ec
gmlJGUT6Bq5rAhb3dJmT5M77vt70VzokyDEHRguBwWAZaWSbMkDqTE8F7Vn3i59t+HcpMn2rJh7X
gMic9+oje8olY/3Jri8ug5xCgFAwxpkVH5JhlBVXTVVQufTuImj4MEb/u3pzeWxWekVgbM0+RmIp
20x5KTT7dANsftT8LlLnRbcwUXM7WX97fT5BmO4f5uSe/YyBCWQ1wzOFNa3IKZ/n/2iMgxmnCRbY
cr2eJcmnxveY6CmdrUe7OgqXC1CR9o2DZ8nNz/9Ka6MN+9NcGBjMF3+TvSFVBvtw9eU8byGtAwDZ
UyXc/Wd/gxS+42XLKcEqYgK7Hg/vb9l/YQSnVuehDZExrRxCXO3+qw8HZnc1S9UZJErTJJ2teqxi
3tEbWstg+xefpkkVec4qWdgUU4dismtkvSygMiajnBaK6Tj9/89WGwS/EtUQxQSrzRQDzbFRKH77
aHMSG9IZZ5qDoA4GMInpr8kVyBxaqkqJIRmYq8C3kEHRUo2RH9OsZywh5Q0ht6kd7CA95HTvUo9A
b7DEK3NzXbjK8rxqNmGxPh1Nejdd/H7qVW8hMpLPQQv0UPHnRoRUX7A35JZpZ4uVWjv14iM0625x
4IWV5cV6Wp3mdKISEaSgGSW921ziXk+iKOtP+i8oXzT98AYGgqJwJkA5fyoMwM036bOfCI7giYMt
MGg4X3eiGwVThDifnBI2HHfmwgFLOlC4e8Ad6U2W+/1TfZhyCpPz4z5mYVL5K+15g3Vwa3htTB59
R995aFbTpDOJzRmqxur1goX+gWTFofZ/L0I/LVWP2L7OhNLABj45E+dFXoGPRnAdBm3uPu1DjzYF
lZE9buDqs49Mr/SG91H2LUzxH5DehRBLx23MyaMVlFpqG4jC4APPKAUzvLgoAgahnL8/+hHmYOtz
wQ3ulxDBelHapwYtAmQhH0d8EMJ/4BwdHVv4Ue32IGVStz47zRRgQoVLhOELsfsSHIfraB02pBSB
FCQprrdNqgcJh/GVHVraBvo21m+dMrkNZQ+6D/z7t33ilJHIk0fL/VM/oliYKKqjUpdHebks8RxX
qNLiPzYQsSs4NsA7BmWjK69VBka+uocg/29+o6JZ1onQPDXvPg4jaIzm/mbKx5rYmoYPukjSdDDI
rqbaVyI3lnTgGTiA1SB/+PDlSNB6+cldxEtDiwYwGPLbBkzwGYXYHshSIKpToKz/zoYtOC3TG/9s
5xUNXeiLZkMnIvNAOMtwUPFf0SQszbhzkSzRaoJ7NjoknYXni8469IgX+xWIMLfYDXbEl6mP3NfL
RRu8kiFgwRQriRFvYLSDLeIeSGMh04eZDa0MqvzaTDv3HbZxESij557c3smPknDIjyN8b7REpJCg
EqXq18/dJ2lRMg1j+/O+MccgdOlGQvRRix9shL6GFPs5TeQIA0Et2HBvd2E1a3/9yDkvcA7YN8kn
C772G7hTdZSSrnKwWShxdb0LnGolsF/ekIzjHN+WOYdmDGPxV+fSS/GZLSgMLbFP8wHpLJ0gtSLP
ogjdrcojxmCErhIZWYK/6WqnBBJf6bo7TQ6fbfaza0Mm0oSJmF29KovkwlZv+y61E6j4XdSWuKz9
29s9FsNNm09wVBjV3HnrxYzhi4kPRVmkj5tIJazBmTNY9l2+OeZi1DJiADXk9d3gLeIQMyLdElkq
SdqCirMQ9U0uQQ+IF+r9GyNFKsDQ3mghq5vOyODmJkdpWrF+Bq3XZ5zznIhFZcKpl14KeLqZxRgN
yxINtl9WI/4OebE/ZA4UkYc9kFpeU45rUAsqQwbMglyb2Y8qL49Bm+2FENXO/coRcjUTj/Dh0O/8
qvlS/XwaaRHQV6tunLqPInBXlLakinXqq97wZw3NSJDhueWmEuRB2QXdTPOee91uAXzWS+G/crcv
eAhYo9pFFDCMoE4oAyjK1t+YEKRPTgHYfmBSL2RhFxUa5SEjy1P0c4V1Y0FylPNB36aPQlWX52Ds
jiOcFnmfLpkt5Jqpppow/oD9wLnTPFYKFZ9vrPHhKgf61K2peIAwRl/1BFaSPiY9Ob5MbI9Y85E2
rP3F5iYezxzeh0RmLVxSVbmnTQEr2kpWLxVs6Eb+ggdYTHY/81nhobA4t6PaBr7LL5bwhS/Ch4f3
1y3mkJTHfRqhEQ4+ZOG9wnCt92Pf1Wnz5iVi3ZhohmM7SGH30MS+ZYSzNZzkFAebEI7faBYhUGR+
aGmyKMhAvqFQlGUzEVoFnvI6xmil/qYuqWt+d/gRa0cS05c+pRxkNMCWl11m0kBsvVCajsIOl8yT
g62SmqTP//GCiinBLLuNkTLJyX+i6b9VwB9H9SRazDKjPZzXLiEFVaHi6FSphY0MDEpxxjnFwKcs
MXCx/B4eZ+wBpkkTwqkzuHQsos+e96QqfEXeRj39ZN2yujRrJBgZPRKMtapAWEufZb5nc+TTq8L2
nvXkUnTvzMx1rdIvGpBIsaYueXlkSEkaHDhdyq97jtrVPhdeD48w5tLRA93clOO/UzLXMvjwFHiN
IznFOjCsRB1p50uNFIs3/AMpDp/Oz1BSSlWyJ2d3Siz++ABJWdx2ekUCIOgPxeC4dez6buYO04JW
M7q8YlPX319PWC9Bk2W7FpAlA5HJ8Zf9DUK+fJR8HTqtV1kKqyTnYl+2kSzVsAZTl06Um4lr8pad
I6s/4VJ8U5CBfTaKSAZ2JJ7PWNcDsIfnNPeNYphz8bsWyxjQtf6HNloZ/Q0blYDOKbvKvO2vOFXR
PoAI72wpXdw00NEwck8kYBAet+PLI+eEZZg2MVwBIA5Qh92GX4ICe1p2JtaOL2xyplMOVNgboTab
DYxldFFj7Bzj7JrbE3fo3ycymkl9v0kZHlEB4AmhBGlWZV5sXJgftN3qOhZ1zWTr6HbJgisF7Fx6
h5BFIh8uiUfo966G9872SkvKS1dy8oQM7qo9kI/hhLTWOB/mARJ5ElmFMzWE80jnk+TxsgC2I7FL
88hbLs7z99t/qgS4e/XrRfpvHlPI/Czlizl/mXY55TlXClzpbhO8gEnnvVujCNAsrSddStFzwR1B
zp0w+iM3oynnsRbZQHNhsaeVIdNJ5+wBFwWcIcbi9LWfPFk46xs1iTg/YqmuSI3zi3Q92IKeZDpG
2DHpyGSzhW+fIWruV2wZNag8bGB3Tpw+57LOp4IlLkAwnsCCCr7RvYnphNM57oTGC5MxYoFr3CEh
zE0kek5VWE9QIyOgtwoNytvC9wufIrW+IxNpaebCo//iy9LBulzgA8sjJZLDiIfo5GT7U38o96us
vkC15X+4BS1C4ovv/GNR0PID3yhfFLjYfe8F8lr5pTHnD88VVXU4/rfzN2+4xs8d77nxY/oBGIn9
Fsa1xGxyJi0i33TPXumyHkv27Wpbyj0pPVZ1Nq2WdbpC5ZPkAV/wUdkZT7Zz0vMb7lB625htyVc6
5GFR25GxnD8hhfcvHDXeDScxmUyYKdNd+F715odAHmThDZH+PJSadOmh170bcVkA1qZxKySw6HNl
W+ekbo1zEG88AJwFBm7LDp52cWu900YEs/ZzeBo280e4t2SWwia+gCks2JcQvAJ8LDhWwe9ey1Ky
ccRgdQ3v3AY1nN/njaxRZLjRolxav95j87ImgaYQKxAxeBlblQMMbSAUOj7ifw/t6QZo62iWQxwF
8Vzw0eyOsyvlyuOCFzAiWOdoOE0Y2C6+Fm0JhKcu0FfH5Kr9UhINOQRU5VKMfECgdAMniyJnaxzK
qOTyFjLtSRQobdDo44lJH7kRqfSaL8vLQGDgkiOkAIAGks4y3OT30i8sg9Nab6oxKqe86lAmd/sp
bkebiFI3RPSKWPTnvxgPAktcDoh8mnvtHhTTeLMl2apgiqvEajLXjtF+JH2SFUL9ShzTeOms1OWX
tL+DnRseDFNv+5XWJLX9fDGjQcuseXS6/lM4DWaeNLVXYFOxnVz/0SqMJb9SUwP5TIguFakPfqVs
rn6INLFhySUGiwmzXoQ8Tss7D6ALGPNQDF+PSxbgAxsiznvzwG4bN3qNH8aEl9O0A/1mk1l/IE3R
DWHlXeowTeT3em+mAjncE8fjaAhwvHJwcBGlfZnPcD4+g4bCD4Fz5LqTgyxpVIW3N8r1ovNK0WUj
kn+Ii5t45fy2B+O4zXdaOie8yw7W7kuPElJgOCyJIEnUI9PhRA+MXD466ZdO2qTv7mC+I2iRxNKS
KR+DhmgsZU0iI/YuLrekdiqh2AjWKI8FVbS/ZTl3llSSv1RaQUWFeWBRXV6Jb3pLqQb9Ib7ThEPy
1XPu8PB0Ri6WB+ALs99AsoveWZPQB8Q30j+MKLy2JslJwtYBV/YyA1YTIyA/Y4HfEKdBj4VSc6P7
C2RRTY6eL3OGdC7r3cDJaul8vTzvk9HBbtFGQY3iHHwE0j89blZN/Z6xo1zIXRdkhC82JtQEkir9
hYL+4DBX6771lBTrbfTG4TOT3eFiCBVhUP7TeYbxLBpp4HDgFWZ9IXOwIAnQk7+N0Upz3ZxBuDUG
oYY+TyBGp2cutj7MjABj1/Obf6P5uZaCU7q2R0YUfINOb3QaXAFB8hPWtCmu9G0TWyUSHC73wJoW
vq4GiVor5x7hqiy6TKK8bQWQhCkjpOgFk1MGtpbMJlC91VWG7Uir4vvC66PtlyHiham19z9yvYQj
lRZb5zDj1umRDk7jPQEKAbPC3CZCBgVeGakfoggpRVOY2NYpkpK6+RO+IW0A4YroPvXcwdJcNLnr
PfTFbpyln4i5ddXMfBv62u1mY7/2CxYdMUu9fYaifrUGOV7mEXLmsFq7APV+LKoLTRN9cqZxW++p
VpmAcOR1pBU0E2fO+jifjo2AS9YtbGQloBqV4uLUUJqhtlgXzerePHpFzSgA9AlMGScAOk8i3Au/
AIEQsOJqCGsWjDD/6ikK3sKIuzWHPFjjPKiyGiA3Uxgt4mdkJ1mmf9jxsvJHa80pEnx9PAC6YQKm
LriVFjDuWN22uXHduw/L/X0PliGCrmhjpPuLK7UL2hgSg1LmvIGTuIqG6/+nHtyon5v8vbMIjdmT
TfaXQCg6HuelbWKyB3pEyoywL8lAK2s87BMrVIRQlRCvt/S3DbvWyiELCZTbdKA4X+nKXvHqjFms
C1t9m6PWvvbcMaD7/WNw8DtzsDsUOTiLaR/A7fgShj0aTAjlGF7ONcUnLNzM0ic+f4IMQCLr/nTO
zHNlHvswXybR74t1hTwlcKpVYtLn9I54EiEFkGiPNJIKDFVeYvZRnjvcscGmpn8wUveLydMlhvaQ
LFoT0gSZETim3q8DuuSH+/yi/gYqYD83WcATHGonQBQ0otnIedEKJpWK4f2UenT6jAuv3mEz8csV
fpfCKl24QkHWWxQTQrJNFYTfv+Pu/gqmORshPR9eYgUnxFJAHKWcCgXtW/DHhEshDobC1Njtocg6
U6cAfboUkCdhQU8GRGBVKfGrIHMfu8UpG+aUUuodBX/g3sCyi5jM09USWgLwbaK/lFPfKTXlqDxv
1l4dW1scObz8jXZKxpXmryA43XToLs10gJsrKVTkMUnzorK809fJnIIt7h4Okeq3zmPKdIIoaJfJ
zx9rvPFLYDNTWDoplf4zLWLRJIlSZrMshyjLWYoG7ZOsRDvnG05hdRSim3sMVelSqeKuqnkWsVR8
QS/Swcd0u0UgGlDoSjvcHClKgaNCuMOc2nzBe4LVYaiLFVox09TsYf/QSoHSRuff44SVYX5igSLi
SfO9MCt/24waC+4U8N4rTzkRf3HT5yLkX84Ay4yl/QjgqrXMyAOFhBJBRucNJmY0bVoVn1hb7zrO
a2iGwdyheSJi6JlUf2pXQGLachxtBYwJDZKoCxMyuNlUesOQ6H3VFY6b1M6hwM1mG+5aCKayWDH0
OD75HTZeRMEoyg5h4/04TmqPdhlF//Bd4F33LFJoIjjw+w/KXy46yyupsjX/PfRzafs5GZeBv+6j
C3HdmY0Gjtz0BXQ9Z2h130aCS2pQ6eW0hx6ppvgxAipDPbMQsVJRGqPGF4Lcyjw/H+DU3LgRVmiy
WnBrqehYKROFs2UTNGFgIeqKurtJlNKVjMpLPzNgQtGJpK1Aewk/B+ax7xV2cmCT6heBmuraQmmW
EaeTxiT7Lpuq3t/3Y1IpNWGnQ2UR0jmUYSNHLBhtJ6jQv64kENYIXKPxbHoNvnUs3PaXdRURrKao
5DpiQHqXgpSP6THQUNtpxYKrODbMFo0NHzwvGT0zE945mPE7GgSjzlkfS7opSH/ER+zuSnf18Iyc
Hmgm+Oz37mWyUdtdSPRmMbxthUTSS4Pg6HlT2QNMPVqIlQNoFFeuBQt6Rt3e+XBb/YrQPBIDxaZL
DER4nulK9twSWVwnuOywtGBryjWQhO0YP3vbUVdPfJfgve+qs+MZX7pL3kf3ebZyhU6y3pZi5s+I
Xms4SiwJN65vY7uz9CMcm8uSWbNKpVkmc3tMSGRRnIyByKBFOqValni02jzuUvZ00ZbzjcOOMjjv
8EuXDDTJPRbGpD8896ID5dOljKxsX0sF803IQklqx8oCSsBZoNYpGLOAjpvhkF0YDFfU5O5f1NJh
IQXhuxkYu1GVMfAYVRKnJ5/69kE99qacsmmuRFP/AMoaZ9yx7Eoar5/B3y9fRacWmkvYA38oFT1s
8QZVy3Apxu31fu9pAwoLpPiLLcCO7Hw7Ca3WHgd5u4PzER6rQN3prHSmG4vyN/6jsHTUwQtCJcrn
JA3c4cKcS64z8d1faXvEO3WnE93qQJ8TtC67CmBP6HuZYj7Z51vW1q6dg/DErzT4lJoQ2FslKBFl
Uq1sc0x0ZWXBDkALMThvEixy5dcrP9coClGpturMkCp6Lm6rlHknj73dymeuyKBKmuXru+rtwyhk
iIM1oXQuksNDb0xTkTRrLcLTBXbaCR/gmyFGCHbMHnaVqOwUQ1LFqgHMYunuotE4Qy+m58e/nG+n
uYvsPNG6+Unr5UqzNiw7do2V9cxWUhbsNP93/Z5duolC8K4XCSHgG5JPX70/zWuYqFGK8pX/IPys
wjViXKb7EsjienbB4Hbj572E8cKABlKKYWOPgpAUYvzDqMZK0qXyQyROhy5tU6qjyLmRPx85mpIU
QNkyoAH1L7c7ugDagTV08YDWxQ7nO6x6ThpkZoi7JfP+FORpn8RmKCLwajkSjqqZIm0uWmH9PGU9
Vnv8EMNCFyjDJm9Kub28/pCLkPRto77735eSBwrnbnrebqcvnQFZnL2Om6W2/Z0btJ5X2MeDdqZa
2YE9wO5xvGshT8ohlcZTEdFEQ/3c11JO09pBbKBPHXtfK3P46L7lFvVpW60sT9sVgdDMt5Txo/D3
7bmhP6CSChnHTQ5mQdpJSOp9B9q1qVDj37L9MWXQRgr2nZ9AfImbG2qZd/Xmt39Wms/EOvUWnPdN
fsc/0z1q95TYxyFA/QtbhjOyzir+WGwQgjtIURLceG0xkZ+AEUzaBK/G7Cwub2xOGmppUFp7eYvY
oJEBOvAIqxYvRtrobbANeIra8s2VQspDNn3yuGMdwpx+iydqxUqjFH2+bfFwkbIDiHDCMbxmyxfP
vQfwnaGHW0SSP6qEFZlbfgU5Zem/mbrrXp53jLs0SxepnPan0WRqqUAgSvUwNXZbRMd9OWXcthRk
nrAFuh7IEiZqlxZ+KrLy2fhtnfc3uu4FQLZ7ipQa2cPd+KGpYynqhCuavvV9AnwuJ+Ri7IUJUQG/
/qy0+6belLZDKQx1Ntnjupyy3BuVZs/khyMrbHAZEEQeRiXRq6roeJjzuytbkukZmYUPJ6jnZs7s
mZOHfoRX49TjYCj86KLLZuBNbu8dBdtXQRpXrxwP0LFysHbzDUttWuBcmIwfXu3G1DCXZ/psIWst
AZnL2kiCFbY1v76qT3g7HkNP+5sQGMSQfRAVTpxm110Da0p/vMUs/LmWz4j+kgX/vI7XoUeXFce3
NwvBoW3QhPXj4jVewPGYK+t/rtsOVliDD2K6RfvpBrGle2B6QCdBkW8VyvXdfhOqD9fOpFIoL/0J
8xu9/NxnIpHYsisDVRDK0CU51m5hlbQirvBT+QcdRau0kNA51WxRClSovZNX8CRFMBMef0tucOYL
40Uha+k3WwWOp+lEkSgVEul1nfTjATfp0SRxhNvWecPHQYwu1rX42aixZVZtq9DHsVucZorS6zxl
dBwQuozlInjy2tJtxl/stUfH/JYgzqC0TEtxmM/7U6LH54UtnhvtHmAJqd77yCj9/aH+sZiKjhNo
bMjQw3R5MESFyu5jfWiPb0WS5cqeGUC1aajoaE5lUJh7PBzec3Ann+TQO/QbD4jPDphQHvyjIQlI
FkBzfvEViVAdszZSpB1A4meq/zmsT5jtBOQ//ZYnBC/txW6uNZXEqnU8dLmP9jfDlKNqJVR1s78x
a/ExYcQMu1CbOL6Zyw0387wWqDM8M1rpszTi/F8OApt9PP4Q9S3pQeWGW/WvfN4IlXtcPnVHJIFh
2B/vP5ldfrorGursrvGFbLoW9CVhAorbc63mewD7O/7rNB0r5D1NsSw/6ULxf335dEg+N1M+K51U
P0g3M7KcinfFvwGcY3R3XYdUbtTgcMFXfStus8txxWpiT/2dAOpw/iUMNUAXNwy4nS8Q85HB2Kh+
QBk6jJtTG35bY8DFlbboGS2Leht8tiePrx500Phm/ckd2qGqPnuT2JMm8WVlhsbB385z8qKl6xRs
V6Ei5BkyyPrI0uPUCK4d9kaH7wL+xe1CcLhEgA8Yyc1LZnJ0+6A0UygKTA0UaNNlzGIBNPgTI5U3
AN0gx6122EeYX1fqka+aB+5aK86c2r9IHdNDIl0KpLwiT0Pj1cVr/wmh/cFekT9phQpq5JFPrcPy
pTI0C9XgjISO+uBZohhAi7PyyO1r/PnsVnoGXzbczeinWjx5uJ4N28+j62CuAwXVcKj8PA2Dey2z
OehX4xi5aHlsYi1VCR6lN/afy0cXdnvd/2wfkqVfDQEAIpIWtTOF5EQYJofSRzi0iD/zMcSls2T0
jb4eZWQ0lwcfoA9xeN9URIaNsmq0eELK5cIRySRh52iFkwbBTFDJb4d2fVHE5XU2x87xVBNkZYC3
Cahb7LcNkKCb3rnp2pBG5LLcsIZETHvJfoXKXf1dXULKCYNrfeWeQMfd6u1vJauulC4mJgY+kpLa
5FFNCjYWktaUS1z8Bi3vQdWRQ9HLJo+CHwYmXtDVBgYQrhZdiS0881J7IWSzZWCSBebqNmfdJapt
0j30+fPbl6n8ZnRuBlEBuv6swsw0HlsGnQTAXhcdSB+mFB28stldanbQP7i3TSdmfwGtqILzjhsE
5J3ZDEfuYXI9FoXQ7u0xeSAjN2EwqlhVQwW/9vgI0BzmI/gaOmTgjM0346VrOm2RAnWf7kFUYUVP
8Uci9ScK9trR0exX9zWym1s0wrBMPh8W+T/o4hMBWkq0RCFBi605WA+jauC2EdabwcELA1uJKoRy
rO5oyWykCMTKPBKaoH8c5ViR3/tKrXEoaEU+aCpJgB2xQxQqvRuzjrLEjLTtv9PSrHIS8gj09XEb
nKcawhgHKItxnyns8j3s/Fg9Fxvwqgyz9AHYKzlne773EgvHMTQiqaia6ydYO2DwICVwWDr1lscB
gUWuM2T5I/kkWQCygnwaSUgu0zxnQLAuxNexLlLhM4hYaiuohurrkuWHKe0A+0iPLa1kDK3rj95U
eoP3I6M/yTesczKqeHNluD2eLlTIbql4F70nwJuLJIQlzRgEqvhrA+wkrlGu5eArOxGHDeBnwuvP
K07ZUizlg16p3hx/g24XrbX2SxUgXk1YcmFenVqUXrC8NoZZEEH2Z+5/Uk7JlFhKQgsEoqKx6wzs
IB6jssH0yVUfwocMaO/Fuq4glsEkkHEcaue+Tz0sX5aWxuZAinTlKhPa/KH0kwH2uTrbdN3gFym7
BCXWDWBSKtb/4cgybdkUvDlXVDlPFrCs6WuZ7XPZEmIR9CB5ynJ6QvuW7IwI4C1AqRDdrrKi6r/n
k20Ljv3joxhWSqWwo+rudlw29Iex9ILik1jrWOmRUUjirpwWO126f2KaCNtrnz3F+vPRW4JISqHu
M4Xgrvz951ZDpu4JiI5kul1oWMo+b/E2dzb11E9qbQI/meN3Zda9MII6/npWBU+YlChtqeRwZALs
9888jsLYb1Q6twc+Z5WoMAw14ngvx/gKO+du3cItI+juHnapq1m0Ya0EJxT1Fa4S1rf8uV78URq0
focydW2Z81OIq6yLr6EkCcR2eazbiW1iPCacXoweLRI2+V/6kEuzCF82Tz3loM2wjAotY4aHrtyI
qcoFNWM9xZKtE1MqF0x1nZfVV0rwdL9UQDpvuRaLK7hd4331r23B5+lRO7TF3bSHp/JsFGLhBLO5
Wops02aO2hoZSVz3/x2GIgdA2i1uqwPDVw77akN5uTkDX0ga1AvqOez3MotPppJPxYs68LLmuXe7
UnWGXck2r9qfpPrzVuFrgRJwvNRBKeU/S8PkBuHefBP+2N2FE22saZGqWd2N9X8lUY7PzzUHCI83
chavdZnJQINsbYHk7/bfDOM0f89pC9PkWWmmS5T5Nt37CSn8r2dtGmsjQHW8KsULRRiVs/s38O50
BWnvhQ8SE5iCZsH+WdYLWhqKYnFRFwL2cTOPCj+4ij6v4LinIxPubQsM7YljxakO4rBSaDWJGJge
FdwJFrr1pFhSnUvLbrYLTAaR57+5DYoOucTiD3uAhL+873LGy56Uayz0cTbL+tq1ulBO05y8JlTn
3cCgHr3pvZvSUkCfjfGsq1EIkQdd8NEXg+tzTwktRo7J86nXjstOYUkzLHsPXxrTQJNDFLrdnl/x
Yyuks5cVdmHxrkib3TnRdYZVQ3lHTY7slUyEGTLQdV8hx03yzh/mMZiA6RScdMl3qiae29R1GC/e
kXD2HgWM83zOsbO3gJvB8Uj352P/rVK0+z+if203mLjCCkVmD517ynn2qt8JE26AeWLvf/8UeLoM
h9shJk3DWRtG0qwc7qfuV4ZFbwZjPBy8e4mShl+UspmELVygbEapMvhUGytgDF9JQEZMD5GKId1Z
0T2kddhUU7jwt2tQkPH3XpW+En1qEU9XMpiBpLIpNsjdZQ7cvgCz8s37H29yoNTdnDgVJU8vTZMO
vvlxnWq9SSacVYAIjD1jo5s3dOQXtflFakF8JLPCD0nUMAQ8+xmlw2ymIxzzTmvgh5V1otAAs2ny
G11QaPJNaYrYP2Eaic8nKrxgj4UpOemDhRQcRPvUO/H0EPU2LcHPdzNG7FPL774ACQzNAubE9sS7
TEc3rxD0953ffAnLrF4n/aIphECSjXDVZKVdZH38NcuypT2qLQB/q37JLgzgrMCXqY1Xj6J696Yj
S511DEkdaCjCgYUxef279wyiM/+cF2398gEYLyc3oBx/b1xMmxhJvJVjC+dw3/AEwu8ttjCu2VsY
NLOHhc1/QsgJvr+42hpry3FGyLqvvgH4NyQ0YLIg7m8zDuIYpfr69YP01dn7PtE7mxbfMYQefKod
E2ZFj9HZr8XODnlK9TqFqaB6jl2n/KFvRx9EnHFBG9EAdcRcFCg5VhEdvUeAdPpaibwsWK+3R/Om
ukxdHUF9nA36fRez5mkzdCgz7s1C5IhbeLjpp2SW9v2D5ux3BSv89Ce+4YP1TOon1vVw8eRwsk2c
uPSdCJ6m7FZM0OY+UKu5prZKwL4G1DkKSVmFLiAfZlbIl2VrJiX5E6R8ZNp34AGJN28RadWViyCN
gpiLDzrCIzfg4rYAoLBX/7eXcG2Gdsp5H8PCZuuoe86bZGnfKf3FK+8m0Fsgla2CczcoGAaLtn/h
YGZUpsre0yme0M27cy05J+b02aemv1X57M2rP4hIH7owyhSaBJ1trjlAliD5dydw+2ZJrBmWl5N4
LLTp9vvbal/JyUXynNn7RB9PTskwXgW8RCASAAn/bRwIJzOCy5L10sZrmiKm7wKbbtI0Gs96YTBU
zcSx8De67P5qsRz+rA+JEA4SISUqJl94zvAsirX39Hadb/IzT5jwz3/6abCetwg1udoyqKSu3QtH
bf8c8QxayD+Tk2f/dR3ZL9+AG1jhhOmX34u77l6N/SqLCbLquh7kCq3Lg9FikUZlQF0A2nTmRyoR
oEZhwFt4gypc8JXr8cD+OMzm3F4O4dSXAJRdkXAEfWfmtWG3DJzCNkbdkPI3tTJgNz2wph/L7JAZ
954jjLb98Syjs1aT/fjmsSrtNr6SM8sZTgT64Ht4B2W6W2iHwahyG2EZBMudu9s/GDuyzIZHwcjG
LL6ubQtBSutMbz/g/L6Jhtpyl7q+nvQdoEzTNjWRckiNXw3G4NvjPhwJGC+IAmPXSCmNNr2NRbRP
OwZwvosQpoGRSf8RfnZQ0Aw8uGY/F/8pmOjhcs76sXqED2jHQLr8NryVOVTxpY02LP+vSvRzfUw+
J49LiKLx08UhKyTJxenXlan4+FN9Sq3huUDIHHtolfs2eD2gHZwdmBoAIsZbZQvF0/fSkcc6sMnD
THWGwDhLDDsVcYkHwVB8cVB9JKmcNKdSlCk30/KenOUG6ElrvJ9KPvgmoSBEFQyXMkyol29PLovj
7cL6krBtHJqsn79BLmx+11Wvk5JiogyiaCjVPrtP5zfX5ec24edFOHyQDwFbSIhYrYqGIpfjJHlI
BXnkrXSuS9uRqVhZDRnJBMduPzMYzaNgp1e8iwonWTRN0zgK7loQmcl6Fz2Vj2DxCw804lj8RZPT
csdLZGXMeuDN3G2BTklWWfrHXEidSzRjH0t3bKNC5NPesH2qnbJNT322Z2flxfWyE3ApIWnFX9qT
Pc1sLWmszmD1bvaKriyPef4ltAFluLiCoVeZY2q3T10caYXovNTwwOLlJUwgq5D7Tw/YGw6LLJxb
FwBjU44Bzg4NQahxuqbpjAqWnuEfqd7JFxhK9Noxpcj+AW2/+2O3WfxOKckL9qf9t9AZrAecmoJ2
at3FCObViCZ9jF/OKoyo8GQkLLDuXw+KQ6JyAggc3NBxQXF/rEuT0F75AlgpLg/qYoRAAMeM1suY
W+YU0FHpIW9vFevffIPJOeO0VS9z1EhwQJXb5BcIRrAjm1thpyJZL78wsY8tb/6UioPj23GmyMcU
cTMy0bnW7Zaypoj3t1vgro2JHiroFUVtsiY/m0vqPzsZhIYpSlTTyNYu1hNK0WobK8rUyp5AaDTA
1RH6ZhdMFYylHxfdz2tJrS7Sz3+YLNJhiPNSRUJQrqwUA2Il/iwK9baXrMkkXVeQy08fFV4Ko0qd
I5DSZffFoZPT0ywWYHoCDjjNN5AMRh3jB+ZxTH31azfo/BCf9NgZMfQmVdr11kCNb9aPo30yCyRK
WzSnyr6poL67z3ltAFfg6eKxxMh9UGpNTudVwmzECJ/fhcePpPaFln//73ifowp2QCMJ9RdOWMcF
ii2FGxQ66liVDb+vENAgVJXap0VXW5j9eugFxpYIyyC8ZKk3v6apXnFwONlF6eJG7C89CCJGc/if
pb3HajTLbJ/aVl/OlScxYn4yjz3UxWfNLvUxgGnuwTLn/n1G874IZDasXhRRJ9pZTlNovDwZEb5V
WhXVduKnnJ9xOd+bUYMTZR8fstmZs074QFZ3LdYnWLVl8zwUEOtrSUvBhIEjDgZklq1bGd3N4nTs
fd79aezxMWDhjFXE9BzevLEUfAKyy8k4QyTlz6G35ktfiStezyorV5RHq2yKaGLDBoCk/17YKTgB
O3NwmTzIW1rNd4EQg4O5AcVjzTCz5nnjN1YYLbKm8BSGedbcqq7tjaWfbfSqfWNEalBD7OozZmUa
iNrxMyKk7h7R4/cHjADRQseEtieH9wgojv+lE8z32d4gI1j8xFrGQkqMbkqC8Xc0QQaMoSQzkpNX
7kijdDcszTwFXEs2KMgVrtMAFLKjTCGfO4zebzJeLsebO7+EDhIZes/w/K+XAnqfntpE85TEMqCW
dZiLNXyq2UuQGK+vaV4iOyrjNzkb1UUPfFazHoZrKQ9rnuOykATjMGHraPj+U5sWIG0dFw4RvYuG
OBubnkHES9H8IvJFEvYS9SoeNB9VXpa4e2pO65gC40Hza4/KSquuGqk2KSiFRUiNET3Zw3n6iT9D
lYNB5ZsVfyXy3hvSdQfdpEI51hpayamGa/gG5uqNS6RtFt+qOojUf+0cxk83OPl90lB0iJuhvFh1
ACA4se/F56RoETIfJCjG8LYRkFnBOwlORvhgmHJm0SFY6X0JmQ5xkqGkTU014nPZufkDG27cevh1
ZbnV1EJhNI9Bxb14Yh+SLXcZVU/0l1SPoZR2FleD85bt3czxFrMCk2O2SE9YmGVrheY+rJj4Uqm/
kFZwoTWCHhEE3wUPHEyLpz0hju4HXKEkG2OlWRjHkODOHIqsCHUbVdMOfxPFmJVGMT3DbFZmJmKB
v/UOU2/8KTNLraK8oeIHxacWK4vk/orPHKXyI0z+/rUSRDPcYH5rJ9N9VuCNS2obp8cG62ZsjN07
cM0OdpPKBJ4WKDWRrXpoah/7JdYHModrSi0EOP4dXBSccVnN/X0EjPi/tuHDsIU4r5/djWkfST5R
w/vGyXIFJEzzTzuhgeF5SVBPhU21qOZ4iB6RULGBCOHulogOaF8mV3kpunUQ5jex5fKSX3nEc0l3
uXy0JGXqB5chcw4EEon6gHROVxRhZhhYJ17ZUcftJ4RsAmL7t5FYkYirKzBR0TQ/G4hGnBLFVlAM
I3UeH/l2YmlS4Z5Najnhmq4Db6PjzdxSkDdl5AC0XwyPFVENDgnfhiXiSJk+NHqa2/diy7btiRj4
/ZBYcVsYBs/2j61VZIcsXgfztk6Y6cRMCNp7Hl4XMmmvwP20MDb9kv0ei5Ji+POkuaWXZQ49e42a
Ct5J48Ym1rKR2PbID+VARm9EysHbScr3KjZ9AfsGzRdwzAoPL56mt6q6RvuAtSTRzM5qk676hPwV
HAKWA1ZWj7oxa2urpbbTPWn4/0Xl8OX0p66ZWkabBwI14t08mUEj0NA1ego1hiEX69MA1AHd16NM
CvcYNDySXcKANgXrAOmDtpAg73b2K/+6phEyxzp6ss0eP4nGg9yL4+wfKOF1c6oka3P64m9vmKHI
z91AGX8djSTgtcESQlkik5NIc2SKUOix0CbR6E9lypCxZcyFa74czihrT7sI4LgTnqpoqE5uMd+d
kZ5u2yhIbhNQS1fh2CkUWvWoelz7WejC8ve96n1nMihySPCTyPEmNHWB0TXaHoLtN9+jY1tlPUVM
WKA5xVpCSzqGA3gMURO+eiLs2gVtuulVWiwoYss44z7b5EuVTpa1nnYlkIAG50z02ln+/C+2SaMx
76rQW9SlofcT8Vmh4RljVXJK111n/PjlozthtiE59NtRegVTVbCs+CalQ0jjXRkwv5rVcS3I06ia
R+24eYXS/JDQAnby4AUNKFCikgEkrBkWW3v9QecHBSnhqGWkrkRxwMh2vdZ2vZ+ef5Nz96FujGI8
eKR55A9Vh8Ua+PHqIKQzqes4iklUo6ShIzFTD/HqNCM824Y4n/76J4eiokuyO4L9Wx/1wRCejvOc
gzvqXNG5bMLqYEYYpGnEVhFSwsSDnVSLER6Jtftxhek6EYFFdXoq37dV7CDCo3ItfDQQZ0IGjyh6
XZoDuM6MwN6bTrnqMhG7fk80A5i2vnspar4DTz0sIYMMG+/C8hfERlbQbSHG2lNCkaGRHB203YOE
oNOB3OmzaEqFToLl24IQZ2tRCsInxVGnBxA05MLoiEWF/a7QmKXCTCQDIJDotfIuGutBOqVwPANF
vsF+DCLWHd1rwdTAX5hx69DqRd2KhnEi6+1MMQ+mrOrHga9Cny2Kofl3wy5ghOokDg/8pJcGkinC
LQRF7wzm9rfJ2UtTd5nRm4rUT6cjwf29qNlWF/ofiE01u1BTFpV0I2FHqTLHToXLB0aLGClg015x
SNd9zFAx7ASmG2rv8Bs7Lr2pMy9w/HN+zPl9hr/uprw1BKeA8DHZicQCE9wXmhRpFmkjMSJX5SlY
ApjopdzL90ql1NvaCy8Nqv9XOvM6mkZeoistGnodkwT998xrgYJryw7Kfllc+BEviZF0auW747ct
ShGBkmTJZOndt8a/K1IbBYoF4eS5x4qr9rzVURAkq90MNXsTweZt1euPP6oXif3AIy8G3QJtPiht
5OS3z77QAx9rCXxlDjpoytykfx/D+j90SdMwclQ4pNAasfsy0mOAXxzJ5AFDpB+scndOL0Wib9Tm
0BIjWGlx2mGuxBNqPfeVLWWxfAX16ND4yjTdCbV5CIjM7tD8M583uVtcJyFCmLI7+5fU5Qqfd5rg
pDq8IRhIyf9RM3NAEytYHnsJEGfVN3YojmA1ZMD8yvg5TITgeiMG163KuiJvFfmKBOqDAYT4GUZK
ObtNOAm1AhKm1xpSKCuDaoX8WGKkBFYSED9s6OJyulH3XkqKl4PF7B15/aeOPwkyOF3PiWmiOGRi
dxDYeCVBpi0EK/rsTFPu7DnhMGHv/pI3le6pofjLcaZodjFnkrrcUVHnl9Z3UqQ9ihr88utOT1EL
Z87Tsrz25NhO9i6jTTFIzQI5xEOi7ERPT3U30B81A61+fM/QiKhoATuo03dLryiQQ/dac0UHad0z
V/+jo7nMlS+qeCffqlnSnmH1G/NuXAKgNl1UlUqiFL6e4OSRm8OMtpsaZRgkYVj19d5+xQiBnzhs
Ouiz6YFNCex+GrWvvlC9pSU2PlgNA+Lenf1mdGP+UnvLyB/cMsHrFhLkjl8KsipvOKISAm2+pSoo
sKHbEOHvWudJOTRwteMddCGv2Pwq/CcfvX94Iyk0HUCxULGIWM8/jlVhbuqCWsmlBQB8JR/dFscp
Itdl9fzKVvuAppmZu80SlMKw1lOQpFoNdHHbGYbCwD1bOuulADYBQ6xe3xdxYCIn7sTokvW3bRun
PEnqSJPhNgrtCr6DOAIFV1aNEvOgMKhKHXCzejXxBpI55wEUI7ZHpyyS9A6SolBmWAWRN9xSxgb2
mFXTGR1eb2zmoh3uj+1+Gc8GQxe4VpzO2yvTnGMvLEccVatWZWgdHL3Brr8WAwOS8gBt37XgRVYJ
D+5qh8/5pf7DQtAPBEySKy8zTuYj9BHqSS7D/WqXo2ucAfU3jtLd75VFdT6zNRW7btZgqrRgu+Br
0d1ITphaMDfmbHr7LcAZ+EfbSexU2V/uMzrer/tBkN/3ZzFuyy6NiAng+QvjMuR7JHZs5pgO6LJP
7pBmUUMnHJggmwmGUAydMsFFRfOWxbYU5mu00zi4keLl5+dwwBf0tCCmmue0rbtuclzYn98Ln5JP
+gXmh+Xz0tIhvsIwjcFQA0CYjRdanPW9WC/HDVUyG+kX/hytk1D2oi45uMjufi4QvMELWILrp7Or
SqcFLnu3SLAKS8g5chgN9em+FWotR3W1QDw8K0Ys6Y5+VV26NLsZkDSBWopyNIegbUXji2fdoNIN
7xSLRaO6mcDGdBRi2glzf8yXiflPVO0OA3GMGICO8jACpzWcktOdezWQkoM/0hm3ESo0LeNfL1i0
YBqncxsZPJo9aT9TvlzxTOA4XonL1MFjo1Qg5dngaxATzM/BgTwe2mSAX5Io3wHL6UExKEhkoLFb
wtd7ZuUnPyojFZBAlpeCUWQLPbJQhb0CbFkjxfT03a7xCG7fbW3jBPpeer/Cshsrj4bz718DCyOp
aQ/31V/V9Pp/Xb15c47C6yrW/opn7xEhZqf3H/QXAcUM+ZHv+m7W3DMY0Rw1P1iiGj0ej/7tzpJy
nG11lQBcBF+7CLgJRYrd9VQaKqrP1GvYbaknWuOKR3D6ixIrty0V7wxbYRi2dFmRpIAxv2YnhMRM
U7f7+F3xir5PdRVixpb0r2dt3JVjzAklExK/QFGAmOC0/3CYqt7kczQFFwSjR98JKIoTP/zzRJYh
7KGUTsRCw3VgyrMpFv887fd4pXys13cICpcsZb/HTFO+ft4HCe/vOOaI6PPhqrHBF5P1g+xr8rOb
SInie1EfM36ENcvmwQXee/KbCCCQzn7Rmdb+OVS8FRoxTC6xl4qYvGkmd2XyeTOHA6vlG6Dgv4c9
bi6sSWhBDar8Va+LWG298ao5ddzF/Nk4K3qyCDi3MYUO2VmYDw/AQ4UHbbOyw3lNuGMQ8HIOUovA
8fvKuzfatBP4Ii8aDpKdlnpNcHoxJiYuAAeuFaUdLRI7FJDxfKMRVt2vJOJZzuwTxDdSrY7fYa52
sGUdef2yVf3p4LPYk7qqbL3w4TWkN4mZ2bWPA5hxXV0Z8+W470Z/A7TzzKJ5RzITJNPduZRwD7yF
nsx/LpeXuJzNaVTDrwjkoTnVPlJF+dh5BeYv5sRI5Pe2dXn6GDjRS4rYyaTBSgL6QYkHXnlCmXF0
53/YevGall7+tF721N1b0JBdeqm+Ta6z6k3PlUO0KxGHqD7O6VCm6EXA436hEzHiZU3IQbD1tCtJ
3rd+/bvokGl4iCasFp3S1UMfdDAY3s0bsmoI4rFlW7iiS5ZQy24DybYbn9fgcN+W8uf/Hxu2VNYs
J/1XUYeEH3VGeSolQqZ/vWm5ddJZXVsrsszEZbcQSHM1Le9WAFXaBwiv1DFulC77XDKLlLKl1EO6
zAZhb94rBBk3cRdcnwEfb72d5loDEsnpztMqog2+ToAYKp5WyV+I/8cTzbTRUeoRnWBSufXPCEGE
T8YigAUNnrUP0w5cvF5pjCnZQgA88jVIUEQjji0qEhz48fnWHB8Qwado7kiT1W6Gn4Ez1e0aqpnK
g6pxwJP0BhuglRwbau8SsDIC2/6pzeZVjLwpnVYbGM3fYNxfpfz1oDZ76ewoJylJeRE35bepl0Fc
oR+mqR5hggsezW+D71px/MeXqMUwTqVI18ijx+25y9JpFVi1rtpMopZJmOhoY5MkVXJdxcZ2IXeb
PejHB12+YFLy30KQV+uaPRCAEi0Q7VrtaqjNfJmiDecNt+TfIEcQx1TXNzkZ1buFm4zde+XVWIeb
9ZRK4ln2ziV9x+2a8gD25KbKMCQDkQ/gIgwyuCZeyH7VEP8L+s4EFyWRnEhKouyId3iArv8Rt+x8
KKQdz8LUc3H4q3+xS/jhzB9sDY79qrPIOhgV6KE7qYWldusPFGJmG0XsIX8gWBdDyDmhDMIM+UdX
1im4V9+h63Buf55COddTQDl6CfvasvGtYPsUPT4G3VgHqCuus+eY3VkpFVQK9jFwhV0NEOz+jXJz
jf1yzrMI9aZep4NWFVrYKZGypfpX5Bfg1pE7Ar+s9crn7M9i15q4SjXaAk34M0JjZPpt25jhWgYD
Tf2Ya1LeKn47CgvJkSnx+hEg7El/9ZkAHOZ/x6pAFA/bZZHZH5sYfZwgVWSOX9BoCz/EGS0RFadi
lkdggAGpvAhh9mD51ocWdfcCKg+1vC6V1ZDKqFxyrwVo52sVbY4R0+qj3iht4ne/lmx5Km3eefNW
PJf8SI+9VLYGHlKAYMS0NLDWKCXsoaHL7wWZ5pbiTaPh2EL9hTSiP8zChIl/VyxQmtVSVl50gs9a
ZUKSchgocVn3hx+VlN9qw1PbfJ+XqGW48kEQTEzDqdROgee7KED0HmCE0Z65xieBWdjQvDey5nmi
cgv6DITUD+WsxxV/z3IZUcncB/2DQygukvg7xuaf/XrTNrxARnb8bN2osjT6a24E9kWNDI178k5Y
oIG+Tpx2cMPm4oASAg/Fj8N+60l760u3qhaGjPW0l53jZhlcIAMgrM/Op/LQ/5FHippN4n3kaf9I
R9+uP3ZiR7t2fo0az6EgPWnm7AkuUG6BRCD6O4Nm+AufHfkPCJoQnJwj+XgyILmEOK6lhTF+/xnt
uyh1Y1wcfSBFm/ztOYgrO9Zu2T0QfeLX5iyO3/um7L8L3sJi4PXmuh2o/0sIJq+4HqH03rpFXy7N
wg1UEC04139QDmDZP2qkouh1alL43VE+buI8553GCfrM5rNRdRA6ZJhwU8dk2sJLObmSgdaL1ate
sV2gbc5I6N6P8rNd7WsPmo2gm3JuELK41GsZkobJsUUxVJ3hYKh4B51UJ0q8l5MGEoaFuyZ+mKZa
I4codHfNSznApYJF6a1JHCwkpddNytxFqR094GsAJjJIVrqWQGN685g5ptXjxDSuUfJ+8lUwKmbY
vWIQ2c4Hv0oUdY3ITIgXLC4cIsyIzPmzZFnU4GcW+dn2UhVRFRw1UWT6rWZC0fhrXxYfw7G+lwCo
/y9kpZ1Y5fjJ9fiycS2UYPqmBk/tBhLd51hnS08R04nfhNTLuw2VVbx8VN3eSHCCO1fdhIDwzeJx
GE/WzDUG5dnGaO7iSuTHqRcBpzVzcu/F3ucPILMIlOcme04OmHoTMwPVibuPHUffqG7difNEZR2K
2AGyrPs8uRpjJHoqAEjVBriHvpyk75HGr1w0pG3mmg5bWJp+7F433lbZoOx0145YE/CgSqKcHpsU
LF9MLDPRViLJJXFzlnM0xGIZZP0FwHApfm7odqN6Db33Ws7rLGDGNSMDvxVEZMZjtEQpwZ91vDSm
FoncBzDImG9EM/Gi6/eYewZTJYqMcG3cm4P9RPbYuKfiHTF471i2C5MDsHHl7g91fIUcu2ez04jh
jgPL8w+pMGez6+p0ZD/L/I6YtbUAd0eOgASIly1U9fJHE8edPmNGlA4FjmZuua3MtF5QUhDGJjSk
zaM2600Ru3hVowcwJhEiQs0XQ40x4NLUx6an8agwRUmVBVQkDUshu28R/vMv5HWz4Cv0R5LgVVr2
6M3tMbpYYKrmcuC7xYdOWtpOLZA8FvWlBe5tE2DkArBDaizo41K4cOSWPJRwfTEGLBxtTXFKaJrg
2MZjxlftB+zmKQ53/NAITr93mAMmZ0l4BYmN6e7JCCkpvEu+eYQi4g4T4Y1RwrY06NUeK5q8Ky6Z
RjVqZqRVQkAwh/3hQlAybJz4Z/hdU+CFRdDpEi3MIKlI/+/2wKS8XIYJ07jVVlBpGjfCF3qZm2Dk
n2jBykZv9/CA2mKR+3C2giNcOfI3nQm60qdcpsg7FG4UNOPDgI42wFiiV40dEU0zCtHKL2HI+hBK
X/yDAalwYweDM8QfpR8BFEMM9l+3xILVDchlkHm2Rf16hHHDDGasuxhytGGERgFUWGiXSnTcdFe0
+cinL9qRNNO5c9DsQ4NRAenZhn9EOlso3KjkqbQggSlkcuKZ07AOh34WynzfFDkVoC7pjYPYhYdB
RfyUGvTPKRV7h6tVJkwDI5QQwyTcdac+q13zrPp+15O+ikkiePepIMfEi11VywZY9U1fr6pihkaq
p0lDPUcs+DnBwKvlNrgZFl4bMmWSNg/C6aCLZo78hyS/NCqK0bfyHoix/pD15m8CboZte+5aqyg0
B773yWSLIb/mNe+AP+DMO2rLIqOsNHJeJmSCDxkyO0rJdNXJ8CXlj/Qi82su9iTu6qEsnoBVKqbL
xzyuP0bu45CRtQKnLU5OuGUJ/hp00K0oqXx7ta2NzsqxFIzW3AI99trO0mxSbeb0/C5SzyJ7R3Ui
mZg3uKiWEAkBl/9Ockc6KTb30HS9HpqXdvlnAEkgAuRYl2y3oNnfUkb0I4o44Gu2/KcKG5vAmVZH
meYwOvXVbWl+9FH30rStLvrdrFt0H1fgGnwO3cCgthBQAco69J0s303ENXX2KVN8nz62TG+PyXEy
WdASEcnMaI98gmQHLCeScPNpOU0CFrEzczb9XDYvibgwjw4fiV1+pWwUcPeqUtprLZu0sIenfiOB
iyg+gPg4GvPDKWi6tLFvTBXMfK5H7V5icLQhW1F+zzack8fIHJhoJMl9VpyKTqtucrB+TZMrWBgw
a8Id632Hgc7UaTnTjzBANg7ps1kbH5qv/6GO0Z4MzYktRWaT27enqyUNu8Pb2WnugpMMuuHVJRNp
xg/Kni7hVa3cVnJgoQXByTatc59WSYlbyIzy3vvBrrijyzkyrL1q5T5Z7UaYJWMmf0gd6M5Ta3Jq
rvw3GpzaLnkQ9fDJtiewkGtb46vDLfZmK1F69mhZjKbaMNo1aYtzhUDb0aLLcNCz6PfCG9JBMoDE
wZFMwEfld7CCDOCY0UO9FCFMPSgb4KwD+aSFfIUnggy/mzoiH1TAT7sGiRNA1UYFKduO92JUDjH/
ETt5jwzbsqZdksZdiJ/cDYYSWS9GkBMW4B8RIaUMaC/7BS05fd12IH9vJfmwZnGDGLzDOBd+40Gf
R/vy4/zrd31WGeRPzm66ju/VX/XuKjh1TEIdyCDGbQ+j5rC3CbElBi0p1mVN6YhGqNaPxLej1w/9
gpW26tEicloLpBYXckMmnFx7PoDFMblhAfk1NGGEK5kZWN6uQhLn9BRXPzuvU6upCAQvqgWgIuUy
Of1kb6tbDL24IjTmfKqv1rnvKzNwAgB5A8OgqtZzD0EenRhOahIZYv4RL8r57HsT5LTdz/LnvLGp
REKlqmpYHcZkknBLJFhB0sW3whHEsosKLmJtywiq83M1xawLb9o0x5C8cPrAj0WjyE+v6PWpwc5V
8daiIHaE51J1wvGGe3fNX+Aduoqz6gtJ+vXE/K8VJln+0wmmnzMDMXzMVjW1xT3LqID4dRSKc/E2
dWftWrCmjKz8S3iNUgy49fWPAcVCZ7PpfFuY7z1PQTbZgAibUMdP/Bz+hiTCVRGLQRO+AlPTZ1XM
36EamfZxI9z0OL5CjriAjM1/7ND+iEtJJub63iuft24dpms0vwfe7g9m0B9kzOJPMqJBGJzHYxFW
sN8NIWQBj1LWOsrfrH+ZRbttEITTIdfSJEeL/ZkUefrksZk193vXQunphP+Znp//Y/ldmkgbHhuF
2Qmxv19FlfgmZio0rEY9rupH7afdTVIzIKHV4+Rx/JLIgUlXFAlVwFRP+WbqBZfb1+dkNo5QLygV
gW510+vl23BZA7nSy/wjf9V3C1KFarRp9JWbdDgiLDOc8rG54gS11CLx6GFVSrYSsnZdFm6kceVh
A4zOfVnNcJDULNQU0uuSstMbK/rciMK0EYt7EAE9v3K6Cpv5+aSPBMIuTTvRcUJUD82sOwkNvKoo
jZj9KU5aiK4nS/LTld590qELsofFNEFv7XDjI0u3gyNovCETzfuWo6Gg6Rh++fQ7RDC1zAK8ZXf5
9yG1Vy/RS7g2YH/6654DBQIKRrENcpoCMl3Y5Pctk7O7ASJmkc2t0PrTOlAmLkdwWDBgttAJU6EI
r/tmRFKm07ttyc2tWDuPKZyTggLP/NC8wXiC6q/Q64ru+dorVPSslS/+VqE4SRGHo0bFSDZU+F6c
dd+d9xQoVJfSnR3y//dQbngFOwRMsYUKrETw1delgYwJn5QB/pEbUGM1Jd5w3C5x8RsDt49SHucZ
zZ55jdruvMmoPLbfleyJrjlusDsK0ZD5awtDFj1EGcxrOhMTm6HfT6SO7/RhL+xRXDfD7akGooZ+
0YZzkDadheCafztVKYikeOuUlOT9IzcyKYYneO+our46MmFkcf+dXG6MY+oHZ7+87fJRqXU5UExW
LGdm3d4vk2cxY6yvk8LQNCT4HFzFv20/Ekw/t7Ar1IQV7D43XO1+g+n2Gb5rIUlvNpiz8OdHrpJc
VTxAaPvklIEFbgnCUwdv9R2VVzLyASj9x//DLdQWLGqPQolPs00HtZNXHhviJqjLPlX51JOnKtym
aZwWXcVNc4VLZrZIQFW02Nbmy65PqUsoDal1qaQ8BhJJuyLK4UH4832ZPXYj2B5uUMlg5tNV1N3P
4Au6N2pbqqoxR/nL15OytJAhvGvmrtxOcCfH3+5gVspwVajkOs6SFprsvZ9gBOuQwX5DAk7bxRJP
Yzu1l8k0A+3QUojDeN4kNRry6ph37laQCBJJXRqQrwz7zaNHuLcbh1vcy56wGxNsO7hSp7jIip+8
6jmVlPt/IK75nMT3ifhV7whXwy0J8YDKKfqFGCtxl4uopxB8fvCjOwk+a/ddLehuY7KMju/2jfWq
L0bXUXU62tgVZLBeyC9g/WZKCMVX+0EYs48HKwuSGNey0sXeh3+a6aO589hEs8/ewPb7fw6NqK3E
BqE9as8kvQQyi3tfQgXC34HPNsGxhH0XrdegnkgTBLKXhEIjjiQW6PXvusUX9JbJ4KJtzEcbqUgk
3mRFakA2ZQf4ZC3cn3BC2eoS6vhNS/2hE3qaMBsrusbpmFDrvKPpjRDxBOQOaKzdGzlCp+nWoJKc
y6c0zAuNUEPP8GFGN7IICyFT43BQdtkgLVlL59TfdoxCtw4jpX8glxnFLWHMa9A3/PIr2TZ0YH+a
9kcQ3jGlwarjZ8jvMNUjNelyt++hwXLyibleesF25xhqVo3FQ1g4NDiD/N1rXsBam4jsUxTLgwvQ
0agIJquqWNcKkYgT2CGLKwEsSn/a21f1qq0dPAufhKRhmirp4F1qDevTYgUMPidz9sxWQ9cY+LM9
MI41WG6ExK1t2KopnHMNcxrp/SCPWYn65vnm3aCIn15SsHfLaDa3WEgKJ2HEJ6abIQ+Ez8scVFik
o7lIt0Feo9PfOUUn5+qPyAUeOzxgxGqtHyH1tcrSodRR5ckgYtSn3QHxfhGoSs4zsOPC+35QSpVP
AMofB/Yd2S1mb1xNp/hwvnT5Ktmk3Lsqcdz3HJKWC8xFpbfxrv0ldQIJcM+l0HWFRE5t9o1ucqDH
GO3r+WtD8SarLN9lvT4T5DUbkqaNoJ8g7bqMHBGuXvO4h+cxcMK7b0ve122pXd+QtfSP9cU7GTPJ
l/jdau/ej0brT1wbuKOWgjnfl52GqKhOIJcm1ybrD8DUjnhtdbQP3n8hCtmQdYhIJA5sPFMmkoHJ
NMS0I1IhPEO/CFEFmMuShPPbczpyVMh5rMTUomrWTNL1kYF4rwRCJepkFD+wCO46krcK1bWsRm0S
dbB1hAp87btZT3bspR+hCf46keDXj90WQ/AkYAoIwOL5Ph8AJIrn9ysKwRJArRdSyrRzB6zloXVP
irS87czCT+pUyoSWR79VkgnoA91/yRiJJQLj5pZXQwETafL2b0tqOB+gMokqGS6sRSBsrudyXWzJ
6uMr7H5Xavcaw2SF9qdgt0GTC+BEA0VhEftAGjQPoSkTd+fnvLyoAPxdc3BtlbLlL5LqjGXjihlr
wkKbSKxHz5HZxi25k1rweSgeRYyOIkEf8KePDnhrVKCX5RMUZbFVyeaP9KRyvudTSpP0NNT7Pe19
POAsuK/7fbwM0D1TMgMMDrHDpT1GgxZCXi0HcXYFVE8K1xxYRIRjWpzwuKDkRAN2eSZFQLZG4OZz
ce4Bg4Qy4B7J175ZFhSJrkIXIcQGO1eqtjHPoOolmoGxZBm8zsvrrZ2b20lOySMsclbQsie3aihJ
sKTYEpkHzndbiuoOvwjB9ckU+pjmme4NU//EmdqeNQprVZe9UrJRwwOS5Y69IwEv+o+3amQ7eate
l3jmIDSpJIN2wVspj77TJAnVu1Q4YMFw8Ix/hYI7oZj2UYTmnerbTth+4Putq4ASSHytRme+ctO0
eY66Q9AgQOzDLcA16PBxhQVDDq+r1PmHVgoKMktaKe6Db+RPXTd9RE4eRDeYCimmzPZjQiD25KpA
lu+qUKIzvD+QJbJdeDzZqumubCos1aOVBSl2jMFB2dGLjR0CSCuNnLF0HFaGdEOmVUDNHQWRWNuX
+sacKx8/5uQsBMxqVYopG/OoSy1GZAIHw61zD0oN12+O1rbFxH4LAclF/hMqJiTiFDNcIuhyg7H1
6la1QUyEVXBhK0/GowB0vWxs16qYQ2vJBeHma0zMXuGG91kg8wstoLWqlXVAtjjIy9jFZgdwtVD7
SHSKCLJZt8BtIzrqWGMoUBJalG9CNsOH7x4cE8WoE8Zgh493qL79Ycg8MDNb2+IAoveyyfeKA13B
Iq6VqOGaJrspdNPXj+7R30b7idA02LFJMRB8Gcw4un/M9ysNbhnDcYATFgAvfeoWaQ5rV3NSyKVE
1a9OavIO5Y0faiupE3jv2r/DvZJ3wOs0J0K3yj9PkPkajtIpmXlsv/qxPKQiDPUXXtJDWmIJkcys
DTUEdGcFYHfNNj3XRTxun3i2Fxy3TGGlkgLu12u5F4254vlLTEbSKhrDm+ftaThVenGNeWx6r9vk
oMPMVcM6doF80r/OGvsFbSFJ1oNff3fE/c2NqwOCW0r0e6MZ5NxQOoMOAApEpvrlTalcNDv6tFLr
9GcyVk/BkKWgVqdNcwogDUn06gf9U/pOyORIMTfYhgfzzXAyDa4N+l4TgxsuQTxGAPufrLI9gf3T
bk0NGijRBXs1V4BulMEVEXineScP5iVZaCriwGPQXvUKmMntk3OpICzK0bSwfJKz1cMuznuZBX4v
e2O5wxtdaVgsJ7u67k/N4w1MUEl1Cc5yC1QZbgJkmEwWVXPS7DibZX34iYhDwXM4/MyAxNwk0pft
ZX/NGjon8t4iniWsrhJU5a5CR1J3/1rvEP2aq6POToeDvsCIkIbtMG3kW5f0wOg+uuiEGg1ULPv8
c5ElOEfQ2rws6dG+rJx1iTNDtK/mYUUZ92GeGsVzvYxSrNTQYejAJ+gCLZ3JJ1zcAZ6EsXy1ooI3
4VNEfhAneXwIvd21wjumQhhuawKiCZRJElbMznM72YrwO6UrVrqJXGA/gNh1ySBFFt7W79MBcsA+
ssZZ3V0hDg2DdstJwL9FYP6g/jU6suTHyfFLWYCkKr88QXEPF9h/mryNx7WIsMjq/8FaIGFcuDwX
vK/BlvCHv40xrneXP7satWzlCj9AeSsrsrz6KtPisqR7DCkxVOn/AazVV0HJCM4Rup/DV0kKVZUp
/Eexv/gUhWukeB4OO9W+fMrMr6YdIVRgIsibp6QNK+NzH130bnsbzQjoZcHXHsg/PBQyXk40oUDT
0k+SY3486XjsZWFh7CZXc3TQh1S1Dj53UZTBJIqS4Kmr3+pK6TNXFhhpDudwCfZWMDcW6qceRM/i
p6jAwf31bNlWTcqMOtkinsmlU/6WtrLrVLtrT3atNyuZi+3U3DT+tAJhx2PIicSnBVn6PEENHHK8
uV+OG1DvjZMWi7UGOmNlVp5nvo+4FRGR8iMNh7bbMbT0RO+Z15lupz0+paoPFnfonStE8W19T6hV
qNlVnENRXNJOGtFh32qRBlcQ8K4QVBrFNVXWk7AwVgAOO3LUYdpElwzI5SD+6Drk9bYQwWLs11Z4
kpg2JWK0Q7m1H/MzOmoo7Z1fVo7JNjuI0kdL0LTUsZ0m4Xphw+SkeSYzEluN9dWZxRsbIzBifYhP
+2fxBpf74/pAvc7nEjIGIH3BczJA6rPKI7T+3vbeG9aImevPjQPiDs9NSWT1AcdVjeDFdZ//NlHV
D5O+72JcJDWA9Jx1Q5pLJP4iEYR+bYF5vKklZSiIC+e1nX2FsbupHUvP2cVyjE9QQAiDle103E/1
vmZqL8e7MJtPaUO4khCQUmqteotm7rmY1Ec4H54dnD31nUrzPYYOclvL/bykN6VXjXW19ji24v/d
vdMAgCynWeyrayg2R+tFHGx22THz6auNSkxqrPz61miR58QRcZE5hpToRvMEuoXGRP29Zv54qds4
yBedTyaR/lZxvpw6dnl/0viKtAmPZCqYr6BdERPXI9S0Es7/L8iAJBb4W+xnc0XNvD7VMLomr69x
sXN8mLinMc0p9lmVCfqnBzp9kml1M4ChBURithiFdK6I13paHAQINbGrFqLhtn8T7eNH2w6LP2ME
bhJ/60YXpOLWFIsFj8VY+bEvWvObBYg+itgAHt36DWk104578bujXACjRuVS2/jVrfU2m7oKicZu
K9j2CCd7Jp/zYGCZy1/ieZXmNFCDI0IF981uDsGRCFLBzIxdss1IpwxSJjNS+ezh6Tx/f/8np12k
v6Ra0XHP0ha+4P4ezFsb7oV9ABexvlcVjXdajH5waBvVtmP3/BavlVbTv9KGD0IEPyrYLO9mX6t+
f3CnEyw9RqQIDPPriQ/y0zffLXN5TUwod9HYIv2M5CCHRzwiVSd3NhEU6e0/bs6sEPF1CbSx9uSi
lpCfXyL24lmGgeH5lyT+hN9+acWES5EKubypSbdBT8Ju84V3vr0lai1iixV/xXxVyc2JKIX3eawg
YBOoyStf3/LrYGhVlwTD964w7vNSMXYWpi3XOiMkskfmfdbWu915mYbqWtMdiECddd7ZTsmCOdIW
fb7dkCzlqDvN0R2IJ4KAyq+PgqUp4BFsaZtCAMb/vvMovPkl7EdHD1qC3xuWiIAUn1yVjmD0AFOu
rw+H8zPoU43cg52h9Nk80eiw+G1GCP8xSvUXG9K+YRDUyj8hoJhH6pPASgiihcBEoYgA4D3c5kjA
nOSKWbsr2rv5RBTQp2DptwPS/wbb7gUiT9TGNzasRCW30jHTmPU4b7/vyUobttDcpxrJWUBhnbVO
fMgAQFu+IagmQTeeTkmNNf+sM/zlrohLPtFBCm02K1HB1CMGHQTdtXNT6J8gpeE+7pBameMsUDSe
R8muNxAy9unm13ufomYOLG2zgkwwOuavTc8u5fgYCyWu6jMdKOFOuyMkkPEgDPwCSejSQyNLCn30
SrmGobDlH8G47g+nX4O5BRJS2tD/g6E5PAuW5/w9B3nhvrqRvXXyKJkeFZa8W+GvUA9RzwpPJDMD
/c3V5gCtp2PlhABKVeQ46H5IxB6W9kByozHvGuq0ysz9MPc++OvJyskRtJo+cSM8FoEewA0XpbQd
SvcIaY02WmDFVw2Sw6ON0Ji6epTvU+ExjVpNI8JDZvfoaXP+fSq4IC4TzwoNZZolHPekrnZtpZOI
xw1VdBW6aWNl4u5p6bqTxjMMw9bKOMZVKZ7GqAKu+TK5Xt9RW1tSlYPsx94bTpy1vqL+UKMvCgo2
w5GIc99rVS/tQMKgSZwvFgqJG+yGyfDhMfhxJbe7uRAmGhttVbqyEzT0TwST7w3D2acMCptkd0NX
IaVnAzQQLekENM2mJC7rLaxKgbjCU+tn5i8m1QEuYoFe2eYOkiEwiPb+8GQlpN+xORfAFSjBefOJ
qRRxKMTdTR3uxVdXEai5MS8/EMKjSYMA9GTrVusP6vIJKJhIVE9K+C6pkpnSTKZdEAWIlxybLQUP
5DAR2zex3HEk+xvkWoNMT9qlofmJaTXuJmbSyzCxB6S/r52yl9njtem4/pGMoAFnSLpXGiGMcAhR
5Rgnair1xwp9tvxS8rVOX1vtOl2XAjiOm0ftPjaBnN2+4E6bQS/F+mwCIDTSqU87iELJoRj1xF+8
n8or9PavpxBy1AbLxxeR8325fnExbNLgXaU3cXHarVNEr8cmfYqaBfgnol6f8VwV5y5ysTsQdGMt
SupIxMIj+2YMjD6NtEPNHdkUpdlSN77RLkibaOSzMhbsyHqTlLIfN/Hj8PCKOI1/BITYECDGKuc3
mHapOo9YAgrlvMTMWUPZP7xA0z51pIYiU21FrcjwAApa/IHZXG+BU1AU+Fglml1oSzU6n2PT4VPx
FEQY9c44ECx8jcgN22om77VQEzcoaaO6ZC2tMRPbFftEIGoRala62Zf9Z8fvedgrq+WStoBpX3I1
GovDddHdpl8axfduFkZRoKSrqrBuzfR66AF3VuF/gNqY8Kre5+cp7Dv1X8HCagoMadyQKwhVtClm
P5CEf/6k1WhrLQQbrPn7zrFN/CHFX1CvxeY5k7tTlITd/EWXQZQP9HVX2hraovejwya33xk5nZ+v
1J7l2GldpFd+eccEV7P/lFO9U+8DpIAtsGOqzwHIK9g6dYuk2tWh1Can9M5I1QOeBrEGAwzw9rSw
OKU57/GJYf331Phn2fxBXQqyqngeKHnvYM3oVb2H6/8aVst5hLrxq4WAliQ+d1j5Ng0T7JWECt5+
eti24uYbuM0YfSIIvV5hxzsh4JRlMQAvy6Y/hOFL36TxkUsXlZNRWiqohc11ooRTWz6Q2RAAX3e/
oikwumdoDujodRMsNoGH65WX3TtCBQGIAVenUqDkH1tOYmbwhqgJkxzzFSdjb7UDJW4HJl8iYyIH
5kD2WKsQfLmFxDPOHRaNiA8PVlvP7yknmCKzzekzKbrs15APt9oPoSJwa4RCkiMLy1A7reV6rfmm
SYkTxqSugQfRGnDF5eM6M5t4JXiS25m6Z7ByH1Y/yUHK9WlEzDzsPXIoxX0Hd9YOUMPqFJZA4foY
TEoBz+UkT4YCjkI8Y3xtrUwnZi9piZzZX4Pz4/Q58r3qGy/Oke4Va9kcFJx3RDAEdQM2zJP/olag
uUPwtC1PpJarZpprSDBcjjYEd1F5RImr+D9jHpzCZaV6oS/SvdeMGIwcN5aC6zc1RMqOZG6/yk/O
8y0B7gDSlNJTWxhrh61sTbPCTVqkmrThFHga8re+qPOIl3tsrOmEPa6Yp70B7GAJ0OqKTPcRUBbX
2t8oiEXRgr9J8n0QimpcrFEl5oEkGQlgckQRd3dG3WV+BKRJDVuvttPn9rbZsckUsCR7VaIGkLe3
JqWbiizGs9NGViiJ8GRhQA6TqL733/7xiAkqsVqQm4XIh1yjFsZAjMrmjVnItXgFdeZDAMdvbfGq
9dN+HHgNmC83DhjJQ+hZ1V/inT73v2JahaaHvsp710lLX+y2MyV6uUpOM/dzVW8byt53b5LM7+LJ
ivXX9wDUzcIzRQfaWPkfwpjMTwwqpoiwVe2naFyepS581YnNiO4tF8NNU/8OhcYItgbMbzv+bQ6V
yGVbPgt5etn+Nu5gG85witdoxjV7oDlCBF51mk+JBuJYcbXfhBMnIkKqjLKvfX3Bk2pKc7w9tl+z
djqtF1tF9m5uOg9a1gLCLGq7OiZ/ojpih5iwW1TXOQkQNuZrG2SI0/qJY/5xEsM/asK+DMy0uTqt
YSpZI0UK9L9uF29eo9lOtsxjnYSDW+5Vulqb/Jcaw1i2cjI12PQpwxNSphyAnHNX1f8+Vz0CBE0D
9zKpaeYSORNj2Cx1iQawuKKmQJj3a8hsSCk54keTUpmvnleY+b7P1xtzVeKR7zJhfR9mzLXwqJ1n
r1p9HechEFvonpHpeHnr62H4NdXr/Z79LEUtkK8V3FIuse2bp0zYPieI6AP+x/mDJ402+SaeyTAK
E8jD4TXXX47E7TsBZJMrjPTk/RNt0YMX8I9sDheufX0vcjYc3sOQZhNAomYrHdBICLiP+H8c/DWX
SeERSaHzx4uQvYTfarznaf+j4TmXJQGc78yEutxBZXmKsJ+4hzxIBGIqbRImju6ec0KDFLeHmy51
Z8aZCdoK3KumzsPuoYQ+i5VtcaHeXjQ0H6x5qJJLH+Zs7mgh3mv2ULZO9d8e9kXar0wz+yPlt4Qj
DOzVsgJN7O8V5a0johm7PDOvDFXAPuoUipo/EK1rxso6uIL6gTyG/oRBJinbUv5eIxlqQSJwj4jG
GMnMkwJ0NsipuLMQKzqyHumCgGZHrclaCarPhcI6kug3rFsiQCwmQ3c6Dye3rCLuo5PPyuJOBvgP
g5txat/X71/ChavJO86Tcll/gtYQO6/943fmA2o+OvIOEfqE/pZ6Uvdgm2v340EbDAki6dPBzpIm
CNBsDaViFzlt5Cg1YTAaj1TpLdjVyjFVUpbeikLs6hNKgH5ySAl61sJi7XHXHaCer7FYSPcdiIIu
Hqxf+gF5hbQRoPcCQ/gT1QI7F4K5e7eI2SrzW5pxfdlWqY1xMIhdkdTybt3tHi+eiW+8GnSz2pEN
R5rWDXN091E9HxuZgL5TBa6AYUqrA76Q3pg7VwmkJey39HYVByblC61CDzyhYptakGIoT5YWOduK
yBpq43xd/dNLzLJOY+95lNSOjFdvrrY4ydS3+cEVItIizdqwSI3qbOqEM8UNImhmmyNpa/OW+zzx
m2QXwLmEkM/W9s3PSTYru3iEkS3b+/M6763n+p4IhfjjgwdCz7f2SbLtUyL8HxmGf2S2HEZ9+z9q
rsk84XI0RATjhJarq1+DNytvNA7Y/Z+dFHmxD3v3RdhthH33eV/Uhqj0cazZs3s8LC7iN4iEjsqf
+gkU//gfsjW5MfQChhgS2EdFILsr/dyPedmgeJnuDQTWJbE2/3jhCzj2PYe3zss588l6nsw+cvLj
K081sFGj+5crlhjTsD4Z4+alfXrbb/JjXzDfGveTbo7SdCNdeCBpTe7vvgS6kk5hHegLjdMoyrQK
pERiMb42V9rXDusViUljTpnRb5+0f5AjZNgN+HQV2GtgB/IcZKlG2TUFi6sNU+90lmHWf7kl0pVm
aP9Ynrn/3XFg+P46lP0XdVA8q0049J61xhEREQpjaOBL5HjQ1/QL27OVaO9Dt2PXNZGjbsuNXOHj
20CY14UQ8+Cyb7w98dAZX3GXhGqKPplkOf4P+Z1DXmrhEmq6ou+zkXFHvuKbW8bciNmlo+Gss5D0
4wgRc702Bn+uqC/zp1hxkn7QGB1gku3PJ4afSOcQ05Y2icmRsYtltPWF+GnveoEPGDCVl3qkaoP1
mdhs0Y8DiTeDTn/qBPTK/tNg7P4y15ROfDgzFhKX9OMf/1HwoeQyKTMKqXcrUnQIRFsj2nxlmm4s
0b/mJ54GJviolrjIoGhmKI920N1zCnOpeDyhJ7Y1avmDnYQy1F/KhotfUgu3Qd6WIpBDLxTHuAeq
kEdt9ZTBzsZP/LlCbaQz01vNWxgdXXeXSXKkZalr9Mo50oPxquYHlsXqYrt1icdRfHeo6G8ZpnQH
620bbLBmirghTKIbOSADMyh92AOslEnXHZOqZQJDea48PcUxcx4eAzoUMWXDldvOeJdCNMsiTRnM
WTxetw84XoxTw/AbzTQzjh3BRlSQWyDkfgcW6LG2sSnjG3tVKsEDoEI7ngtJwj/wFgJeotAmC77e
f9Gcca0qkMT3RO3A5c89+zfU9uFB/Gw1vEE74AQtigEWgxUVtTnVWGmF8jUsZHnMnMv0eALY6AkV
HSL7B1a17FJee558SVFQb1e7fsdoyQ/XCEMEsHnup15tGr2lTBnKpjyWxEiUg51hPRaa4kiwUVV5
JptY4RagDszEhuxk72GsdwJcucGdimwlG7tTjRq/j/sU4VOsOJsZ4d1Tz4++0lBRVaMDrIivsu1h
fBBYCXQmrOy9OZRE3B6cNf3HhJE5eZxNV6eYPBTRRe012UtZ1z5aMZ1eNDyEkVOh4DIHyjIZSZjz
rfUArvLuheH8C5WMT0+MBKm7eZS3s6gBgv1PDCfyJ1F9S9xSTVsJXzFiGQ1c3gBpLsDIUz8SaAd7
NiSdaMDL7HLyaZDapeudY9C5ZJPnfSXOiWF+LOVtjwnkTm+4aPS8skC4q2mWf7IZK+g4/DP16sgO
BG3++EbEEvFTdhhBEhkXAob//6+LpmJowEVelGyPCJDjATutEE/G/RlrM0PlR919iYc5o5ANSTmU
i6QSD+ZrT2nPtml6f1C9GHy0tCzcwcgxAaQJqBVFpdfzsWFsiPEwTkhGiAkaFJDmQCHVlO6y2a9i
exWfVPKHjwc+c5oXZnazbkHWEcI4rQOvofhMkt/ly3J+ycoy/r5rwIgFQQk5XqVTrowLlQNc5Gtr
+RFKPpeOIKpW0ljGpzKKVhZn+Ql0JiBBWQnsj/8AFH+/+sRkdC2H3fUd0b2jq401BFtn0QB+pVMq
MaLLZY8F0QtKNwy/7M57QfnsSOrpehA0X4ADL1+xNdTSa6gI9VJQicOk5bG6W+vlG2oyu4NCbbV0
Q3MJpayKIVu7t57px9pcprAjcdTmB2GtZeQDgMmp8wGdrnZUOVPE094o7WnNhFiStoB5f8lT+Bfn
BreZx7tY37G1xDYrEio8yUFzhH46eiiz3cLK5kfTMnFAAErW4w9gzGKSaFam1vgwOOvPiuocPwvm
0J+dJ6pmHXuBv/1aeTP90M5GUUIIkBAm6GtnAL8eXy//kRLRYrPuWZIlEheIIrS2YAv/B2PZDU/P
WzC6Mc82S2brDDE91tNk4rEmmx/dfAUUIjB8YbH125Ou+rbnLCsX7jcl4Ewcn+2+AubrWbYiDbR3
ILs8m5Hp1p8qhJf+PvMn5MIBP2ZCH4X8PqZ9nb0Dj+Kp+Y7T4+xFLNzTK6WZu+1lBpamAkK5DVxu
7nagwQCMhTCYRHpdGn52kie0HHN6NlBPwemLDJtThCI1IUNz8knx8/E0OttokQ6Wy7CdZyBqm5QO
GL2BMaQxvasG4uRCS0kgXujYMETITi29qXY9OpJxHyjMqu2Ke+5yknM+gCb03oWS3oNPMY6q3OCT
cQ4dqojyvF7bWesV/vf0ysiyCCuBam47WVhOoL9RpSh/bsDHQwY3ejiGksKFgFC6hawVuMV9XIPd
A56CMiPCbAPWRW6RbFhO5M8gWTHen4MqWYXlQzH/RRPV71CdktKMcRAuwn553Y6RRLTbeC+myd08
5eQxrvMMmfzwf33F8lxRXpR43jGFpnpXZw6ZmZiYw5g7GQ0GEN6y9gdXkQaZV7IyTxSbPE6m1Jrh
gdN+xfxRyQekc8W/4LA82SGTr22M0h+Rs191zJ7Quhb8xIKbLPVzNjKnOmmsjQLrRwinhJPlzN4B
tYkpL1EyguiMdz2kNsI6clRFlgUW4HGgD7BG+xuFKb6d8FXbR2iFLUZ5dpVPJXtGPEj355Wi3+uN
P026AbiqjNXfYJzkTXbG6POuP3craQefBLO1kSH1l2GfihgAwIZ6zYkGHyurtzFYXx2Y5kB3RuU5
yR2eN1L3IdmWoPm1Gy9PAW0jINWpTXRjzfShUt3dyebM9+/3HUsRXVy50FY+quKjmytmwyVH8EmT
6dyCl5Od5lkBTW/93HnukcJe8OwYhsS/K/X2X4p8XQ2cYiQ/BX0C4+bA4xm/BMxMOocKT62q9ewu
O23PYgUSprYlVZi3s2SgPGwi3IVqUp11PMI+zGBP41BytsqQlDYsmCI2pi00pP1q8Tm+M9UHPN+r
JXOY+cjas0oAt//C94IvbwGGMGtVlpf3q8fn/2DWHTChHfuSvf8TjjK5J2EHL2buz18+MDbZK4wy
Bot8+86ZplFhJQAlnUPYZUXWPVwGs+UE6wZv3G5xRtbw0DtxStQGqTAxwhkB06nfYsVFwtawVDMl
GSNC0VhCnznDTuKUlm5t0dPvONesQzSMxilo6xiXKAGeMn8y6+t/tN6HMFXhrj9OqrTZ1zM5aCtJ
6JlXa8p1S4pGLdhB2N6qK5kv3QGfiaqAG2i0QsVMlTrqX1DV34d7Of2K3mjytQmCgtDsJYBb+xkV
l8eVpSoh0gyyxCd9xFllmrmNBZhaxA1oCn/XhdQTuJsYv+UaGrKgA+DDV9ydXV1yxPGRRuVarn+p
gQlFRw+MY0ECTwSOIHjceRlk1DtZgm6QEF0uzQftg7qpWRnZAG2gCZP0f96rta61NMyrb8cdGQIk
XLK/0ijkKN1ufWqwmcANApo2cqquVhfV0IxyNwN/nNSSeEOi6B4SAg5AsaYAqK8zv9R2RtcAW47y
a0yNAypr8+vC1upEep6fx4wy2MM5TjvgoFEJ/XNyq2jhfpZPj+tddLZfyCRO0wz5fvJGnePaCrXb
ltwOuytXat2FNLvNc/x4uf0U/DFWhhv7HwMLPwFQFpeKd7jznYQXFD36FNFaqOhazlrKDfM7wEmd
D2BRO2PBbddS628qY5XBGyspWLAQJ6uFbr1msoLIbRkC0oc8Goh31eJB5N41StDIuXklgGTk0SE4
snuWce7JtDn1C0nTbkasU5gn2ODnjoL0RigoFzXfENIY428KZQUQg91FtBt2JpYmRwQ4/ARSwY+u
Ce2kbe6LC6d4cyR9p2WejzgLXOhkTzD9QRCvLz5wmUgSVtZuNM+YCvHUzzjOwuRCOf6EuUkELCjD
AQKRY3wp9WRfMl9XuLOKQwa28PkbPorVRFTsO+WGzq88BHC91HBTDwwzf12OaHDfN4H6fxMHec4K
dnGbYbZopHIULv2z1S0S6K3jvrnDqOOBtLZkeqCmNSatDX6jueukAjn/cURm3Ej56Ywxtae40+59
onZlEwaW1KWzFGgBUY6n5cQJs7FGOflYEeKa1ypcBYUvTxBxf0NKti94JfwGHhi+QI4QkiGTR1Te
BsRTUJs0Ojuwgpph8m5tkIkmZFjrTMwjNwQxkrC/5VIGZMJfhpM4okzZWxVaN9Ui8pVPJEhD++Q3
VbSxexd0s0aHX4KgAB3itSkzWn0hV5ohyy2s0HiqgXIUzKg5rDUtfSE79rSGfH2ZNlqirW4olR5l
kljZh72Yh1YU17bL0f9Ql8cEMb1kyVYiF/We+vS0A8Vr39cSAx29gNbmdjbZNi/n981TPbRmgdWn
IbxOugWKFM6jFCNF8+5ZZcZkEUjupNJtd/qGFtewjWGJ8yqxO+9QdrG4dpS8lfAsMtV3IakMpe6z
IiOjlogkeYQP6tyziWfXp3jDuDuafVShrPuixtz1uQqggbSRVOHp5SgsiLFpv4aEInQoRy1VIIYs
qummhfVM02SjkHRmxKHSCnxZ7lqr5W7+ErhimMyiST82MnjQL5CPi//ubHeX6H2a1Ec38x4MJiHp
w+Ejcmp+hB/Uu5fYthXX5mDbw+6u8dR/04Y3h7XClJ9f4fC9slQ6+5cbmBLHswvwl3LhBm+7jFzX
4GZ10ucA/EXVyl5xU7679rt9pUo/l1szNeq/LRAMkbIRixWHoVwz/NaQpV9JIn30Vf/Jf6LDKBCC
FjmULMirYQy8XBmh/vXZi/2An3sFGTN8TSYrryv1nYFrFGsswXqlIKTOeiiA6mDbCi3KIfNaieJX
kSh0nPpmR+P6hgHQQBNeg1DeuQClq7CGwhKown5upwt9ZNo694LiDTq3whY8Tw9JJA5hAaVKNfnJ
peovcapENBAtYE42t2U97rrGBowZj8JoUWYdpl9LZqeiZJX3kbTN2zlWcedeAyU2SpMa+otRnodi
u+Ra1suLTjEEQ/V5V1Ab7EG9kpFJbEIII5aHD9OmTH1GRuc5SNJQUxBVCLWBMpFmLUqFPpQLNIhh
T5bF7ovJmNVEW1CJWjJJmnMw6L29bqQvBRWmSNOgp1AMARVWTEWzSVEkqCJ6bEnP610xCpsu9kSo
JDTL64/EuxIzEW3BfHdsv575ie/WiA35bBbSlrmWamJKAtnchwK2yFdGsfqjaZyEaOCj9fysJujk
/FpHLSXlwkEYlqGcMgO9y1SAaK6vr+Q1uaBN1xlWT0S6e6ClqAg1QS7AsrhE4Yvi9Rc3EnZp6HAO
q8YalBF40W1waAqMK6V6sCxQvCGLH+BHM8+hVf7Ul1ptgV3M4TAtF2P8vmMNgENifnd5Wit/VjdM
/XlLLsUyCyQgDlf4ERDhWqelKh0/1HbnoxsM/4ElPc85Uzcu69HnFqFW1NxeKDuJJjLv8ptD2BHJ
naUqkjcRr2wnZxKpJoVDSkPedflcYWD5YGl54vqI87CqufS/r8oa5YxJ0ZNLbwNoGuwhKkGM2OCC
IMqAaf2x+99C3D1gSj++eNO9m7gCUZYDfgNM1YNO0M/cV++ptrZ5zah7R66Jse2gEO6b2Q2K9oIh
kWrx89fuF1h/RkXO72Y/564CrV1+QKTKklhEbPyiM2Wkkom0uhnD7hNqiBoULFMvqOf/u0Vwcq8i
nciEgVkIoNahCnE5ZnR061briaAUQCMwj/3H7WI+rweHWh9rePDKWlXFVWuPXdVZgubsC9934HMK
rsHryWknklN06mixWxQ45QuvBYpSuPctFA1vhFc/ZGgraDuTHS/lGcTsT92Do2AG0WGzc//7F7y1
SLpqWK8FcKlY2LW+IBttUxo+ffN/KvbsByoRQCZArYn0HSGQKYOamz0apI0VD5fCxrrlN+zU4KaV
OFb1/76P9MIVkemmO3XUvwVnEDTR9K+gBDB61HpyUOi/cE8mT/R+qCd9GGikFCkXdUbGrXHceduN
HfYibu5dpbzWMF4KlS1H+Wz5L1h8Qo6IpjVw+ZaY798u+NhYAS8jaUdjAtFYBsOaj/B4qb/TnjmP
qwpnxLxE9ms2yjF0E2/bv74ZrtvVpKmVkjdvmP+I8fs70fPKhrDlV9mK9Ri8qwV4Gvn8Ktjwr2SM
eySpDnS8yRZzWzrfzjgLi37Uy0qZ3hYILPcjxj2IoaOm+XbrqlVZSAOM5ho9Fj7pqRQe524sRM7v
Csaox+hlWwhLqalqJwRbrmYKyO1gOCJpVjOha4FVoS8iOJtWLSTzzBooa1LQ3AJ2p1UeQAX0m2U+
A0YlxPw6njB1CYJ/QJtRZaNWEP3DazRA97P+E7dSq4y/NdAlxIxLK8YJisECAARuvyudt8QMhZtF
a2kAhnTUWLrRCJ2g+q7NbfGdyGSrE+t0Yh2dF+JQ19+u5FSftn/239E2vr/qs4HEpapNxHx8RdSz
8dKazWnAL/hy75Pi6mVPRYiYNCuIY4dsrFzmVRMhfX5l2Mhvk/vfVibuQ9sppHJbPwBVhHsykH3O
DQoqAUT7CfrsgaRxDXxGrY4Z1ymcMdLdS7vcvFaL/x9o54YO7zZY+rrTrDkkHvZ932NP7na6xlS5
G0IwkwaIQO/q3RDAVTkAyKUU/9YQAsy2B7ObJ9BT5XuDPu0sjccmspZTnspvyAsHycR4EVY47I8p
buQKT+GbWN8XY8AbcjKuMgUr84vOhk7peDy+WneTq92pg/5+vcFfgA8ZcPNjdM1LxXKv7QdJIlwm
uXAbT3hFlDgaBoxr4WxGbL3MTtsPY08XNbB6acZzsLV0NviHc6jDfngcHT2scUMf3M7IQj5BDswr
ydGC5dWdd27JTB653xyz/8VfP3lm2+Hn3NB9PJHtIJhbZNf0BI66kGH5Vogrf7SC1z7sHTSGhMPm
DhXFEfoARO3+4l6oN+xqg9EwHaiLaWNQs5yCEQXpIEht5YS97L3z/3Z2Nht6TfnLNzQSzmQUBQHH
GzJZFVP0BCYYtv6rgczi+3/cnnfX4+60OaxFcpywiAw+N/0OCIgpF3gY43777DSTnY6UKOzKW0lG
sG43UPEcqsQ6oKBqsiKBPmUH/bmodraDFtBKfJmpWrrjnxkcdsy5OBsZ+m2D1HbPIxfQQvKbWQZs
8rhyJNQQSofK2g09C2ygzhNrRYp6n1xXYLqSodkBgJ4bVu3Z8DkKbdv8DUEAvUuLc+otCb7OfuTY
OCmMzSiLwVwT2VmrcJehwnvhyvcgpX3y5tOsjtTwE02mnMZ+yln1IOsTS6JSJ+kjH9w4MsIo/W24
8uPoni5xbJjcAvPex1FWivzkdlOiXarsuzem3bJ6AiKB4sIdPK4Vfz+AZ97u3tpKxO7O1gvWwPf6
2cPpkwctIrqYOZdRbF99TCcCtPLD0xTgPPK0fjlQKE+mJ/F6OsGQ7aIp60CvwMaWx0JT9Ijx3tVP
Mk+sUr/aGbsAbZYBr1NsNU3Nsmg/GxcXeA0lAW0AbBCoJbnGywoQg5zhHJ/0Dv7fOD336DWHbxhh
0yhdOFHlH85+N00kh8ak7TuI9QqNCpNazOAs6h3q4WrcnFeAe+Uci0PUbyMHbLxlR1QJbWEdtSGl
yCn0c34H8wMx01Gthl9JBTluz+YGSZa60tJ0jSqxKSwYuPXFocYQpN7visrtOzhV1sf+VOxpksDM
8hA1R/zRMgnLaNZ1Jfct8h5V6Fo38ngEahU8aQuItvvq0pgj6bReoDm6In/WDUJhIEB3uaqJ5OJu
PJb0i8/qs7e5vT55hAjAFw8A6rZoaeKXuQrxwq/BY4NEYIveS0L4g2pitoUCPDyqZ1clj5m7JJX6
hnLJes0YoBabOaUgW9PRYOr+peEFNMbyTT88bLgLcq5Bk+rqM3cDBybUnACgUoR2NXqrYv2keegK
QIM/nhClUgni89wAtPdVwlhWbVNNeXTCOgpT+qXUP14ftopq41OLc1fRCuFpatlSuJl+hcy9twGt
7STIxyF13QBlapG8mExQegu6YCTPoUEiJz1PRLspde4SBaqj4vUYpAoNVIV4fUm+4PEIkht/Lhzj
cpYDOBoBu61DbOd3+SRSctgPzNlXiCieqWib2NxWGXv2gY37gXXm3wfeuL7dQtX1LeDoXGOzdaLh
7ciATMRKfCyqwBHgKEraZRM9Tih8ZeesHxMkQJiSJqCyfwPljO5EAXeWuVbiBOlMNmmG+R428WNE
LQ3kg8RFyViTD+5Fan7u9MIAo98zFKGY5Iv3qNKow/TIkjqCQdtn585liYMFlvVV1Ort0yPMDwAS
2a0EPgMNu00nrwm6jPqZLd0CQMBUyzbrWOOPzV/8M7jolY2jw/U2udnT1Mgm6cauncG5vo9/1G/X
C3WdJBlkGedf3rHSWsfTU7H3MiFDDsG3rk69Io9hZ0qvs0TydjUbK9wpMDH12URTYYxnRNU8PJ7V
u22PzgIfr75JdyMZZDrBOO3UZAGk3cw2veecRq+4dewocRiddDmA8eiv4AneAKuTBspbQfmCmxqx
YZsx09Bfo5/Pkjna2PPH+kvIM5mhyhvFKAsiIHLXsEnUuCM42ShvwL+fqnePZ1Bp1/+cVjzVFb+1
u8HhGwOOYiolH7LZSTfd91gA7g3SpWNHFtBlbZO5iy8s6xSsdEm4AVLr4ov69jWpwReZLzXCvGJ9
mEEbOUMjiFmlNNj0mcu/Mtt/dnuwB2d9OTimUXuCrX4xzMq4AzB6aZMcgsYjvcvxyYP2Hwa4WKVm
ixyYe6hcoklqLStuPqw1FtpWTd4c3QFFdyNjiZA4bxEZEfuMTPG2lPFTnGbUbN31qT+840Wwv9H4
46dsBAjH6kukEghiVzVwb6oVZlh9rkTJ5BkqQnIVa9XnExzF3rJx79UkVgFCzfMjJKLQehiRVmFC
tpEz3Uwo24r3lXJUKGYX1Du4Wg0ZXXbnqm+8gK75NLfe9F9y9OqmV5h5PglvhQAVHAaicHfnsEut
aN8TsTM7ilDOIeCUXWqt/UONUeHKvd3/v/gN0cS+/KNhdHCIf5VT5VU058Ecnh1dXmgtDwdhtKc8
LDPLBHdFtZ4RxJ+aMlxk4AOu5M6+EmZnxJcfUS4aVerSuwuA7Xck8r/FHgtTgP6zYgqBN1N2QYEy
mnhoGgb3sXDmaNaLfr9BthnQtk6LYRolZxNy4AzmIci+Rz996VTiuG6m7sXW+ljokfO9/8Qw+GXB
F20Vu4T/1Tr1qMlEaU0TLC2hwxzv+8y2EJRTGKciUyfuzW9wsYvw6pTUiWjrHo/y8penAa3INp7B
Z26+JStgkASkOQ1BqSp2S9UbZkFwcwcK+n7Jr67CTWsTH22/fqaLE4yaWkxkBjRDg/QzWGP08u9g
zrZ5NW9fhsyZmnEyF2gbGn/N4rQIgBOZci2UGiranSd3s9nJG9W6hqKFv4tELpdsWEJWr19ajfjw
uXRAMtcjEpDSOGsJwb23R4X7QTmcszaF6p6+De7bd0f6JydDdIpmMWFNB7B375+4Tf4Vf5Rbmr+P
F+9Brj0Gu3gh9GOdJ84BVQtvSkkqeXbUezfOHCOa7S/HpSm+eou7r0iSRdFuuhAcqeNihMp3ZELz
rcLl2Q6wtGDRaApb4u7t4qZyQnkW8sLn53yaEAeGtls+AuUlxDCYNbBWwjuUyhTKibX97E7NViMt
0kM2sLz04S/4rZ3EQWTKwAWHpvMMVmwmGmQyzVAuDxENc0rnlz6dwVCfedhS1KfXrVAenPazXZSj
BPrSyfT39zG9z0C8mm1Lj+8CvPSYWIM01qzrTK5aWeCTk1xNPAuVT3Fq30RJun6XKEWqETVpPAA/
gDrlUmdcdFQ/5I8Akwd//tOfY5V46zkFB+fEJ+9Wg8WV5wFmqNbNEdg37FbQTxn0clqhOSDQ2UAK
kcNrFEKRBGMsUA8pK87pFHRLA29dn4zuOXz1Jdjet17tomxcrT92foWA84rP7aUVwgeV4H0/9a+O
xIZZpdGwb5fuXHxd8Da443lmY730EQiZHppqCI2w6VztIZpF8s7xXTGz9gdTXHYoF8Omx863UU19
VMCOeleIl7IH/hCZioq7rc1igoLfv9AJP7WeejUH4kDEI2buMQ5HBpYKLFxss86u5oVQ8i4S6L1J
X1oyBcIhU7/fDFCnDSn6JYEW7Nueud/B559iPtwqLn45fxVbHxYWIgFxj5IDY+c6LaLVB4Tk2+5t
7RFkiutm3dQ0CX8tcmqGXx0b0QGpageUVo0k6F1rUU8KZ/2Tw8fFU1Vt2+dgYuMUU32l/jaQUcR1
oCTdBpkf7Rz0lt0ljLBsiiIiBqTXSgDUQ6Bva6JB3JqsLmpwrYisoPyPviD6nijWp3XQv1LzFFAx
Hu4RIXUXSz4hp5GVHv1RjNCITsqbpM/csOVFUdSnxz+st6huLRtML1iL9MiOU5BXglA500Z3BxF7
cb8PZX9t24JzT+nCOdqtS/jRSoBWgTqUM5JRrW6Hc5nPDopFh8kLnRyYylnqvoPW3GfcW5peFDm0
NR6Im9zvJp7AVOywuukIWBdLMt54I1YUASHkjJlYBu92KR1TYMn6Y6a+3Ijuh12GyNup+0AhCjom
0CD+EI0nWZBHR9KP1110vdBOqGG63Nz2qwHv04n41mylXU/OFUhTzCHN6LXNFLkFRmokcWqLAVML
OTyMQbd7h7lQMqHFU0fvEU0EJWRAJitMiPfvHmjjSw3XCseGy3D5oIT/iTSCipLk5mo4mqv+QWGf
toPTv0e9rLmCNVNp2EjlGEBmrRVlFkrYHohwQoSg+yFqF3QqMQOp7rh1ImmQnGL0pxJOE5kRP7Gc
D9KUFYudSmCksixJvM3UoKItM1llmQ1i9USQFRMN7G7JbQywtnyuDqhISC4XB+/oyhf/kXlyDbAT
bniYmp9OPfTP/Kcz2iS9w9mH9u+7qkoPARO+mge7/fP68W5knwDc5SDsHWL8WeltLe/uYxxmRM+j
nuTnH7x0WhSztDWb2/FRZ99ATp/uGQknhQSOjbFZjxpLAhYb+Nr+JEmYQ3Bqbgstf9pNEtwJMi1S
zNHJuImdH3NKeVWyyT7PtcbmSSRrY8ZavPNSs1ztbwH/Tm60cp11QunNCQc/QlTynWpNIBweX6ln
6Y7Aruf3mI+4GGd62PtsKepA2batwOfwBOxKqjRgNpUnPl5ElyJ/uZjDRdSCle6Gbg6HWZQbXwtn
wSWg2srbtMrKZVZZLhFMhgVkvX8HB3/bUk9yuHlYoFYY8enNirQpNFY8FMr/0VDAgFBWvcu9Opwp
AXx8V/z4k4xvLtLatN9hpPF5vXlX8VULSLQYNLZn3x7pzW5gtYf9tdtEl95Dm5e7OqsCYEGgxJbL
JVg53RjJq70umvRv/7h78FgsKqxA+xzY7JHks0zITymAfGJT1ast2rAE64n0oiql4xRQ97uIbWXB
Rv2O9Rbfwkwr/IFkZSD2oHb46DXqJSJDlfztKqzC6tbhsrHVrjFUaZJYu98gTsTBHUsVUGXqxZeW
aeG9xroAgze73j+oVZxLYrFNn27YCHw09iRP0D1P3WzuuTUbJy0OwFFPyB1yAMxjl4m00JDahYfM
Y2zGyCMEutNXi+EfAqgTJCU5ApbDixhFOwX+Ik/6kS6UmWNEE837xxRfElNo+rzxwDIbgxWqtUjE
Ypod0Qy5A1xElOYqwnv9NrwSxR6yzRSiNVkLOHuVqOTUdcNQr7uRCmUm4KcsG01YgheaHmo8lk8p
Q/IVCGkaJnpYLlXgM6n9owUYUoGU1eWTgQ2eZf8isQspfSQZtGQCRNkUf5L/LBfnUxe3Gx14fkHc
Qm03qj3LHKGInWm7VYXZUa086B/sIpBFuexNy3kF+ji0uUqzvuIXsEKM5E187zyONsJXVpJX0f/H
bN6ZC5YnprHoSGiRulNlsobAiHd49gHa9ChtVhJH1M5DZowDpRbUwdYMyNdhowYDi4iyqoMLtpVa
F44m1pj20UrKf7JCgVcJkKRyl/0tBxmunwOn7x7cm0QREbcyDRKI8mhe5AJs7m2Hhk078pcyqdbx
k1jLWi0cq0RkGYsMWlw8cyyNq92hiVCml1+zaF/qAmHfVX/0spQA5S9G8sa567TvkBxtEAxC0GXu
32qTFVlu8lb+GPi9iJAEYsI7v686iW5MPhLEOWJVNspTlFonBz0TYZlcpcb/3Rvanea7V3SDeoX2
Wr8pMjiuK07COOIPDtOzE2w/IJeRonnOO78tu4gppsZ9BzPWEXsfTU1LkJBpYPGH15Bm2+nSfbGR
qgKiVUaen10WVCe/ZgV6kh7ClANUh2C6l4XrNad++w4VEr4eruos/3xV/zpPAcPQ4pfQ/kYpjfJ7
pmaKKmi+4TKGd0EhCMv9HVfu821coUbJesKH/cGYy9S0YigW0L/WGuJnM+98AD6/MN5VL7zw71KV
lG4lHu1O1WVgxs3JOyp93H3iutjpCsZL/iwy63BMXkdzAYsFMY/N1KYfvYxaMCfW4hCvnufQzmVw
ZQ8kpKdPUQLjvbL0OvhIjM/gr2ksCG2ZDqkP8t4DeJXuVClHbTsxatCWvn5cj0IrqV8U9xFpEoyy
11OAO0M7lOKLkbxtURqKHYa1btozww9BhMfTYCtBS7kZENgD4mPxCTXkKjEr7h1yRzQLS4gyhHI8
PIcKp56EoVYIboQeenNP9PodxskFlMp3z5coFa03Bz0CkE4X6ltSSsPX4OpL6/xTMYcrU4r+na2w
jbOrxBoTSsYgj4lk+C3dnrOAhDmkIeLGVPpi0Zzl0maN88VDFfWSPWGEmz9wLt5mCdt75WwZXVDe
9A4TBLzUXvpmhF7tcxPYtJ2ybiVRSGlJA8sKUom8aqNS4QjpRIO5dpFRDZ8l1tp/g6GZs1bu3hja
5Wn3CnhW34QPbqFgrIK2tDBYZBgHm6hC2kmLxEI7Nry4wClYXMzrW3KzdItDZXTZTwF1vjU2OY8p
nYtJXfeFBjarQrkM3Y4nk+/vais5q5+SzLozdbkfFI6mBWHOK28yviM9x7X8I7+aUBpqKizSs+k9
PXN3N3yyDpCrfoSGWTajvS9coQ2MrYk2EW8EhGPNHMVbrGzYwWJqwecg+i7gZoCCSIjH44U4HHZW
HvmU2AqsRWp6qfIiUmiTnqWH6OJkvytJYdivnZ5p+iQL+qRn1XB80hcpQaC/uQA27Ey9UyzoIKp0
b2vz75Z9oILmbb6mQrQ8f3Dve0dtuK1zNpUjRih4Hv+RVf0lRcPsEemR/WH5i5k5dfmlalmsogZM
z2QAH15ie+6K3f0EypheXRbRdwOnJzUrPiYoYgWgNkiUCeyIhxCebeckYQPcsHcaGqNBM0NOvkOC
u/6fHbrS22ndclH1i63i+UxLcs77IjSm4KgcA7wtFXgxSrJB6I+9AQaEniUWJ0WNMAdgRkJvUzBb
SwyDCJxUJy0ErQ24KPnMzYBF8xGnDLa3Y4ejiLuiUs6mqXXwy7h4XWFN66iJWX14LRCg5FpBgGVr
F4bH7uwmHuYhai4YG0Q/6bXVPRhcgYf0RuaAYNCAsbkZsgaj0wvVvzTN0DO/9oYQwtMD8Y+1tNY/
HZVlhgCxMCIVOIsl4v4TwLazB2rqC6YtkJCxJ1VXmJdcCj/Rmf+FTVkCRKNbaQZ8x26ZVgaUaZyq
NY8nyED/91i+VBAAssdLw5dsNRU3VYyANbiQMMVYiypmaeWozzgUKiw3uuEzltQSyeB5R13Vd/pI
OVMsIduJ5F7xyv2ibSs0f0h+MQov5DQJnY18JSu2V7RAntxl1Ww0J3Zu9VxlBq7ABoYjEdKEuZQ8
/7gjLodaCUn6JFVKqPb13gyffoEIVPqSGaqd6uM71eCsOvsbNF2MmpblumAo9vPrv/pNtr9m6cqi
iUJfXrGuhW/uRYik/rFGYTaB7/Zc1isu+MYNTyV4K8ctjVTYplmc2xDovbecxKy2NOdztFnMijP1
x0YUfSwtFGIU0DPfIKj5FnoX3Pk8uMK44rXOXgkvlJ4m42ecqfJ30dI+OOLdpJLA0Bu1IE2rNf54
/pTqYfNHY+fHSYR+Tu0k9gSKdogU87oxKbqsrcDmLl3Rx65AYjWJ482cCf4tmgPjSi0RUhbyj/lu
X93If4h3OiTM1kOVItgLZwxmaXY2/bO8pnmHdiZxB9g/8f0NQ9hlw8hztDkJsKgX6+8hXySOQf6y
a0NpUncioBXbWBHroTMo2o5LHYAQ5H4uZCtpzn49of4kV0P3vSAZ7RlWa4mBUjySinKqwjb+Gm5g
L+r24DkyefZ8jEpnIkJwx1t5QfHI/F/oUzkMzDNCxMGbO34h6WJMmd3w3qqLmWUPji3RWOWNpJLP
d90UV/mCZDKKmUj+whkQfJIky0wnnv91qnx0JiM5t7cqghwApB9uIKKnA4ke8tY5q/6xZ8B370/H
kMGQNcLzeBjkX8611Td2SXJHD3cQRM19ptATjNekEQ2QD2HLkG/67911mqbDKJ1TAbXSqCfKz0SB
zxLJzjvg1eNcAd6mPQeE28c4wBj5Vog5TbyUBpDXaaZ9CUUD2GBKVQo6nWDBkx7NU/KGnJ0BK9kT
J7nVi3sgIndNreB9rkqZrPOZ9adAESlc61nDm8fwqEK7Rrgai0c+3W6ZDFN+7tvsTRfa2iEDm+fd
h8SYyqfgF+gj2ivLdu2hRxGs/siExQeuAqC9l4vRAULA9nFIB4EuV8AFAl1Bd9rAYFe3awa5GlbZ
QweWZlSLHF2Gd5WDXRLzvuPa49ynj7srajsz73jIet02JsBv88c2WAYRhVaZCOyKCp7AO4OsPrTw
9REuS5oTsipedZhwtL2c7rjgKmGOPyg22wOH9/gvDnYD28o4MXpWOc84z+Z26UxRCJXwWfehzUpk
INqSS1+kGH/dkxU5iw6YxYZnRnrbidebRgJfHMehJ3+1A+80jO8dKlFYXH7U4C6HtrbieU6j8DgI
JsWLXX7qJgZWKZtl3pHR4L49SDjno1ozH7VyVVfPT1WsnUY381cglVwQwlL2F6oC3vpM2F5ucNE6
GtPVPn/hnm6nwnXRaizP6z9UZTnV5Mzy7UMRReURBtzoz7YKLMrRcsW0XuXMi8QtA9EGDeMMp+hT
7e/XzvtzOavA5H9OnS5n2G62i6QWi4PS1bd0WyDZC70gqPT1OtiuL9f6wqhCRRD9uS9mwhxr1agr
9DWkz2eE0+ouhMw0W50DPgecZEjrzMwnQ8fmuSo5pMYxrVUAACdD+H3U3rv2hfd8cPK0KX+lsuMS
8oYZ6rU/rRefI4mCgpqvbDkQo9ioNU8KCozpgXNi9dF2SHLeHulxqIHvqZPurCf6AqdHDWOSBdis
jw+3WwuEgWX6SrJjU6xJXOlOblRvHhUZ7lg5CRHL2DlUZx5GpOMipVEeaNecqxRCvOwWZw+qARpR
pKLM0xqCwCLed5QEwyKBj5LMU/7AEFloLYEb18gSqarSLOCI05S59WjqWsOqzB8PV8lySCV8NHn5
Qs1Sk/6Gvr8l3+bajAnydGZXqaEIrgYC6MJDFy63vJUJZfS0OSYiPk2m97G+lZmw3CtC4OMqYTuw
1v5kaACQXWx+OwgWY2zh9mtRXF4rPG6Hga1zcFYfkknPzSEBEg7h5ZmzOOVajDI4FzcCADzoBT/J
H/5yY1b/UcL6g7VwLwO19kDa9h3V4BqDVTyJKW0h2nbfpJJn2iSa7IUIIC6lrgOw+6tWt0t7RpJX
GWx4R4w0Fa2V2GfQSalqBYvOZeuPjBM+/hLqQUdcEURMM8khpYLq9MHR3vvY6s3M53YtcbY9V/Xi
1HO6shCKALqVLMq9MucGfsRyXyvIXpl3paDqpWQbSPEMwklkZWAAv8aL9H+CjQ08fF/nN91u6wes
EIZiHNcpvLm97o8uWzOk/mewVjgdQEjOnR8eLD0qvnZLJSs3RH4YWSd4qV/kdq/9lMd20ePSWHzb
IrK46avbUpmeoPprA+41UWZuGRHXE9TxXbChEmWsoixIhty36V6T9SreneLMq+bivRaVKlfiZcRP
jhLTtyfihg7lntQsYwklMgSgf9ESSIoh9XDANLJNjnVZwrEnNWBL9/ZHoQjVl40bxf4YfcnFRd9O
/MiaZ8Bb0c6gSV0oL4sCyrHO9T+3SQROZk7DvfobOONUFLsqYsGTrG5cVC0k1dyMM3jTmFI5Hol6
QkHgP/PdnWCgnrlYOi96GXhh1Yf5SEtMElE2FF4U6LEAbHjlZTP0ySKK/zKCR/dDRRJlIAxjT26u
s80BikNgsjxBl20jYsNHJd31DHaF/bRFrkz4tZKGDHd0xYV/EOso6/ZRCEsS9urSEP7NjC5qoQzT
MUigIItHDmMmriksY7VBtkOUL96wwc5c4NQJ1WJAQoeL5o3w6CTp8JFNsxO8W5sU5DAKlCpE5hpB
EmhnnU4GyNgwMVgwUglNLUSiew4lvTcqt8uP6s5KRtpBqAyGidy5z9A/LJZWgOMhtN2lSniwyqbQ
jGXZYjXXTYwK5mPME/3YQ5YmyoDPA8mIgvIPUXWYWIrl0zpntyJORZo66KpHrPocwM7m7It6HDS6
A2Cn7DudBFlZ4iLTR2ap9qfUdelKiJW2640V/xuiyYYW55S1413dSa1svnRgLjBP2g9DXuMSFenB
g+PImkBploxBQdk0PPbOWwHwbnIY0KWGrjedBvJicFirKrIXKpSBnF95mam++7QJcrrHa8kO3imI
zqeZUhRE3jMluBtKQQZRT2bM6FyTIpqonkKj/b+JOMiH86mr+F3MxEKjD4HnlFg7TQtxgMZg34y8
vo1kaI0+Z76P0bdkNcJpNzFHzzP3BtEb1FCSNtQ6IWoZl+G6mgYgyVqdzJll03FtklA9yH1X76pJ
nDTc2ZnYbg8Jl7aU+9GM1ZM5bAX4eUpzj+KEbtQNiGHHz8VtaGPwiCMLCDxQMmI1d6no812hbV2G
nFLCcsw92CXCBb8YMmmLgT2S7wPFIjJmgPT4NGdoLhiwqajXXMCIc29GungGDmyiYJ0ZwMZWua2G
hSf9HfT2oVdbKq1HxrfEs9AEmUskEkNOhvsAIfYeRScmwuJdLRYzRRZHM1DzAVkq/7bSpYWI4j1K
0aEnY3GGvcpmTfxorR8YNaT5iodHocV6Unc+y6YZBXXdMftkepw5hqSB1dxbm3GgYkywsGagHDws
4tjPmXzgSJoNCj1I4E/hnFF2uShzld/hFlTpR/kL/XU7M90BbmrwNTIcIMJ+eVHdQ/sb8RSbjuh0
P+1YtxZFI+Lo2v7eA7yKfvKNzWHuThP09mp8AL/709v4le1aWPnRlHEK0GvRpD40FVtQUDjNsLar
7gDettXYLt4//Kns7bLPQZShtQU2DhnFUfCeqDZPUnrZUicDxm6nTKsX1H6PemylJEhRGxa4ekT4
3XmZpMzbz9ggP7UcZmJxLdrRWihFn5zJiYE4TAQinXwv1QGZc9xSh3WL3B+DPCDvzzkkO/ogwm3h
kF+l4yqXjrZQST0Pmlddeubmg6bLEhQpqpI+UrykKfdyxhMcIW3lJ3aJ4zHs/OxTjbQaBqHkz6NB
64tSUByCm/ZcqiZGPAOKpymb8BkQ5Wsha5LEPZAZG87phHs+2yscyqMo3yu2ZrMml4z+EQNjzVYH
OqsJTNZGhTqzCyLDXgmXZdjjKFm2np00/nGxi6pMnXZ0JbDBHJ/G59DWjSutLuMbs2xJ7YfJf87O
5v5tnBrHSjyYcQDoehOI8HNpHQ7uH6rXpAGt3XVxOe+JOHzCa6DGuvSQPhi1uZGYrBrkS/GGkhm1
abON4YpwILyh3Ymv1BP2r7iHIBYkv8p5BK6ij+GM2Y5WRxLXl7+3yDr+ydd+0mA5VbnGBx2mWahw
JaOVvsWSWd95wG9RL8hxYkcnmBBRPvXlg9DwwFFvysShV63hdoZB4nDv+Y710NOHLqoa1/X0Y0pi
4F82ZvM9RRyWNWpvHAo07S/Bvvc7FHqAojnV4lNBAoaE3V72FSF2g6sN1j+HZ0mQWnXi0Xx1AMOM
R7LiO0JXqKeON+G9GDzRGD56NCaTe1Ujre+4DQALLK1rfTeuE9jo1cgTMi4omilxNzXWuw677uvA
/VOL1fxpRL7q2JrSEPNzzMFPDkBDkkUuCv8x/liIn6OlfFil4w2rzjfWNdh7RbS7H/didFkrzShn
HNDxcdtZ+4Z0mskKH3D2eCcp2lKtHol/IxPzLUXUJ9fitL2nPF+i28mQxql6g59yiOe3IlgYZ8NP
2fbiu2JAhxI+Lp9bu1v4fDTQYw+xLkF1IfX+/e7RU5pIxVLv5G6fUtMMj2yiB0Cd3HCChsO9qmjf
2ugTCJ4HR+f4AwEXcqiGo8xIaJWXLkEJiUV5YmBbBlOCxtgh7Z28h5rBiJ23l+O8zFEohjLu/wQg
S+VXdtXrRUs2ghh/YBjfRPQFsl5WguAAueq3ADEI4qEC2Gd10DmwGCml8Cbktl/fAvuvbtIubAqA
bLwjy7ANfzVZpf3TKfV4ah0JnhFwmBknbbPO6SszwT8fRN2S9vpptjDj70a7PF0w+842BgIhmbr2
nwzRDVGwkkTWtx47uDaMjGxD6SZ+BM/f10DSdqzjLJ8h65snS0emrxSFvnye3MupPoCiAnuLS4UM
XHqPHXb4LVilRkz2HKbwKqVYu0qU8Kzn70lbq9GDR78wys1fty+lZsnU6PEFlNINq7VxMdMjTXlY
NFG4whiO/xTPXj+jDLzKQ4k0/vcub3AaDcz6rlR7t0ZA/yYwsVT6DwworvCbLWsvIapQqTSfFE8B
oJisUWz9DRqQdoU3s9YYEtEDx42mGy4h0FzibJa0RwVqdnD5E6LI0Xeyjcx8XGOifznnchNiUPw5
2dOvJWqB8LCUUv+5j+5pJlS5VJVoDai8xfCBNvw+CrUFXOk2oJwTQbJmI20UCNMH9vGKf7nAhFCa
kDBd3QxgxF5AaNxVxnbZ97AjW8VMhNXhxy13PV0GyMu6nKY1mxhRm5Q5UidfUTP5nMRst6KXAqUs
J05r0A+HZC8q+Luj7K7GFOvmRWDAY0xz+wVFAbyTNRodOAlkNqMYJkC+r/faAYs/rzGp8x3bRos7
5RGxtY1kLB5oYJCs1nuygK45pad3/AdZEzp97bKVeIbLk+wN6b3znwAPaJqnsV2QQSF5+lV8nkNn
l4swoVWHMuR1KbNFnhZVomGh7ZgHBFwgLcTYNZMkIs0FhvOA2CS5TPT+A4TOG7YUkHWHW/4Uo9GW
VgRwt+U9bFGEfBlhtG1cla0ug2c+xDdlVfrCu3LcSJz4rk8Rqfi5Z/ltiO7/1VHEvEcJn81yn0W4
JgQFiTY+Hp2Eu5XemjXlueEZbxXm6vjA9wf8jFXPQBkm4J1sQyKwhDkRScg+kjJzWeQxEf3cMNbp
ZlGB9BuqZir9Q2JnyahMw3ADi+X10hBjHSKhx9uzfYKGAGVZ8XcYp5pFz2t6rh4XUbXs3RFbBYrc
y7y9MC4D/yvKO+JI5jOn4PT3M88AsB2SA3Bqvi2uQ1ECCtUlyxuVgP0Y3ID6EMlI1auoJ77c7Y1B
/2OXWYc1u08A4rKsCfnoqCMdtw1EtASKvB63beaEZ4RFqlQ90bMvU9eYgV8Opc5KCmIm1d2om+4B
EIaCLhP5VPtWEckHg6HQKETQ8V9/0gGQm3RwE6ny9BqXaMHulY7fGqZ/6RujLC28Q0k7SDdRPGcn
+GQ2vyDDqdFGQzZpPm/kg1HfCe31V6pYGgsMlt8Pd7UDhHx6dMjJuB8Xm4Kas4UtZB4t8rvocH3f
7bqrSWrWVni79TQjVvmZinLBGduwSGVld9j8RFa4R4utf/46cXD9xIuQTZdtn9FXgPeIeHNy6bK1
oRc4zC4RDGpWSbLXzqYiUcFB2ynm8D3NJUACHE7oceETYcVbySRTE7zSrwo/K4nC6rJmpzHzkNT4
khN5PH9tJmfaPvEGKPJuGjFd5tXjCxipN+fkIWnizRk/tzcSVlx4p90bkORUuo4UuT+L0mdnXKcj
F2Nwu7tuBIR/cfoZPR7mUPCbuXhIclHprsUvJL/DfMTvtC/JYzy8bH6T9MPfKBqS+RvetgdQdAyG
5tuiPmukX8g8y2qN8uDIk4KavET9ZU8X0rIg/MPVwJdvu71M21l+LBeBHT3p/Jy1HzBZHzO0r9/1
heElj6QYvaPf1ARVKAelJ49B+RvG6uIZtPw96EjzU9RIolaudnQBip6tUV2NvounM532a6mplmDl
dEpF+R3cnXdhFA2m0rS9Pc3AzMpz8ne7pXkc5o1FNWw6Qj+tL5NU9J9bwd1QpI8o7TkjRZ3p3TxQ
AsfiwOjZ9ApYE5DZOA261JXqeosSsro+6wwpz3WOppwe8QKd68rw554xhz9k9z9j+Fi+GuauBga0
43LgGVmpEggR+heZTfIofZ0xIfjHmqdh+LW0egDT/mGWDYlUt5OPfSDixhcN2uJLOFOqxA9tsbuK
6jAVBa/FMcUn8K232+nlBk/Zc6EQ8p+7pKSF06OjI9afB4ZK8oXLxdzJbIyqG2UTB087+D4N6hRt
HA/U21aecr2hVnIz1CN27LttprAw172PTuD98X2WgeKuqCbYnYuHDZqeqbC8hkibXICO6ipgSZjK
ey/PlilqLxRejrxdvBS+NhgwdEMdeOnUmv+tf51DmjIxof/XFsGsmH7x0DwX44E5Mguvfd0StGwp
MwlSaRuakZ1XU0+V7JsFJvnXBwBmY1uv6/FW2FpGr3EKTlJoG4ksPGbi5msujANvFVKJRDI8F1dB
HDK2mlrcqcgKc5UFR3OPkXsr7ET/vIlWiWsg9ykkvrEXLYFxw1yQDoz/3V66MKHFBQoItI5I3bvC
eJ/Pjrc4ZMhUapt789oUSDt/nyA88LqnJ+fX9nZW+xTgYYQGl4CNd6vJk95jpR7KJ97Esc/cfTqc
BhPCgE/sdFSfczuwReqoLjP6Gcz8GnoKjfknFd9RXQYJW7EcV+xXRGhVPV5TcirZavpktoKgQ4Gh
zlRAQigVjTUy1SeONt5eWPiFzKUjaNKXOa/f4EnXx6r+Y/Heq4w7fCY5PsdlZ1zfxBxXhH1qS+6Q
6mCHuaoza2qRXEdRnQIbhUu9/t6hz2aFcVGDRPttgMUSeWEGl45PmkDdvnZJov/+t23ENgISfWwN
52xNhcXaIwmFp7YnkLvendg8kLw/BeeiZheKPjNyr+WlXyPgjeEVrRg0XzFX9d04A/rtr9Dv0gRM
NAbwUh+2BODpsVqkQe4FZzyjA4g5yFY2Tt5pnAzBV5OzHIYsLfMgDyMoBelzzNm3pEC3puTZOBiW
Uufl4tcsl8RobP8uUgTwSjDHBwYr5qP4nA7HIITyB/Lr8XHoH4gfGiRs85p05b/uUhfJmfzv1DSm
0qqOXzyVs2DpRpGHqVqe6+AgJwFKbKRKDycFn2iGYgETw5JXHPT9y0G+ttdvA1dFrWpq/QdO+Y87
z74U1wANibhmH+sm6OtPk2STGPy7s/rOjKO2PtyeJ2+QH2suXh8cj7mSai5zbB/KjSfkYdS2LRLE
i7S7Q2kH94xvrIo0dTdrjUj3ek3w9sxy4L/aMHoEysLLvplogDgHlT9CgkunAxlxcHXvnOunAHmL
bgCs7D8rqSFuSFI9t9rYWMw/tMHpIJ4sPgZv2F7BsvRzLuk48UoY0kbqu3AqaueYqMSU51eW+xH9
qbTr5ScAEV8hLhVciC9WfO5cddEWmLfOGpRZXYtE11CzuVNfLQzCuO+/9ni/DKAvAon1/TZ6OEjf
GFIA61zIWJZHxHeU5zwDumxu4l/XrSuHpvX6njaC/ZMHdKwmFYXB2pjJdZJcyDccrG0ez3oM/wbg
OmZE+xev7l0yRG1epKzY6afgWlmlIXkrDAPiXHRw5YRbi+NmkeIGW1nVMT9vlOxT4TNNtibzlHN8
4V4f8jqrkjbKwX+lWsAwaSXJGfWqa/JX/BTxaxqo3Rbux9kR0+89D6UvYNi8vjzEopCo8MuHZ613
7gsv4Bqf2I8ToN0/Wm6S7YQKuUtJQ5X+M8Cr2oFY3KgTv8/dTu5hiQqxzosAo37s+QZw16CFjR5i
EG15n5VKxY8+aZ8qJAlrwBGd+d70U+p0K5i8ZS3MpdRpaya/zMTskS3YkNRIGjxH9bBjV9B4VOvd
518ybcCBNoJASTkCF8E74lQKgnMigptvDFfP28rZIzrBo36sgefMh3nXkUW9MNpgb6uV9y04zegN
VgSZ+wj2yGrmH7iTT4vD8K3uXZ5ViWRlpq73i58Q1+Uh99WlOCe7Qom6evIjfYMEJzIpHlMcbQ4n
Ldh7xrKkZH7CFpAmOJMk9ge+RpdaD/0x3YL8Hoo4epFqdU9NNAcLKwCQkVTSfm4NkRp3XXEuNQE+
NV9a4GYEcHpofn3l+ntuwBQ3cb+r6KsNbVWCCrtOpM+2G/5e61biW45wqBOaqxVqeey6OlPYMJQY
BnfOJtgNHQPRfYMKKsveEIoJog5yg5S4A/RG6rk7hRd+j/p4oXCzkGnsPjwwbqYgPPyrmc82aBsy
4SJT7Moo8aox1/9EDTXzIANLD9FFhmgEjvaJBzTch4iS2Hf1al1gR7DLzOjZvznvn5X0sIFTSxcU
gsScQU4jakF/rfSXbH1OcaLeG+A8LjozQOSXHNdcHnbTPRoYZtjdz6qvryqJLy0fngVM57whGWv9
k2MuAEufmsXyYYubon/RTNsCN8LjzctQzGtvXX728fFSLJW948kUA/fDvRNwiMNnIfbjv4S9N7NY
o97cBMeLrOL/ko6C4+k2URWsSseXXvsF0r/OPtgSkYvhWgnMFa4BhNZGmj0lvYjmeVCu/zblXd4J
y32RLHcNqKi9I5P7+3tpSfLDYQeDhPA2l7l4J/9sV7QWD7IEeaBfECwsP3BtKRm6Kxl3vjRia2In
zixXlbKBAdbn7O1e/Kx7LEdJGi3bK+vYHhiynjV2dR/zgR3oWA+fh5pyytcHAap+dhEIuqVD7Gmc
4IeDOUxSq6w8KU1jFgangLlrUzGUvjhdvKmxjicb6KEr6/a8Mlts5qyq0IEnSxnlVPutLCXw0DT5
i9EfU4W63phS3o8+EHLqXr9fD1dC4t/S8j4LAq3McJboixOl9728NDMUN5s5rHFc6UoDqiIHG2wh
1I+9rPZpIxh3U0zVKirLumRb3FleAjRaQVJDE4q2PVyl2LI1K3kZ5hm/p6Gtiqsvb7JE9t/4ws1+
1oWgOUl0PWuMq8EFx5zNi7S7a4hNW/+L8o1tEUn6KrPwL0M3UTsL+kY9RcwZxsSyvLeAJs2m4/th
QsEn2HVwQu+2YL7+zlqrYj6yS+l3058Bqx/5yUjPe/TWe2y9onfbn3zvpkdSR9kniwIDlU6Q4F6f
boUUaEZqDQQknqIn5O+FIwvYEWwa7TmymWpzGMi24ddercnmBBHBipkMdg/t/lh045dGyYbpMCpw
osJzRfLFP6+MXMvDKtHxEMbK3xyKuMo9u+a+4zkt5KJlBaBZGaQiBaUJSzC8gzvSzGndbVcyJO0h
7o9YIO+UfUkFlXa+FU/jTI4V2XS9ecMuiv8pVMTWYlXrGcWujNhuPhIG4ilQgTieln+ELV655xw1
RkTVRFZ9hRmAwV5iWYb7hcFdBTaEU/HplTTS8BWsscIitwd4tHCPqC1t9B+osn6nrNasEWjSpebF
LG9nkc6PmThThXxCJNSrVU2dcGVggjNka+TP/4iQedy/AEwYizxL8nhUnN5GI0b1wdCxmt625QCd
H3Aen18i1jXhLkEY+0zr8k1H0qpoA8xTjGzUB8fdISHNG/5FySdLO/Mc346NXslqiivcIRcA2Pw9
loNw6K0EZ8qCuPTZoEkex+3kOiHFuGqFTitQwDXagTKxcnM7RyP7DjAwLcEjgQf4INlZlU7qveFn
Sq/FVLktYPyY8s/KoAYGYCQGoutpsHqXp1h8UAacocMg3dzbTu38+6iEttn/P+Z/TbiKv5JHlcDb
amchrUci70n3ZHsFKXDXmrYeZ4rSR+wluFgM7grzLGo1KHT8V9p1xlcSjoMjjlgKlKCIuxGvsDpS
l9hLbcYqxsxToR4NDwQm0r/+wcGT5pMS+HTnLeDmKVuitw2PbtIC3Bi+fjMEI5TY6jJV1p1b70so
lDW56K/3hPPhCH6Kt5tuNcYBZIOUGTWoFqAQkSk1EzUVtescz9I1icK9ZxtR2cBapD47mRp8PxUp
oqf9nfUckXYzCyLJRsl+9SCSlEaT8Ra/r7k9wNVbsm1XYGeaTwIwGtON3fwimnojgM9pFFDMatjx
Rb1I98/fbGgPPySH7IcC8GNyB5OTFUZGTIgumexzt61UmQFKIXfk+VIMsK2v6bw11NKUaDh3bfe8
AuWGKdnm+MfDJGEvVZfthmpwutkn5oUrVoXdEcdyMTi4P7UbYpqtO3IC6StfBQixXnhpS3c8dznG
k18Wx1ibStla13lmij8WHay00RGWoITXH9ZZn5/2Io+sF4dz2BA4Zd+WLMI4J3JEmyzZ1Vp0ycHc
4HnlMfM2Wk6NXa5cEVAMrmIU5nEE40R0iMJly9OlWzjlyfrvHXwF4JnIGO2DxZLTntNTrds77Ua6
Dva6VKiJMUC3MllzRq2YKA3gzkd5U7ztBiFNLJPf3nNppI99JtUIVbGrwsRvoadlK6RTj4dP5mkI
UkyXMLYOpBNrK1xKC+m6/Ro22HGfuKEaPR4YJC1wgcG4MX0/bV61ZIAIonXQbe61Fu59sTAbYaYt
MPNCNfuQU6dF2YOCtUeqUTisceMcn6oYEeejdzYHIYZCOl3yMJBIeaf42HiZq2GoN8lZ0L5Ol4P5
Yu9IZlUPhJjzpwap1rSGy705Ns1YdZwj6MWhzYxUHu3kb8TNnGZXcfg4Wu+2uHoDsij5pcCHf/jL
tlV4AvtniVO6ECvQX2M4m4gbsaHytCcaAN+uMajy5MwcdTtyRi/3ptvtXLd3dVUxVTJ9EOrqeTfe
7qUQxFcjLIp640Nfb28BS4dapkPBZjKNmRSIHxh2jQSZGKHJSRYjSphKbgZPiIPE9TsWe+aPextP
C90fh8Wekl6qvFcJBWkcJWhEJlWbwPafT/tCcP+WfNkniohaWVpEx3Vc5syCOiIq8HcpF8/4ex7g
Cbq7O/T5d326qZEp/6RP3lWEqG6MYKUqXrUA6368l+MyglyEPr7O7Fu4buZGsmDbJMXSApwg4Dli
BM62nsBb4tVdOgLQH4eSfaoCpVMkox1UMeUhnjART0eOGdn7k9DRSFewjKEtHOpKT+HpgC9w9sF7
YVGmaJrpV+UA9nrKFs+fwYWlWLYT1y5Lv+gVd7L8uXxzLV+1ecb2lkJg1YV0QWal2RtowHhUSLb0
/DRxr63NGBvxH8681N5tHBYMSQoeePum0BeLRC5iXutYBts9FOTHT0/Ce1xIF7wCTIwCW85WrLyw
+MI57sKhKJ5gcLutpoeMSo5K1HzRkUxZiK+d/g/a7H9tKL58EnRr8DG1sjoTJ4S5+mrIJfXDenva
Zlip3xYMiY3QwEeQEvBI8gBAHVXk+K8I96HzY4hC2881SvTU0NnldH+XIB6+FWZiAvQVBUpMTY0A
YfCu5aBPbhHuDAoouMQuyw/h3Z+uMBwycTqnPV3Wpmr0luyEOy7w51BcE2aqrMrMbZSj/vYQFPiN
Oa3cZ/oXbhw/y/SB20kTGjBk2zFykFMA5VHLx8kFiqCywzoteXua92A4qHDGi8vPqXTAdV+RVH3b
aKbJIr4yFeoBIPydXucHsbyw66VBvSqPJ4Zn4XN3k9Z85BrEdLzpcLY7d9O9iEpgblRbuztxDB0l
BaB7LXSSgmdDqUzuZHPW7MC8e7fkHdMHFG2Rv0s4XyTG8DW4iwxUOM9nKsgy4FWKLUdiIWJFdMe9
HYX5v4hkccj1J1e4tZRBnYAq5Rk5s4rcoIWAK5UR72NXK0YWOQZfUOG9r7eQ7lG3Eb5hd8pCr0Z9
X7Oaut9uGVtVGehOXjT9iQHGDgzHiSYsb/XCdkHtyFacjuL+QODWefuvHnRk/1msTLIujb4jB7gb
E6Cy93sxbSDUAEd49G1qCsthS4SzX4tl61V0Qwfm+JtSGOg5P3pBmmP4QWnwBABhbjC1uHPy1u5p
CcMhXsp+kSlcyy/+rh/qK+Ev/C2FJLDeI+omRXJYVis4+rNySOxe1R+KcXbuYhmvV/JdcWI/tlfv
/sqPAtRC3gP7eTElizqTMld2Ah6iIS1ChkPmuFBLX7pokyY18qPGM8Q6T8EcXJIYmpsfyR4EMzXM
eBreHPVDViUsMmNwWy83K1Y27sliQ4mMzvyfRhBWCrX+YuaTzjt5lIx28XjvSCx0OriiOI1YfON7
aHbf9Xh1Sa95totN4G5RE6P8s8bCwK08UPne7AQmfVDJEI5qOiWQoZeEjQbQ90E7z5SZrLeJa4D3
BkVXgvMLNKFgZrMKEaDRsVJp2VyDK2KBcaE7F1Qt8GHQogud8ZSgZzypqpCqJn7ZXJuqaXFi7YUS
NxKTD1YKf4odpC6SeYWQczBlKsv6FO/5jOyVHH5FByDUgdI3pziQl9rFGfwrxeMXnjeuOoEDDhRJ
EGjv1d9kWowfLopqpGO9GWMxgo9h+UBBMiZf6yjHDs99fStZe78hMXFPJYhEdvZ2NI7d7rnfsVwf
Zv17/LXxLaJtbHWBVtf4pl+2S5DOUl6vLzoZBTEhEKWjmofBtlOIz1EKR3BI1r0TgoluS+MfvyAk
aQxaPmiXtEJ1tJ94ze10XXX0S8dfv1ioo7KgBvYKnX2ewouIdglfOZuxauZGbj3WUw2TJPeG94gu
uLRoYJezMTI5Nh4KO7iw3i1XDKEqUKTxUz6FMCiP/rHFau0PMmS7FQgGwrNgDH4IdDrkzG7TF5ar
Pd3j6ADFzQ47FJhs6V+JUyPh3NDg4mxtjCcuOY/5hGu1oaJlDeFlQ3QaOSoOdB6mz4zQkF1PCDIy
CKaso1jjXxTX6vdG35e9nU2z7lbOf3xCRpBs39PcI9Q7Vg+a1it9alsZodNmJ1ei9r2IyQLso7+j
HBHzxz3W2OJbD1Yk5iISZISZ3bofE80cMUTJbRdRxQ+ZPZP35/U0L5P+fVed1fQOpTMpbKL4EQkQ
Cyxc6EeQwUJKY/y8cS5yATT4fsY9gyERf5m7wobgG++thbRnFPANKRvVEw928K6rlg0MhiK6PwWh
I28a7wZ7qoTPUNDFnDmo71DIlUpcVdlJ2lg4o6EA0l0GLX1DueZ+CKTDhcBnCEibHJ1D98Dbwnzt
OXvum7kQYhm8LwoJRHLZZpXpdPLNuUrw3fRtzW3Kgrg19ALu9hwMXyWTicRUEOvsAE8EB+G4W1UB
0jZkCBxD3qDpVc7Ci1DR6C+zi/qJRPk1ChOR+8tqZNs1EIykhgPnqvbbnUe1W1ouUUsyobTHUASK
HiOX2M53iGsVCExmqwUi3p94rCuiWZ5WAumqhcbTS11QUUFwEHU2Vo4XUHeCsIgEA8H3UPLCLHWB
zOiOMs5FYalngqpeHXeNR/tFI4cyWRujQn2ZKSZcVgIBdg9AkD4XHpQpPL93oYI244VzqPlmguKD
CAf0kaJK2BSMEs82Ta/1xm8lTFx00dcClFIKGvMiHdStcHhu91/H/oHkt5sUylYw6GAkKKJDP2BP
VLl2qb7pt/Cg3FcExLujyWxwDOVOrGxm+1z7bUdnI2x72jxdJ5b1IXZTMnpTI47TaKXLNA+tfTn0
fMdXYQrJ7iVT48sg9oUrBoXlVfRKP0k7LiOxeaf5xzhVt1nVcUHOwzEUZLkZFHr1kgguSLtBM+Yr
fKDcX9usa5WvEpLlqFCv4LN5go3jQp4AtIMTge3lqqWm/qqlVxgyc2kwcSYKbmA+lhWYkRibydBo
3bws0lc0Iaknk7Phley6pfeF8UhfBagA84rHbWnbhWyzfJ4m5X4OgynsLrK2lgZo+2JDO1yQFWh6
BV+DHFSej+AKp6EH4LRm79qilIUA/AYK5qmtCey3eFvorKBM4ZNUkmxta/HLhI83wu/JBh307qDT
qiVdbnc15wDNL96zqeuxqa/sac/wWcfK1Hi2/2PNdsE2Xrm6GPbLCTsRGC9sNzhDoNP8doa3HXa/
j1oar/3bmdq+MpFMz6OzvyO2yNLfE8Kc6kF4iMWIywRQfczeawxVt5bAh1sG8MFPcfzyQPqkHimc
+NZO+3CPV56vdeM37YcaUmyY8dL566KQpGyg2RvackotXdaRnFTOKE99+PWfVJWNt/CvmRzcE6qE
ML5Fg5fUlglFPPBIpHZ9FkcsK0QF0uV3RKuH+M7DOLDVXffkYjFBEwHv7pfre8AUA2aNH71Lmnz+
MdgnO3QqZcXrMvupV4sDZVnmJ33aYFqWXhKvq/ghxz/vNvQWYw5J92WVSgU1MedVcsfzGXXEQ+uU
CpSNTaP6x7XApx4Mzflf/yOUL7wo3z+HBxl1cLRKo4YJyRsSaKVZksrPIMSX9mfbrdkF1i1sF7Mt
B5BcgZNf4Kn1DPJ9OdawcjsXKjeVRMrCHdZBfEq6X7/730qYmeLGHAJAf/C4WErywZSiXyu4yH+O
eMF/CtML1eT4Wwypzx4s6twUx4/LsBJL69u+dME56tuRLoFNepVB+v85uIjM6qgwkKuXiU1CHNaI
t8eVotS0/37A8tMGODxoITqvfGodn66TL3FWwl29lyoggQDTrtjIyNBy41IgE1ijA8NPsfddeD8p
j9jp6+Nj8OM/zZnlIIu1qELl4eQSBNXG2Yo7uUrY46WJcl/lSdyBRYGgJjpWVu3ZdCeXtXxPvQoU
bDKrw/Kr/D8mhqyRjxmc71wwQjEwTQvI2RLFmYB2Otl06Poy0ULyOZCNffMum029278f+1XDxFrY
CY/mm1lt22dJfm9ItJ+YL1ILt6HFdVByddxG8nt1c4ysAAxBwD5YWJsIMak1VK2q0KZb0TK9Th6R
BoH2B78/Guyw+1a5i8OCE90VKsz9/4wtpH5op6P1lzx/ydxHxPJXDc+7sOBGysl4HkB/2m9Cuafs
GxkaYyZ51uyskDCRKj5BlQrqOB0a1gSsRUivbKqCmYPsoaY2hfhvv8L8NHbXVqAFBTdnK1Ci7Jwc
nVxjrInOUrl4bxfCh+A3PRHPLPogilTCcZUvpKKvl36vArjxUDAKsHHRoAIo8N14bV3TY6Zm4s1E
t2961e8WwoEyiODwqxPEQBWwJmTTsTzpJ03xjkldansiYysHubPF0aoLeTu0daPHra4N5eK8M+Xb
oPaJdobEFWzocZpjKOCif4ePFx5WK5tzUaAUjeO0EewV1A9ZBZzLt4QpNZS3C3f0t5XwKBCP/gDn
4MHY5YeXIeKp0ucxJiev0dn8CYfuf+4lVHmnJZ6BjKYzRlzKwav5EfwY75KszJFBTdT4A5S+r2n7
oWaXXZes7tLektvdVFseT+s1QcuEiNPXgcl448L1ypJVZTEJ2oIXBl1b7zOMDcqZ3iCQkoyJwlOq
ebyzchjV8M1XaiYTyBP1TRKLnnW/nlXOqDAiVeq7sPFlac31wPnbZxAHIq0jVMK6cKB+QpAeUYHM
y2uJVW6jgMI6qIlk0VmFcKXLvz1vzr8FDl5LoERTPh5IAVFJjqiaYMlJaBXdopFTUc01kpzFurzh
vRSLZv6JeHmdJ8DpuXKxAcpCxtN8uFGWXRV0O9ar877QqxfAqRP1cDyBDfEyMBVuS9DDzV211AcQ
mMETNApXtLauxpo49l40sCv3B8cDA4ISNewkF7AQYH7OmjfChV1LUGn0cztn7h0o7zMixKxl3duz
NJDuTIxfu+fVsO/M6URopPPz95I6EJ4BSA6YlGeah2+lxIz+r+5cQmKSfspkv+HKDeVPQQMQh9v1
e/Xkb7ukouRQWZakOVxbPx7bTSEozYVplFzPMubHnd/JIL+Ipvdelm8TjY/GQgqaZeJJGj7wshP2
zfM9CJK00sEJ6wHiPPjEKoLgH5PFaG2aZqKm+sEoBdonbYs3QONPhPzPOnqdHk8R+1K13hZVlNpm
S0NPYTRnMKi5ULYpFpc6iWXxh/vzN7afRy9fae9I0A+RdB1P+xNGzYs7DvjbOmqyaePohVZ7V0r9
l11h8QzOtFyb5U4ydhexUWnp9vuaFi5hpusIYF5OoGBkFR9dwOLRVTFasp35r0LGRp96yN2Ur4dV
gZsSTIRL+GrPkGOSXcn0ZqSbTxTBm5sAVyr3O0Pg+NZ4xOOvzvGyn1bFNZHeUrO4VN3Udws/pOTV
JfMEU4bM6Y5dnyeo6r52qwUjdpVnDKfCWcorAXyaZHYLFC/1p2SeItNHNcP9kRJeKkd+ExC0qKyX
FU/uqaobZmzqEPAwAw93moCDH7Y0Wm6kl2B/Rq1uYvVvCPZCgBxK/s9PQ4iGVioOWS36nXnXr6If
lRGWbXypLbqAAvjnLUCdJJa4b4FQeG8qof7uBOYHiKFEAGQBuDxrcaz/Yn8OuUu117enoUxVDyBr
85M92JgH/f1KmfP+gbHLzwVG++/D7rywElpKqdgZ+17jCascGgbvb30NFySnjjLajBmgxB+YktoE
NSPl1j3UB+hqLuIBE/Qr1mLSxlE6qcGhuZn5GQSO1uGhSx25lkhewN5V5OS3zN0WBKHSvjb6vfDQ
XUVKnMNnvq/VniOxcvkntCn+ip9RDUVLmNnQ0VB1uSFywzpAm6wPUL9TIZmDfkOdk2xYh3hpFoIH
8jwmIALVKCjuTgrSm61+KC6QsGudMkhvEQx3Etjlvo6YJVhVVsAakX1+tdgk5gebGHdfcYoyTT1T
lcRbLIx7ZXwr594QuYXfT/wFxZ+SMUGkkETECQLIfzrOGcWt/sw4T1K19yNHbt3yk5L1fG9t3xsU
gHYCm9cdmeve8ffT9YEK7hEUzEmuam2IYppDi0/UfoAgWfQHKJllkDN6uBM7OAdu1R6zP1FHZSTq
CPRN+wQ9FxShLgFLG5f4WrmPI2ckarnxt+Eimr60yxxDHUfLwVOYWs6QQ92K9ODMNnmzO/m9bYRX
HGQ2OrQ7AzZnSr58F1cgAqWYcBEdO+s1ONuhuDLQTlPxTEiHriPUR0BVXv1Tjqzasjg6nIJy2fBm
FgQyjmN13G1wqDOj2c6Y2Xw5akVN2VdGnsGBHedUE3xOjQtQYfZwnldh6iIIpISywDaZ8paKtboS
zx7AnU8TacpRfFDvAEkbpaqBgCbT/f7Y2kN7dC9Za67j3zcCPICiYpL9lFoWG3MqKsrECD3Q0iX6
lvCpUrQgRCCePBlK0ORoPxOBzvffTyRd5JCKAGVbiu+p04L+ix+C12gRAPFHr3x0fbSJhQ9yO1RN
hgfAk343UDsrf9jLwNS6rct9jBpCRHTvafmsceoImNz2jea6+Po9RqLsYkagh7WTXpqE9exsQHcQ
w0huvBUga+uBH24n5VK98CMVg5csAmy50kFVFyEwtP/cyoqx+FlQJPBKFQuveHpvIRijFEDfXvaM
tVLTOlWOpV/r3EGmrlUyVF+6zBuI+lNhuHAHQD7X73s+LkND7T4HMzXau/txOczLXZjeiFzEu9xg
V5Uh1SOo331p0Nf3AgOKQXENrfXcRKMO+bGVoKr/rKEEYwtOoy/9U1xIqtrMRcN3znFzdIyZ4g3d
h4UyJQzvogbDdPjFkhRujYFdFFP42sseKhkhEALm+4XJYUlZBzYRg1jzXsDdGDCC0RwJNxenrFNF
rTaoD1ihHCEoFF0KCLrqZNjauTAghCGH94J/FnmWmfnf51LMJemkSOdGkb+iL+y/K3V+ba0Bh90a
tL0hL8gNvYnbiZJM1XhIfLdZMB4OKozXY2bPLJqqdVEG5oMqn0cgqo24I0kgCpRItL+HcmAkcy1r
m8/tVGGnw+APEbcjGMjJzNgA9YKvCZ4jDLfPf95WnRxjHz1CjOOogfzl50+O0psQH/ing6xALT9k
XwAkCElMQCS+o5JLc0dMS/blEhiacdqdKIniuEr+s0V45t8zczY+smcmPY01uW6CgLe6rs7f7vun
at5kLpS5Oz6yi8tf9J6SWuLrOyFYwdSQE5o0FZT1j1R0uonRXroZdn1uHBPEbCRCWAdZYlpidhF0
+QoUiqPGfH7G4dd+I8AjdqvHSt6XOw+MryTAJ5weBrPtoXOCu5uf3LUA0n7cJnHN5HYZohwnqGeG
a/dPHgwMTacdwsZgaVSaqBsz/EXLD3PhpgYESLqSZWF5h3CX4etswWPjfz9jdGoJIbZFZ/sA2Yp7
8ojRVSQo7qVosLPXEjjqmXQjIMN0fk8c0zJ4Wem0q5XNesk6wNS+4GW0PQ8bY23Zda9MlXcGl2sI
qEaWM1XuGktUT9fsm9erdQRaUCNd5Bw+UQBSAYyZLF7TjhvnuwGmch0RFytE78GNxy22lJpymVZZ
W1KqHGX3B/N3hKUyHPp7coTw0EbgfUR4M9Ygo4fh+PfOPEgh5G0C1pDaoibfEuo8WwkQ//WYmLI6
Ok/7Bo437zxhfKQZ0voMsQe/SWhUX4yKGhrUEcreziAWFpyLJ8eKrWcDd8yeOgT5X4p/6xXx1DPv
bJ++nnoDHO/Y6GiCBCmGNJjeI4m1dn3e8Fx7WBvSpd4bItFHj/1qI3sj0qV9kapY8uExSYW+HfXt
EM5M8/2/Wy+hFwO1qGxzv7gp7WfGQWMGv7G9kg1FufBG0mTmBLanLb9UFdasYteF2dT1mkMgaZ1W
5XtHjYE6UvMFGNw9jGSm+JwFbgYq2GAcl87MyJntN8bqJEq9XD8ycoF3moF4iwpF5e4rDsaDy8AZ
KnjSHqE6vAQstD86tOwjSmgy7fqPv/txz7kfzi9c6kFwgup2wyQFo+ZEc5GeywHzvzViosTZgxSI
2wB10z3gUcnZYhJP+r/KRAv14AKrfoTyG0NwzgJuIZMYthRc3WjQ98YKYnzPOzTjRV2QEZOz73YY
9R0j4tlev7tjTjVY8mUiOA/yMkU9NBWCcTuNlp+IpeVsamY61gsjzdOQgAT8aHqsbtpbKyJwdet/
q8pdnRREnXd3BzjgEjqzdA2F9ZjY9RpzEb7COAB3dgGNMhmB1PSEuZK+j6LipAWuw1uf6lNOy+wc
Nx85Ph/AYkEuRR8rbhxD+RlTCtmVjIpvockemKnzHZoYP6ATxkMVWTGj1bNWAH250717R+JozeA4
JbOcFXtGgaJ6dQZCF6bvfadPK0BtA0axk5SNhCcOGTM8Wf8KSqUFyEwGyYwdj+XlJGkTSM/yn7vy
pw6YLlxczL+U9Hso574GUuAkoW0akDB66dR/OfnR2rQXg+E38mF5eEumEVT2plPfpkJAFcC3Y/KL
qr2fp9vI2nvAQ1bYMwJl2GqRIBcJ2ftCHvdzNQaRZVFN8aoXl2ZLLwgyMQuJExy5WMNdLNjEnyWy
9OfVRdjCBD+Ab48X4L82FJZ0cF3z6g0HVCYOSQkwbUn9VkEqIMMyD2qsQq+9bf7aP+QYXlJcww8k
yyPN3u8LWKsnwrrNM3CqreSkVD5z93sw0xHnW24DJdWINtAu3G/yHvL4mv+k5URHpVDyt1f5Fxep
t9f5PorC6LUQrSrF71Jwz4Ji4iue7dKu05/Y5QwsbRiqEQ2IKkStTd3HvsubOfFx7qMn0fVsvhvN
M+bl5LGCTy7lJgwkjSbYjZIvERzR+2VW0e7F/EXQc/xvjFBFh2aMEpnG15sdVGhVVHur3Sl3HyYI
qFNgmkX2i0ex/YnXmGHY9zFCHf27ciHQkaOfQSjA2K2CHRv8HF1GTxJ+r+QDWCa4U6vHP3X3XIWU
yrS05beeFLlD1WQDkww5lyP+r2jZPZh6Kd8ulfbEsxCzV0j9T3lvwVe7j/IAguBjPrlQE4afpXhk
7aMQ0UJtP+QBRP65BQioaBXhrWr7H8s2I6boQjcV7qdsh98toNyRdG9A7QBuCDj4/6JzPJxAj9wO
EXgKiLkW9GE5TSqpJBJKlZnqn4lb97I+1eDIJDDBRf903mGlWFmeZjinFOsl6nSYFVvUWsM6Vypc
qY5x9FZt0aKua299IGkLp1W6f2/nJHTDMSZeKYUSFl3JGwmYDDdM2kFIjUqaHby9VbF2n0DwnYiV
OMMvcM+UfzQIjkSIV0Bdk1WYwJvCx8XkN07778Wvauu5amWDIiUt59YnsnFSpspwVnGfCZZMlBL2
YYhNyTZTP6HW+fgCPcvFvPIDBXueTi4g1Z3TbzCeCb6h2Y9Lwh4FwPz3q404vkCQiMFrgyf+VFeJ
fg9OAIQ4SuCY9xN+3IH73CKP09tkL0u+Dj0Mj6HXbBQ/jpirZv9+ln0GSSOHFlBzm5t37QeHojyP
drMjjo/MACLnjY8nRYVMAsfBX/V+gtCtf3ybHlqhhwBsmeMnSYeErtjeZky2Vj6sGtgLqgRoQlxn
fQuldyEhEtpls0gkKTVFr1ysMTerhpUchSZg/OCEp42KXh96q7FcRVuT6HYmRm4BIqY+lCgGch2p
9OdBlmCrxB5Py8qfZwDfvQ0X3zdo4NGwY2ghUvKUc4uyx1EkPUpry9Sx2gFqKo7lR4B/WEHwPdPh
bcvvQE2qdx8iua1HBWhJWXWaavHQrv27yPFQTXmYjjMIflZmeTyke+RaeNIqblc7qqBGhEwuD3Jo
caVtWK9azLVS24w9a4sg20jjs1HDtHx7arMo2AaF4v40fx25uuoGyC6Pqb7plfB68o1wU7vav+sa
2w9psJ6Y5V9NnisjBNwoT5yD2fl1IKIhBza1uN8UrHGi9Erm7/puYy0kv7y27QMiBg/vXvx2/pCL
ClnYDtYTUVNS6bLHyGGSXa/sfGb7gjz2xXzTqQ/jbCBiEky6LjNGp4/Q+MnVuDZ4YHnHZwkB1WAj
HgiXMbSJxknHRCsCESPF48Nzj8u/cCRftGf09e3AmBKiFwlIcXpbif+cmttaVrSFTCnDcqjVgmt8
yIvdDocfrRfKWrn2uMlGz4PZmM9aSR+adwe8iDXL8I+tutzaLqAVF8IH6ceEYcKO3ZGCj7ImwXqM
mlMZBZ679piIG/pqtJINGd9SrfB64+Uzsk69lDyYnAlpKRGhkLIfdYplECBBdXsFIGAu2VnTWT73
oR/vVn9itAHYMcULcoxxFSgW46roQ80b5d6oYemfGj2hHMWnekZHjZYm6ZvnFjg8/3JWGRCYY6xv
w90BO/RbJaXUlRhjOuEDYFW/RAaMXZ0l+dNmslP6MciaKXQBpubQ5ojivn0g39S+0F0RfQCt8EZc
zxRonUZu3CKDC4w9NUzPwP/abgBn/AYrbZDleyVI+CJIc2N+lTpRjVPG/QOIYy11HBIH5ouQKVcK
U+upDIujFRfPqUbqxNyCnZxYGe1PX+yFJuSHerc7fD/nNbPlFIov2UY7/FSUPblAvAmWHDzF+W0D
d3j84NbH0bwdMSO4oaq74DMeW2toit8QCHJEUygr/FYRcC60b9xiENQSC3FTNCUPRj9TM5qk5ky1
qEl7727KT+ZQ7FVPudaCjZtkCeev0VRij8euIl0NGw+sxyjEpCx4fZXQ8OZ2QJKcdfGvqtZmpcr+
MEUx1k6m9v5pDxmI8/osNWbnJjc03cnC/6i6KaQeOajnfqc0o3JudZERJgvAdXFdn7l5DJxSkFEY
GN84iO4lvHB6P0VpStdod+y1gwxsCbGAzDWkAC0bDKniqQE6nLCf2ZBS1RDcH/KmvHcToTnF+oDX
21hvLfn4w5qD8yj/Y/JMUTHyliFn2x3d+pAUbjGg3BbuWxr8DBwOkeRpZoBLoMTz4lJTlfptzXbn
lB6FmM/zlZ6lfeW9hVPYx4bX8mpom7MGyYvSQzKKOEIIvlyDVoXQ99DAjziROk+sbgw10wTQhmQE
y9DY+JAqC/48DDNae34G5MXCmqp8iwfvK048iMyVy/3YLXYMQ6OGMKey3P4n79JJWkAG/y1LSmeE
zvfZufWH+0eAxqtH4ZU+Rn5MNwMcu+76RqojbD+iJ20JjsLa1kR1P7N9NB1WCZXEhvJz1YRXfBBF
G9bg9WI5637SvHtVTRLZDB8/m0xvVzL/E2IXUGI9vrv2wydC00Wehc94uggs9MsIQi8EC4u62fAM
uRsqI1Dmw2EW6TBoDglAmGRLhs9dF4q8YzkYRhX3B/uQBQGBsUmZDN/bxw380s0FAjK7Ijer8WEP
/6NjL/KRxSmXX7ncox/ahwBNjVMUdXs2NNQYKUTizHVFyHtsf45LlFOBu+fxp0Ej2Xr9HcAbXQhj
0ud22/46COdmqrudVfgVV3GymvvgqEfxmAtrKE/ChVeku2NjQ1wXhfZg46qC4K46v5AlXqjerw7x
eTSQTJBTJ/SB+EkuK0leCmLIpEWtPMeyIkbwEdbtppf7QpYt/iVm3ML9IOI8ZUilh+2kRGtIYFmg
PmDQ8nDttzIprGMzlG+LBeQ1nXn5rp7HmgseVyTyP0GXi9QUKXVFbC67oaRMRGEnUjAAuvmwFz5R
dVZANp/fSYZqQkWGA469S0LXM0IU0xUlRepDSMELBmhOLvf1dlQxOHHyWT4CnAmzqLMfx6zZnRXA
cNxdR9tGoDB/iFfBEL4I0rzW6QxUDPoX7anjPp3EYvx9AhvwajyeQwwyqnyYFXgHDow2G7NBYaG1
t7VMsNMzwHIuDhgG8J4uRBCmDYgHJ29oZieFOXy1vshCqIm6WeaWo6G7Cv4Q7DTmfno5t4e1xObw
iGHT5upLEymf1ztWamCy7tx7a9pxfByksToK36ZtM3yEWNK0BTZhhLdD8iia1quu6E8BbCOnuq/Y
yHMw2OouRokvWnL/VpfKI1/lWGrGOuxAf+zMLPOZU0nm8rUj3v+NWWC2pT2e1aJ2ynhEcNMNiNV2
gwnWl8oUcVfkBvy5KryZhHTYJFjoxRBd0igYg30PHRV8jgyND+f70nR9vJ5Y8iGBY6VPN9KsBjsR
QNTdsImF2qXvRLdUQKsoVt1sSYXSuWbDMpRHtd0liqHmG6tJAQQttq6sKBZQ/BlixdZPRpshfq1J
j93euQ3MRY4PftELR1UnJvbbqmvOmbFD+/GgaeNzGyxBuHVW4VP/TfYLAAcCfDJvQoWbjivBVkz4
rVKir9Bqm+W4nFUHWXuZb7zMiXe04C9wyH7O06NU+D2/RppJuqqZmA99wzibSNNi2r3q7MB01pGs
zuxdfHjwRIh8Cp1gorHAxa00XRHsl+k7bpy0A/b2er8OjVEmEOgIsURO1hKWyxvf59dlbEjs54HV
6qhnaYpujU3WJfTqxGy0rSnzH2FMSlbudsakZ9BAeYMGQdNMSfEbrHKzT2R0hHujM9C0euU+JT2B
8zFxbJFU2925tnFYuRfesiFP/QOkeMTuICSazDC44Swip6ye+22W1BSnx9Zr3gdOMrYhqVcQqjTU
FISQ3ZRb9tRuRp+nqIBj/45A4mZoR9hASP4Zb+yh6s8C8ESDWTxcTFPcqdZyMmHUBYeuyaOZ3LUh
HzfEQqH7eXca7MuAVp9m0aUA+G3xyuQjv5DMwqjWU7UsgDWSwnLwK4QmcKHiu7xYsicqxXQ/kuMo
gOUryTx429/vTLR8cUyBdX7JCd2yg1CTyvYLFFzs4dsFtOGi3dGu7TDSgTvbj9ojH5BhCIbnNOQY
3qg2Bnxm+RwE1Uh0/RSEul0RuJn7J5S1Dnxby8AbQn8131UBnAjdoh73j97CVZQv1bqeUOaXKQvi
aadCkvS6zawSnPweGk4NPGT8N9aQopu9OYyZCSNbOTRuAh1AufQPXd+CmcPwAXVaSV22LZTqfzJN
ddbdrzKkyJe9vNGhuhN0FQLOWqT3DAGWPyEd/StBmgGn2/77lEBU8K2CbOu5CdjSGOBiYc7xIAei
UOplzw1T2W3Pv7dCCqx2s1gs/0TLpXrUU7ynAliHUvn4fPYQVnkHpv3kIWCWnaxvviH5njc97gza
N/Il2+Ynm2A/sT8GAjaaxwIwqeHa3+kT2LxCO0sjqnChOI6zihUU22VwVhQ1v2EqKQm0Y/yYcuwV
D43p7ysKJds19pMxG2IBDBeNCQ1m8K54WDvQMPH7FzgkAfotHqkeuJQ1quVZZqBbtn5joJ/gCHCv
Vs/IQhXwECjguwBxuzvpx3V3syNQitAIb2gTpLkVpeViP103XBQ+j0FN1hbEjBKTlFAWQL1v7a3z
H8i3pTr2ftO7jqk0g2z1afm759lOTiXbWAlJCRHXY2OB+pzrvg1d1sRpPo2UPINXw28KAI7eELGN
E3YpguPTybZrQCbP1bHNRUS32LXcnfy1SCwG9WpBREnav84NaenjMaI/fWFC+auNyu9kGkwfv55f
NqjTF7Ko/45Mn+icqFeRMIa4hw5qHV1ZzC1cswQsMMiiXTrFLYdqYhR3EektS2RYCwiy9qF0d68O
4D24d+OwaUe5qZ6JG5B3kZrxTHuZ8rk5buVO67oC+sAUtyzCmlqAALMew2LsJ7Hna3spGuTbaaIJ
aZh3TqeWZaphiGTBOTl7byMsSL5Zh9YtAuuC9jhd6p/Z4Q/qiVhBXv4JmPjnsV/smQR2ddODoLN2
U2tPZvR+6YO/EHDAUbNhd/sTOc31oSijMoC0aXHRlG5yjadvWt4c8C7vGuhXbwv/NYQU4bjngOhG
k9pmvk7TSBLiHmT3qstsoOV42VSpj3JdPPv8OEKFXIO2C7gudzGBPO5eu6guvPB+ZpWrG60T9Knp
6OhjyH3X7ku9zOT2SILssE9lGzZU0SbsCCavEBoijupbNyUXAqyMgubKM1NdHHgbGEwmXPPaP6IC
vgmlhPSDVQLiKzPZAjxmvme04njZy+Q5YvLzRPIx8XqJJ8zZXFbcXjVgasBmZIkdosBefiNx4pjs
G3PYz+JVJog8//JvUMuE1GQgstUtxdPElaMGniSamVLXJlSEfJ+FOMLmyGTpMPrSuYORLcB9IfnG
VzwHcZYWociAVEF92LY0iD5AS7LWyxz/EA/IJV/D21/rYIljSQo2UhCuxSYdCJyAlsYDhxwUfj9u
I8O3iOh8aQJJgyo3iQ9lmMBDDkydCjE7ziRZ68veejDOAspIis+Libtmx3XPEctTzGOGLyyol5dB
MA66RHexvS1jx63tM2XYPiN2eqDq516LqFV3ZAL/+g5XTLWCizNklxAgcglEzFScI0b8nsBfMR1x
bUSH7hC5uX0B/FGT8PMvIiETcY1+lAg54ZrR+Ard4Zz5tiB/j1oYA6xP1e8N/c8GoHB86ZH2V3Xg
FJOJ7nFEmBccdf69DMJWUAGKqxrY1T33z5iG0FT37onblxWLfBFdhBoPY7oxqT5lMWE0NoV0tEWu
ezyLOcnXACbny2V+5C9W5l6oOVQDKn7EgKoNbCs4DOUGmk5Y3Z+PrnvQMQ4XM0WXPdxisyztQ7RN
I1PJeQSHbSeVCPgVg18saVN464WJGEkVeYf3w8QgYCqj9TsA/TyoaGws9+OJhVdTxlpVHDT9d1Ey
A+Ky3WOLIHj3ulwsCmfzR5gXjNjLXCTE83FTozjWZZhPU/Ukzuv6rQWj6ocg0XMmS2yFeWqGg2mx
iUtWVmWZ1SoQtdFEvysT+5ROAbERMMyCb3jj+ZXaDMAL+oz8safLmpYw/xJsm6cu2iI8RWLdHCfT
t8vIHPdh0HEv2FgOkjTdIxi3UwgZCA+sPqEfOaljKMx9rm6Ekb8wy/NgE2AYr1nB0WJk17NpjIx2
Sxmjy0PqIy6xKAyXv7nBbEoDUPyJpnmZwpWWOpQYz7Yf4CVYsy2FF+2miCNZyFkM6MR0HvTbjT1R
9Ay56ACXiOQWD6pwOzn3yuIx9z9BIj52BfnUcwcko682RJy0Ld/SsrQkPcoyHhjOZB1xuT5TF+8Y
XtRWkkLBdwvn4N13iYIcTPIeD0/2TTf76vvHMw80+3taFupCClDW+XRtJWYYqQeA1x/eBB8nAmXL
6aHj6S2sLJwHsibtxRnydqy8tv4Pg13EC3oxMASBMnGETupYn3jPa56ueO4VjDn73VGYgITKjG6v
RKaFT+I9aV4MUYhLe459EDswEO9HHln+YPnW0NlcCGoCk9GwJuDGEQp25qNU2p5IqhASZGpcoNcY
Yf1VNN6noQL1zOSm322cC7LUMY6iUSE6zUHaT2FpAo/ebzfNN1jIPy6cFuvaSqgNUDdgiuLMGYDr
xR4svnpeBAgrTTRR/lLjU7Fw2/Rt1k9DWOvQOs8YaDNqXVGq4brhAApVyg8DnHD/CjKuWW5Pvk/n
Lom6yeTUUtZ3c5Kzu6FySQFCjlUaGenjf86anBw5Ssutrg+YeRUVZN+93VY/6sujjTXjlKu7znCN
3TSBvm92ixZsxisKGmSzeRZ/3IUtxDGScey5pSGX6LzteyEkSzvf0kdRN60WotCV883KPW++G/uQ
chfacz9RG8GqwPTh6CEVDPNM1RbZHj0YxhJTbH+XwrtlbHSW9TlLxuA6ZvsCSUxwGDFqURKCYFSs
tEpp3wqTrX2ulNE6XKRG9qzvuCeRW3lTRJJMd7hzE5A/mwy2NDZi60yTbxGoZwmCB9V8xJMBcj9s
31OpXPXgvrkntlber6Slo2UBMCvQCSJrjl2EbeK0ed62HEP3Mw60OAHA5W8UuUxpYLhoPHB+lE6i
sU+YYFUUCjsA/1uJnnkDcvNeiTR5b+jzilOyRLSLno+rGlS0KIUFNSbPrNjbwRRf2md6WRqEY+fY
E8rCyn9mvMSLg+2xTVpV8O7uKc0vNMEyAKuxT4iu1vryJ4MkU85dwnKHvWrNZ2Xb2uxIwGCMrKwJ
jFy8O7MjnSl4Z1YPT8+Txs/f3u7hCa/Tpvu310PKDSz8KBNcE9yD7pHsB2vmGgO7xTt04Obdhxys
9yodzb3p83zdBBqCsxKAAkM6X3evhzbtYjrztaeYtSVyQs9+CBIEXlM/jH4jU/hyVjk2Snvb9/70
K52JtHMkXsWWoHTk8TvHpZuolfNiavx3aSyI7qIBW8TbE3eTPE/wU/oacpxdb19ElUAUbyRuELZa
nW9LlVHENmvEZUxBB7BYXsqV6WnOvIw9C1Sxb5o0bep9+6KXbiJXmqQ7ej4CjfajJWv6JqrWQZJI
bsjll2/AV9KZbqLdngOIHqwnbfeUR9ZqYelQtLkNkLI/d2rjgjcA702sabRKiX7YhfDGJmxmESGH
OeL3W3t6uhQ0XhEbwy+PKCrt3U/arhs2BZEDs+U3rjRSiSQXJCHqXBE2HARI2S+2ALRQcPBcnJ5G
x8pSuldC+Z0ej5C4YSQAZFDtQxSl8wblY27dqTLbbkR0ezhsjroYJLNhrdWxEVPtgJSluG88m9q1
ubg12clmT93xORptCvKboNGy8Ofyy3138K/iS0c0DiaaztmLrdnKHDmM+M06onrL7BTZZepbtfuy
QAK4ttylG4hV4DJL2NqwQv8K4TIbUMpAkjNPV5+YysEUNaa9v9s9BlvTh9oxc2iO1k6zAwZ3ZGlw
iaX3u4vyKFzXUWvz5md2LWeim1N4Utq6sB8m5/s3YbV6Wf70BQVmFjTDT1PXpItnJIxWs2f3QUSe
+ri1Y3oBaFcYHIhew7lozm0a5M+zBmf2U1sKUM+TtBVL1MRACMQg14MeLzwutA9McEiLNjniuDiL
AJqIcSzEM1OoIhLZo7MaWfOTBCmvUV6xWV/IUJpInsNykXGArcbticzK8XP0xVJKY7NB21LusU34
+SMkCeJqgmxJ+UEXT8a4vcXYTkM45jBZAyGJzM3O+vXjNNMMAeZ/+NSoY71CUt6Fm1n6qIkW4ZrE
/6DxZCmNzLtlVw1VVNljfQ0V96m0CsWe9CvUIUDvveDLUFvh1pvgi5P829NEOMHn2zr/BW93hsgB
TaTKVRlE5GbVLur85qZgs9Ojj3kfFmh57ql5wcFJD3dBon1DchrY8Iv+cBm2nmlbEccNYZrBT79f
xE7F0jov7e06zJRr1nn+y4FS/CmBC1kxS7hTGsyUUcU+kvPAa2BJIHXmtam71hcWPqmmjylz5Fq4
td/Qp85Om/Oqa6l/54skf33WAGehqhPSRvUVId/I/04FSoTeaeJTM25ZJTzaeeMeRkhcIX0ItWq5
EGwGv7E6cceWUSMmK+qaiL2Y/+Pv1uJjgaSf6FTw4/KycarVs3VokynmYEdqK9+EMyUYuJgfZ51Z
Dl2sM1RRgRa2XoyOjc4Tjy1gk8TN26EMrfu4UvAQKNxoO61SEw3r+qwkse8YcHKohD5/k12JpSc3
b6pd0ji8Vstlj4U9OcjeT+vq4DNKd5IM77QUrHZyVZaCKmYBnT67KD1IKp5RhnnFEeL2FIJO9MbX
q69DVUakCLaHKaDYTj254r8p9d/BMkKjRZW3BD8FzSydMkWFVm9YleKgbZQMBTUWBRtoQwpdjuvs
1YrLTSdzC7LAIgYGzdk2jDfMRDs5u3U1Dd4JzQ5RmWbvQ5z3GC8oLfTNyqkEAGGAB1FEOASV3vc/
dcROZJeCzzy2O21Hh3zOKWYX763KOfTp/cTWP5lPTxzk90UfUTENx5kQ5ePq4nniENCPh0rhyHIL
GrfnIhEaBdl2AVPJaCAj5NAIy2oP262/4B44+5cofBBzc9U6qDZiWbA5XVG8Ylwj2Wvq6/oaady8
j7gyA7OFc3Zwn0qbuJxfwVRA+T3zNS0yDsk8w59j9FKpniL/s59/hHkH8AM7bU2IEaeb6eQF/FgB
7q9YDpy6RkYWa2sG4xlqCuz/6Vv7Nyv8IDNTRG5DY0+7sd6n82erj3qJo4r32JYjV+oGRUGSUBUW
w8zUPHed3IYOs8zPU4Ufj6L7cb5CwVa7y1fPUBKyKadzJPhRphD6iN9e4+Oflu0atFi+hyrECKzH
9R914aGlM5WXgAFkwTs4qwFWNRQ3wOUzjfYmD4kn/Tz/k8HgJzY6qUChFpdhCwR/2BZvqHtYnceV
2uOvJ9Ws0qNRqPI4xfmOqNnKmXq7SacPcym4jhUDqbiFIuCg4JKuZmf3as3YYhTIZasLu/a/AxXi
UdW7XKicR7v0JyTgyb8oGbajAvEuAz6gRu/Btsncdrn3utSS0ScmKvK6bVJN8rPrHpuDyGnPa+5S
P4FzuqSZDsr4fNEsmacjM+TUt7OY20v1OndrZR44mYNjhiCOPRmHXCwX6biajuJNP5FxTflrzI6k
KpHTPMGJqwMNNpReuDFWA6iiTGaUYPrdy92BWLIeZdDmZn99KQ/Vl/UfaM3wZBiy/UMn0bIc/+aL
oMhsa58/lBEB9yXXjIUCb/8yLzY7Y45tvi6fU7gcC6pCohLcnzkqOaOIXjcJ8PYyeyCEXZdGBJUv
/4nOpJzv/kITEnUw8G0ytSdSPQ9ctA4KOcrj+TTacAKa4rGxLRY+szORFTX9Oj/0dvhFYhAbXVi3
UNf9sHc0QrznHyRxWi/vPfuEmiEzZnlw1EVyQ/W8yKuXWQICgMD26wB2eTVuLiY1Lnrvlen9/5ae
oBy4iijX6qql27It0yD67uMmAuSkJkgLQGArJQSuNbPc17qVZgituUFkom6SDx+Wi7XXgmdxcHZz
Dk9jKjZLZV701SLk1E96G5HuP72EzX01sy9fEENj8B1JWv9/spAJgoviYi425m6vq0hpZN8DNie5
GUWCR3yS+acXzsf1o8hbZ9vheGqai4Y5oP1PwolTHVAjrgG1GREPCy2yzTYowSFIF8CJFrYO4A3V
5Du6xcku5+vrf+tHNqHTiahn5xMP0WljVGAeYIbUwawTTKXPbppnC64klmII2PtF9SJPccTjK3/b
0+SvOrS5sMTKeetqD8batapx0Nt0Wb5vsQHDV9U7Yq6Drev+xuM9kFSbWl/nOvJ+/X0FKAxBjg9v
s71ifdp5aNDzb7cJI6inBZVW+Vi7a9OCkMufX7whVDUCsCQ5xjBnvwnyWU5MfB9765C2/ZczOVaX
IH+SY8kBGoMN9mNfgcU+FF0rfrCZmXakC+jgBnDk8PxgSQ1aGPqxZ2mS817QoEKq2VRQKaCTmTjX
LXb4hxycwdYKpUElaxatttAgvlnMsMZJSpFD2o99S1lArntd7AxtOtwWSBah8wld56jfnE7cX7wI
MFpMyj/GyrItI3/9T6zEE8extijpHgLUTX7al8hniQmUK5Gk2bqt3I8eq7+0uPzgEfdQMjdH3zLZ
CVf71iGnqyqWA5J4aP8JjrQHMuaS24OAOChbodMl7VNdlgEmaapuO71OWwsnY2JEK7OpVijW3NhV
k11okI61Yz21yEzL3d5FPJU9UOp1+RVJzinsRPnGt4aLpqRwQ/+zvcvg1Sddplc34pIyP/DvserZ
vQfhFHs4P5PED9eIy0PJY57h/4g8Rx47zIfhrICYTlob/Xya9b9t9brid7n1XaTSkr51um1ifunw
j9QgUhPzZWd+eCCKYUJ68EJpEbjUeLGXtBll3pDAUNhES0ygy/xbfSvvp9BuEswgVH5prd2tctd2
45FzN7WIigdL8A60JQ1SgJycTxT99JYn9mmRLDfmS+kpfDsEmVeSiUo/e3FEMlQ2n4vzoHnCpzV6
CFwtu/7wSoegDsdF2K56mAeH0y/LUMSTYc77Vh8nsaFxW86UofIYluF7aODUGl/ZTXUFvz3HIHGb
TNo8Sz/BEo/YNzCpzKi8m7U1AqGi2HV/ktoVLk5/In9nwVErZ2/uc5BH8Xgjx4G8q0hxPik6FJQt
+TpgAdc7PuJFIgp4GiPdwYhdWPwxIApPxrqTC0TDmoRacJSGF4ZfowNdGOE0fdnjFgVkv7RmYmw/
Cfffkl/+aNv07Sz97zN3JhT/sm1If6kQ6ooVCJiokCxm4CUsoikbgw22N0ruvUNWlxJkXM8Vmf0J
l8zyLPwOMwRuOwmdWypi7/PTSNUW8tCstCcI9kHzyyP0Iv/YT6uZ4HFcOvsTVQoE5CGakGyUIHN8
zK08Dmzd0tGKNzu1oC12XtW19jlA+VYYhGNKD8+T+VXajorNmxWS2RBUBu7yZRc6juXBcYoeZQ82
DlZIgAITYailuD9eXa3r4qtvulX/3J7uCLBwlRxxuBJecZwgKjtyGnMFqnGwstqxkajtdfJBJfk3
1nUYZdotB2sum10K155PFYsaeTqmiUIaB1L2KFABBto2l/lDaWhqz2bBH+Qv4HEwL7VqbYn25TRN
/ejsX1oAhGkWh6J0YjYp9cgIGl+S0SAW8Cah2TLYVZowkvADzjHjTrw8PX5RjmLNnhwOdKIRexlJ
GBkNbAtB3smIlEH6ERPFZQakEerFvNu/QhfuSXyHRoz6xN9KXAoyfUI8RvXSNFRGPB6Ik4eyRrke
00X+DWrO2aMe9SKO44afNxKJq3orR/TtCug5PpxoNRgl2S+E4Daf1TjyESuMEBRtvvX1GD/DiS2r
hYXcQA37w3LDoFLm/wxMkLIJfPp/xXKj+rkRJrQFS5qrGtBweegJjhlTxx12QfC8Ar0alk9mg+0p
E8pgOonnL2+zs9cA4VKtzPO3K0bDi9ioQn3ltyeTDn0pxI1KzN2MUuPKi4Fjxt+LWl0dNTztfqsL
y5W3TucO18I3PLOLBTxzCnBXS6iVmtpQG1tfF+EU6i32B/u46JehbWuKFTpkz8kRaTFDB5ytH+uj
lsC07VafAGrFKdpkrPCdVEqXEKgA03tgRcsQ5ARg95Q9ZpE+1IgVbvfUmP8HrRgQYKgGZNSdr5x3
X80fOlfuXDFLJCAFEsF4LcqbPPzzRKby0pxZMeS0eM0AzTla2mJkJPc/EDOkNVLUhVzO0cs/cmC1
4mL+hFYSUqOvRAU7MEZntXyYWVakG5/p3j6+/AUKTK5K+xrJNOZyhouhRcxm2Z4rnuGlnzTWTmYI
zqp4anjLd94FMtU5YuHviFYZzv8tPsQlmWqtI/7Y6kpAE3x7jEdiq/F0hoJIPHLnrsdWFW2k3PJu
toQKcjgw5WNGMFgLDwitA7nLF+MO0a3l2lCa7MVWaIFaUDbaWkiiTZcLc1O4sDXZj5xXjf8TYgOl
6dJHi4eQpVADbJTRiQkZ3H2hGclqWvcPCSHVJxelef8mZosXXUFyGIqeeq/kQ2LNP6MDAMuxoQ7A
GoYAsAfNHwnuVqmH3Iw11aHa08U3hAb4SRDqgOg3fnXLPTL6i3K49CJJpSLC7dASO+0Vme+0Rt5d
2D9dNfuHb5g7d4MAWdGOOOMz7Jmpu0i4uUVay+nWJCXREGFgz5RAVB/Vnn3YIWt0BUIXoWHvzWVT
tA2blBYUiJKfl5RGdL9dcH9BKzQpejBDkKbC18adxAEECLxCiLVYERtodBbtT3l34mxWiKl2gj40
dESqz/1ZPjG2qbcyaphoUjv09VxiZqjOlh4+Ve8ApE12dScSv1X/zZ70BZ66ZEhjJzImrhUkZeZc
yGk6LWBPjMZoNlIusvahF8qm75GtE9vCzYvJ4tbi/CobZfjPUQXoOhNYaiw9aSzx+gl4CbR2jMRq
B9KAaAJC80Ol2xdDfoCeRY4wyTK4oEF1NBfovmA042YSuAK3Wd0dRmMXv9l6EL6YCorIUH0S8dg0
dW2rBI6vR7h9vfytvX2wAiDNQo3AOfAWfd+NR90jlhnPbnggDkph8RUk50uW2q0ULclIa7LOu3c/
+2X9FWp/L2t38sskBcx+xlyCiuBsn0ZEuwmFr9tkmQshcMimvPRRlTdXCKVIz1t7cLI1QCoHW2cf
vs9UBf/eEwYjr9JzaaTlcbvj6Z3pDDxIQ0R956BwlUeHo2JiQvvkAudFLXSomrHAYqaFXGiCCJyL
7rqwhpetJEK8RYN2JlxcEgy0l07xVMa5HGEQuT9vAz/FTY0PYDq4NXoRwdi3Hw01tvx0bTHsLcFE
b+2iawFDPijmw0lfgR+ISUINpou2qDqZmrBXzc2DZ5SsTWAvtYfTw75copc6n0NvnEuj2FiE2Fot
nhqzn2WOLufswFVlIyA+y+/nIGYcEXNWNaKlSqbZRGkRm2CsYRApB1M+r1ewNrrwfJCYCQch9eAz
C6/1yQWd52A9qoCMePd6FFrmbq8+KJaYce525tuYXWIAWHQfUmgvoqMPUnc1ccYbJGY0E6doGDVg
y2hPYFz6Tmg058YpmdJ3+fyAR2uLdytwuGNsIuUimiwyOp7kUaKp7XnXrLg2kC8DT19TcJ1vcpE0
DDNexAXHsju85lHOgyE88slwREoGMbAYqqHvxgKzCCp2JC+0lP2Wn27eHKrdgstvjb7OwrSVuObf
pUUdonVCop9YMGz0uWRdc4QYzrKRtPYNb3n3ejTr9uqjTT3Y+Dsx8JVPYdJO1wz/bTaG+izazPGp
N0WvlgoZyU7c8CEwf5obAps89zpKXA7pdLyi8+zhJTH1WZV4wC8sHgAlT5N/4vL9nawzcjEJUsIa
+aaZxrfyqrPfeLJXUYR4tmaYxP18+zik76hysmmP9GGXusAyOOgsyqki/3OdoiGShub705K3EB+4
CFCg0qwRJWVRhqLCOLboSDce0T1fWrBsIKS1aNDl4/rAkgxaqCvESJBlEHw+A2thvORwWtHj05lZ
4E6UEavEL3Fd9o4MMaDoNt98x/WqZ/03CMghjq6WUsbK01rnIgX7GixiZ9B6CoYbQKcnjEyHSGu4
h3+IC0f2KuUhqD2rRQNXimNGz8LFzJpwNbm4Ubqb6D5fUo4/b7p8U/kTOlepnyMpOuxwfKE8LPc0
TmN74XAA4cTCZprQWNDCx1x4R+38qa+3LgJDCwHgnUC/GxMPYDNRNLOP/MpWtbQie16T3R8Omoc+
V/J7Nw6LD3Th5cds4sQToClyz4dS06AO8m3I4DJOhlclUFaq0OSN2zHoSHjmC95XX+o+VMS4Bb87
zDT4dvYYgPX3QYmWP+v3bqiYgCzgmrBv1KOz0XmuSre++fWAmGU4bXIIbbBL8CH4sb1ggsrILxc+
nUbIhDuNLUu10duWtxEg4QKXraj2bo3ZWcuwyaZW6dIm09QpeZEbuHHXfLjLHwL6a9B6pcF6itm7
KpgrrzaXB0KTqrgPqV3BxqlaxytXdtt6KmrtGDFCtHlIUUm6HtF4y7OUfVUOiKje+vWQ/VH2Ybw1
WBxAvy8CZzsS++m36K0JyC+xqU5Be6CvMITe3FrvepFgmsApnCOa0rLEfxKEksdD8txYzY+j7s/8
1N4O9W0rm1elSEdI8nZDMiwME7AuimWSg4Uf67qu7g4NCdfVUjmDtHG+CZDdoLRbKsTeM4b13CCe
sfmhU0WwCadqX8d0O0X1z1lhuqHagvB6Y2E4KuAntjE//gWDVMn0VJBWquwrM7bFTLrtCkgii/rr
LaDYARZbNqHcsLYUMwbWsb1dZ3MeHUX7U/TMYoIgScuJp+UtCzfGwMqXWaP7Hd/fB205a5spB3Mh
Y3tGn4nt1V+M0aTc2EuweaoyjuJtI8r6dJ3Rl8huF9tBv4CTVGpOIGvqIBG1l0VVNZSQoPWwQShQ
SbbneKFE7a5sLd0WppYmpUsMDDV/T5vOtkBfpfyIe1UmIpcURXvWXnx9fZSg2WdUYGHeEWpe8n8X
mfYLKm9SaHMORymU80tmFZ3gC4Rx4iX7dC9BqXu5xyOWIB5nFR5suFV9QwJN6NPMU6s9fGl/V4sg
Xautsy1vGHCdK8bDWxcNTfWFUnXd/OUHytzUxFgWsWFEkYMK3gqU0QgwgBSK2kd4w37EcJSJ2KkB
9EV/4SzZzHUed+a7YeyigY+6ZPDlb94fmeBi1saTQ1PscS/GjxYolrUnoxsPHTGBdnIRHgCE8oL7
f+QxhVpfJ8JzI7jZnPsWAUjPxEX622IOc8IufOgoGunLrEPrSDOVn1HrDCuNHe+CAebrIKREX2hm
Jay3tGU0KyUHiDA/i9tAn+dKWiZ7ItDxIiImE8ttsMZSb0s9YjdXVOwfHyqeQIy9Qc8Nrf6TMQDA
1w8BPlq/HRNdrc8e23E9p/rLlcn+09hLol4/O015MyosS4zSXpXIGn3aXtGOeSn2s1Y00kgCwuRQ
yOGqURJIR7xO408RytdvQ/ZV5YvYDM2PlHTlkDvOxiM27qN9AhN2Fb4nwIqqZVdvlFJgPqD9PP+A
ggeWlpjQBKm2qjdAA5i8cp7xWwyWtOpXuMxEGKpyK7YR8aYy1NBlJ6h40D4i5odYbUP2VgNZuyWX
QRjGUfY2NVfKn+9L9EBtiGc/VtgvkVL3WS8CwdfiysyHMOhDbmsyviNNX49t4/IAZxMdiyXLOUXF
sk62rkhjt/YfTVGE7xGSEd3hgQUxikDoKx/473pzrqLFy0KNcBYHEVXLF0/wZbSjk+XqFabYfvBC
rEbah+bIAyl3KTeeX2jVsA2Img6atX+JlDfKYIzLyeHjhYmV2WSFREw2uhYGDYUOBZOluKVWFtZx
eE1ERKirFCSMlHcGmzGA93MKtjF56KnCHrMKq4UpBnO7bIiGKLzUiiNzU+ra+wasrZXUxcghVfzJ
AAhRkTRwoTaZ5q4CunqxvQ5IfS9hrpFaqe842aUR/CWkC91fzNkSE5agboN9irPexXhON20645KJ
per5DqJt5EwPMpugWzh+mTEXgpN4Dg4dOu9HA4ljlmON089t9IijP77aetx5Mq9mHYnnbuxdY9OX
Pcbt9DjyVBnq01FnXLGpcuesQpxTQb/b+4UMLq9o7GT7SLPtTsdl7/TV/KgcrLr7qWyPswKRBr8a
G3Urdc/F26x5jPFGTqU4xivMIrwHIKpfwiHXiNBIA+KV0CsAq9MGu2gCRcw7BqeSTS0hRKCgBgLG
PDVfF9yEcedM9oWr76ftR67bNReFbeJb9SaLdcMq+NwTUFdFMzk46j0HXDCAM91Dv6O3cCPxX5G3
/aeO0QKBAclb+ie7eRNzXEMvjCeX02JzK3MCck0P6f/0sDqcynbIP8LaH8DAjqvyl7pvlXmu2oo/
HWt7VmPH2dptDLGJz6ub8MyCcFkkP3QKeevCdhA+BRWyRu2Mx/2BgQnjvH5TYHBd6ZI8NPLuyJuq
F3n9bv8sEKlU652HGOqHEy5xQ1dZMOYLg/Db9ZBfA+kgCtGk+ozQPAHjs1Gmi1Z95asgzrOqMoGW
/YSS4OK0AIdWaBBHsTc5H4StZhzrVnxHK7sHQvSdIM5reXQkIyxgaz0dxrUFcYF1GFVGRd75q5yy
g0jhg7r/kAyzDDU8RzfRcaVIpOSmhG5u+uJFNfmrRlkcO1lwpgTLJyLzsGcXI2+rsVsuSW4uq/3j
IRxX1aKEK18lXMCto7Cm7Vl8k9/33ttoynTJiwED/wZFXP//vb1GHH5lWjA62xV2fcQw2pQ9ABCE
Q2mrx+0zS/F2eUCpZLYtQ4HpialGYfuIksan5kT2gUYpg1kifbIsFl6CBs1eYBNc9ADg6Ug98N4E
1azQ3f8RK6cTBSjsycUX46Ri1X7r3c9zJ5FZComY8liUZZb0LXhz+rp1dDgkfzqrVI4+MQu8JLhu
IfAaPkRM7igFOrL5tlVrScFs8iwSL76NpqAP2Tt4amd83CqJUeRsf5VmAMpv8RMdt2ZSPjX+UPu8
IOm2E0UXa+DVKGHG385YBCtYPMV+q3L/osB/hqUARuIX+g+/n0IkqAziAbZpTbwL5ZZix5mbSvhY
erxc2wLnLSn3JzGAnKqkOo4HzFibBP5RDL7guRNlNBk/e5Qwe04Wymd/RS10Vpn+I843qjLQLjbx
GV1X8dy5iC8XfhPIz7pgUsN0UyD9eVEpO2jUrh+sEpppf5q5w0q978P4RsI7/ot8Px8yqQ6/Y+Iy
J8U7XKKBvK2eJsTvdSNXRryLdcg8KYEG+lnvsNxVNKzkxK+omOoT1Trea+w1l68DQCZ+vN+FJHC3
9NnG1ySpQyb84VjHKXV2JpJfWwmjU/8KA17yAA+E8JpN91XBM2m1koD5NCqNLLbkLBHC5jvUFnu0
QRMlT7TpBj6qDs+8m+y8xeHNW2Hcs/k1o6Mq3zrMcvmd71PIzZO0V3tXJ3VVL9NK8fc0DQlXDsGn
JByM4GkFsLAKfPwYUpAP8rdUV7eHb/ckToFMGf426n7EBPzmcIDWz82B46w6bjCpDJieeEOG9t9V
D/mTK2RXi7jZi8jY1nGI+7Np0oe0Nxs/zmDprY8ryFK4/SoGQpbzCWG603Ixrh2H83Q+2fgYQxaj
GIGEK45/E9dY0GbOn8NwxZM5abrlnVNDZEhc3jFcVbx+mhBjXsuGt9POgzINJk4g15UFE+4NEAFV
GprDUEmwLrWGifsI/ezYdH+f449H8ylXgNqVm6+VUZRsOeOCaKW6wZbp3kS7OhIzVx/TgPeG02I+
Y2mNkW84/veFP/SVG1B6NtDaj3JDGf5LQNCCjvBkqf6O4gr47/qpMtQoSc5L5kFg/RaEvao3UMmR
QFv4gOD/3eGwipawUyQ+acZ/A5+Ws2TwjIO/1tFmzTx8qbXd6C7TUe+XWveGp7+toG0g3matPcu9
cQ/F5YejXowynSlR1W8QFJWFTRzbj/sm+LX3vlkklG0QmcpcTs3GmtLwF8feHbNHFIvVtZDjwRTH
65BMCYXmoEnXXf6jxc0yCcJyhMiJR12OkN/0318dM34gDLrcCUX0khctfYDApgezAoOpPHsQEM93
omQxNTy+tzDoWmzHVaOn0VP7I2blpvEVcFUjYTAGswK6IUXy0y5n9zX4CJxcz4PoZTf/ezadMNjW
4xjdVy5gNfln5yRqsNR6e1AkVg5Wq3Yw7YlsaXUlHEFoJxOlCu5EAY3G2RQOUakXoLCGO8YluQ9D
HFiw/ZxdOMe86AZFUH+0DBC6vzu/A2SWj7b0rCGD7737z81Op7p9mN5z3uHdnHDajz3VX2znS6RG
RS4HlSR+1xwL9assPOSkr3qvOnixS4w1jWaZzthk6EoaRV7ZHVjHwF55391RUjs3e7DgSptXp7lu
iFiXvKrBkJjaqduZUf5TMKBagjW8IfAOFHd7VEVofMMaofOA3SI6mfLwfrzh6W2R6H+VCIzQnBFk
ZBBQr5S6X+sQm3Y09Z9cVWqIOKsv0T16cRTEILOPcrIHnV0xv0ih4s3Dq+7RJlFZTezlZ/4fd0fx
lBgdcc8BXwC44hCvzDJPNmumu/Rs5wuRmIHZzmqIVYyffP4ndISGbT9FpYiget/CjvJzM6lYLpo7
IAx8IvaPdREcipK/V2fuOkQxI4ly98LR3bKmZlatcPLjmBP6MjvrN2mqk4R0rCtm5bC6sMOmtGZK
UfyKeewdn/ep3tatmeMC/VgwEevX7HSIzPWfVlJsnhvcui7/6YPybfkY4meSsn//TPQxxM5TQtU9
NGPlz2Hok+6gI0gvQRWOoRuNXSOlsmWA1htOiX69j/Euj9pDSiEzSHzEZVhMZPEpA9joEjEJGwJ+
vVWDESbjvZLfVJc7pN69tBr1hCygAeOr93nkSXZaJC50YCXOU7OTgiQIT6R8TqMr6SDDRReHsnsd
mYvq5uk59Ux2dZXoSm1lkgTH0cAl2bUNwX6cF3kwKZw90/iuu2MGk+uI8x9gZQ7JsHsUKjb2TNZu
keAyyxtxwqkuRNh2adrQdtJ2/sgvfZ57gkMR3vT7dBHhDNRlsWBc4NJlTQMIOjfivzLC9H1EQFMd
j/tdG3FKnbkLwxildXiwaZd8HQPv1LAgM4WkCGb0h6CuaOpRmmH45EcpN4cGbB+3HUr+b7hWeQgB
Tap1JBhbpa5LU4RoGiuybzZFzMkoCiFVogQv02rSYndB5OhGaRHLQi6VGVh36bfj7dpQk6IkTb4P
KEB3qabbzIFSgdskl4A0VvhSSQTpZrEn1zeMpi4R4tZq1ev3upkOsNCnR+K6wUrz4dtLfhry2B5C
8SHl2mb5S3nD1FCL6hgMQRxhGEGJS/7N0FqF7A/aBLkSobKPqKAHsgT8QH+FnX5bKIIh1FrKOPQq
8uUYM0dlAP28/I4QpA+AvzuMgenu5CWd8VdCbXGOrYNS5w9auBNY5DgFqBMVblKQL/k670oEsDwG
QOEiK5bSBX7I12NXALARKNwUD/hlvhlgA6g+kKeewIRBomi+w6Z1BUVbQktjdPi20oTW1gEvvxls
3ueTtl239B2i1vnzKeaJrZvZaUBIL5sm4eAFcNFhOdtIKn2eBHB68HKPAxEYRsx0Zql/+JgfPNRu
99rk+nOHyxHSOAlDFDP2CWqhUO/VoP4I9MUyfJQlExxBSjtl5SyrgOVk38ghIIZ0WFgUb3Hn0s1m
8Z3s+nDmW6fe2j9FJx5FBmEkmC6wme/RsVhwyU8Yvygz/5FQabv9hWj9qcQzLItEYVOUQ7v1PnzR
7wmx8OvzcQ0atf2aAIfFzXsFF4owHvBPTbigbNFBDr9+eExHQNIY+cDGwi9xsygSD5xj8YK8ETG3
Ne9ZqFw8sqL8yjAN/krcU9hNq9oZ1ZLkn1aOD432WuZdxR1jFpwel5apxYhymJEnLkg96foLYdzh
QVVOCuAl9358tOg++c3l74p4VCUS900h5A20DCDS4IXLHorwObRkbhH/QiWe1d69TiGGh3gOLRF6
7OF1rJtOCbeUnjj5cf0oJWfJ9O1NTTGuN/54hE8uNhoPr3HYRk2HzeyutZ475MdW4ICe6T7Y14/q
pm3G1SYiWCd54YhvNbIW3BeGa6+0Tkw3W9ZNiGvKkGoVTruKp67Wj4U2FgYqSCHSSyU9Hn+iP2pe
BRCyQUIJfp8Kk5htbvlxOWBhSbZdvI8YiV42TAq/uhKTI+ympZOHAWPMRgRFTq7mWcj6vVkozWY0
PTAjAoZxbrMCYA9n+No+IIPsEM7sKH91sSP/dKP1l0TYjuk2TncPdKJlWjeoOrZoMczfg7ybleC6
rQ5RGkcEQXmvhOpJat7zStV9EOJ07M7qhgLONZQoX7kV+kUbOtP2d4JauPmcEnA9l3GPbtZb/0Wz
uJy9IxTEwoxhMOfQcenX3APnVfEmhS3TQNB+AFnZpQN8dLrd8oECa9tJ8SegDGqFopjdJOA0WVzF
sVMw8RzS36ILvw8+9OgeRCF0zBnqrAHTc1Tqn+qeos3E4pVKIevaUBogytQ0o+R+opHF8DTwUj8+
4i07mIusuWEu5Wtj+jGSBYIYdpDu0EKCOagi5DvyEHG8xpcjRPJGlQobPczELy/78HHU+X0Yul43
gRSwqnVbr66bcIXm1tvmSZOjgm3WbD5mA3cES0ouRnSBB+JYWp/d8fDHDDXReO+Shn0X7YfJlCtj
1A7CcAmjWhojq3gwKx2bFSsAA4IidaCugwxwcALVe00koNXgRh8j9GdFH16f0Ad+C+A2NUklytJv
ZdfeU904YdF+X1xhx2i7dlohFKBpmB2EliZjebvHVYAyeFsMQmetV3x40jYAHJJE1s+d0vUpUB6l
uB0/OLyJCRbdD/WMBfw1Mcg6cbwZ5VRGfCn+rCl9FUhW6yFoLe/EZeZ76y+Zym0lK2cmPpBj0kap
PwQigpIz4A67klUhmZIClxYIj4x/BpzJfbTSg+uWzs54Od1DQGCw0TYGy1DwBk8s43jwo+MLR38D
lc0jp9YNGLRDZZyZjxOWTj2OS42tJrHBkVOn1PvQMGMJCh6cIVEgeN4Zq6agPdFA452pGZgos8Mn
Sz1slO/BPkV6lzfmTf+Je1So/UixFACNGU+mD4mVrJ4Ctzi8/AlFQHD8B9TOdJzrirwjQMQOwMCi
uMhACLoIEqep8ZBj8iny1hdu2kPZUAXIbseWXoc493Zj6eCsVRWjPLiWGJ1KLkofv/5weHgjlFYa
0NsEjW+Tr7ZAmNXc5gj7W8kEXnuQagdMUoF4au21B3lxYw5l/tbbstq0U/2lLRP6nrVrX4JpwlHi
2SqwjzCqLYGtIuk6Xy3Xs2KCab6ue57lMuYkDBvVZUSR6Nnw+6r6DH7qOk2u3NBGsxtglNhv4hAj
m15lP6ul18MOwrhBjIE2tWEWl9FpVQ0zJlPLNfsbftvIqzg5e5jb75NWBMfW57JnCMuQTKWkfYyw
7fL+j7brD/W2JnMXSeV+uvnN8/+lRo+boptVsx5naQ1SfbIP00AJ+XcuHsQabZ88UklZZxRQ+Mh6
3lBxXc2huadCMlrdWIgXLWzRYmgN6bqYWVaXuv5yWGTB4+MGzOBLLAQPPqO4Adkxt+WqGCnzTuUy
32VI7n6wsViMJRmxRj+dD5smQpY6yfM5LYiXGrja96a5tJI5m8aFBa2jW5yoaNaVX75VwImmtlQ4
y1C2uz9aFN60CSHGXseB8885mPzfO+ja0nZ9zl0wZM7owK9+XCpYIisKHctqodlxESOCKBCr1IO/
ATV1GN9LreVgvBJssQ1ZLR4KWUrWrnZgtWosK1EH89UQwZHt12sELwiK2J3UQ55i8LWS3wqr+9VV
rzMvyM82Yjfq2F5ER24YFruqi7AHtUqTLMg68CwyKtgMMAxER5J21/LPkwnZbVUYR5bV5MXy0jhN
lCxcUC0F2t/jZQnjiA+vI8qsWxFrUeIoLN256uSKCh3hoNhlQmub25Y9t6MWUSZZXwlkm2KHeDFb
7fRDpxOPOc953xTYONy+Ox9a0LHbRKivIEbT2KoUCJbLJD4DGL+fczZkmkkxL9qIdV7HvsxhZYtV
WW0Cg7xQJAegxBi4LTiyveBS9ZU8uf7rrTdM8jLZdA8/5tRow0bjq2VQ6eLjrLOr7AyJHLU/v3dM
HtH+kHuIW0eG6VcXDy7ikSJx3yy8TlrTNNti733QI2wlYn7BYPtk8XgS4a702BQ/BLFQMmxmSckP
ID9+we1We9oB2+LnItVF3aKPYJos6tWbFbpqGxgUmCVd9Lx5Cml6MKoYr2gClh4tDOtRSsV3ip3S
dYE1fUT0TSqG+vtWPe0iFpq0k55yPM6DwF3Xy+1y00kbaU6wWqE0ZgXOhp0T3RRcF9xd/q0kzClf
A/usbdUWZW7zjoLW0nxMkGawYWZc/b35Obyy78s1h1L2fazz6q7/M5vgWPAeyysevc+6855UYbwC
npxHCD4Vknkhn+irp5EVuEUoDCRzegp1jqPQ61/6N7n+wTU9CygjXy7M0goxcJppa88gR0Mn1iJS
29TNRwLgiGI9OIaX301Ccg1/+P5g+V7peMA/vxjTNAGjPMDbdXSeu96mLNeFcMuRowvwo80TcRSM
juuTqhs+sFSdW5Os8nDfvnFA3bNpY04slvE5X7vtrXgsexp1ogUvb4qbjshQBn9WJhWMywp9gc06
zRGloEaXwqXTb+OUzRAmlw2xqSfShZwzT5yM3YPEgeiqYqx6J8nUGSnDfjQnp/aEFnYzvYG8f51X
VcwGgSHdlv92VgV/mK208jJ5ct7qge1DrTn1UQ28pMA+iaofoERKid2nhB8nwZO9OUkEUpUcG+g4
96fpp/56lsITMWGx+Sjt1P4LomeynPWhMMUltALE8suQ04ZBCZNTkES8iwVyQ/l/8raEc8dVPgqv
G21s1zluSonxX8QGe4HiNTeVKAz+of2JqLmAphgbxrxt8/CCKt4YPggzrwwhsMxFvL08INIDH4wR
Tj1f7rbkVwGHd8jt9hHdZF6wKRaLm4P8EE6EdYBY3NIVU4F43cpad/yjqeqWquvMSt7n2HE79qSp
qkXxenquc+WZesmOm77JwXybt7QRwEGfqzWKzq3ZiqRceTGg2u92PxaFIlDvT/aeXIku/bMbp9G2
3H3qt0LcvYHiXI1flXxNByXqEN7dirVJjOyafsvQ4HsSTO/uzYSLZG3OdfVBqmmJ0LXGHduTeotR
rp/+Zx+N4TdBvsfgxlpt+YFf7T1DnxhYVsvs0+nc2y1m8HOAFFio0yfvwVc5RhUC6djToKh24xL9
ScBasOtS/f7qQr7WJJNjxzTR/iVkzxFVhid6Vd0F9XrLm9cgP5LoIQBMjtumqPoOE5U6/pF7I5tS
Vp/2QvH3jrM0yDH5UPNXwLDlLeCkDlhiMB3TcLAd+03fNeFvm5QO9nscWaOXlshev7OuwuJ4yOcC
7Jq4tTq1wmD6nCGtJJnmJupaf2FT1myFFlgdiGGD/qcAzDhkG/9ZY1Voanuxr9EQTbR3XZTbvRjZ
f5RN+2kPgej5uhu4zQsOd1ziulacHG8j3NKlgRzfm0M3CYT3AyzjaSpqDsaGykcmcL/xAl92dnfD
Mx6sGrhJ1+Pw2UkoXhpfBAxmp4gW67W/h8mKSo8sJE/eYZpZ+E5fx2SKaJXRVa7ZnUOVrh7TteW6
ky926FsHkkB5SrPpWfkmUXxDDMgrM1vwvrm3WghWA9Ftr98sZSgr5TnQhFHPcDscz1VUETsLpXcD
JyFMUgj3taDkv0PfdAimKqQEfCJtIijGk5wFsqZM8XcZvEdEyFJ32sHmOjiv7e005oOJ24wG2gXt
pg4ZHuJd43T9jxPXG2L+AUsRZaJtpkjt8mO6URubUerCggVfufNdElczNA+2GvqFGjaZlw2O3ISP
+8PXlyf29DNex47nCzCcI1Gw/3lKrHFVYNq6jzRF2FXmC5HlbxbWhGHto5w5bwVP7xuB5AJcazZr
XeEqiRbEyvlgoPqXeStvX3zZQ5HRO3rMzn4YgmqlLgXITWWY7sciRHsKdYjxLcohu/5ViRmY1Sqz
8Wxl8zAflYBvjvYF8VU/cUe6DKbehThQDdpJ6ws3g7nY278oNJoPRA7zALsXTGf4Y5s30bFXWldy
+Qf/fmVjra+cw43A5qxk/PfUb3EqTyFCnb5SyMRVKuN+fbfiDNwl9j3Y+Qz/qD6aVOT7YRMB+/KU
5qFcWUsbZyPWBQRbLlL7t9HUEIamTUSLZPYIAX0jz9Z8ETeji9jvoXvcD6XCtlVvc9GhY0IRjc4n
SqrModjpaxzuY9d4ZKeyYqQ54Ik5Sby0CioyKLtQ4jIQZ/CWCXV3xNmKZ7nr/zS2kM/DjxBX/Lki
t9wPuEZlwafBKUlYwFIGvUlMi/7g1iN+ESIqwzwoDFLOPCvfRhiwElyP2rg8t4hjalxcia3KbTap
GFEsnYD448OfA4Tu1X8ew/+qpxvBq8zSRimyEaKP9TlfJfAj35LKY/ud6hh3iQxZn1hhcYH3EIAX
yHmcslJaGTQQIH5E9Jw+3UsVJNc7CEOtInwByvZbpuzBCw+OZdJh+zQajEX0paYIuILOhDMc6WqY
PMhs29kzggKBXEazpjExtuV4VD+oDMVt06KvmGCTc84OxDV8OPHhLt1bfgqS4hPUlLUJMsRebobe
esQ3/74L6gJRyqfdBYY+5/vuBqOSMkWWrVDcFovVums8NJjgjVIRS65MvQAm+q7GFcrEHSoP5I+7
12uH4vK9Ab7GyQ95EDP4Mu1gxXhWzP8ZxPvmgJ3UTFgmGMASA8wJKfGIrVk0vapqMZ2/iHEMaw7l
S53Hx1kFopC+tW2hPVJfWg4dBf8lkDik10E6iPve+H52jNi+hK0R9r+Lr4ur0qgQ1aDHRN/FyQmb
xNZwqSP8WmBptuy93lBYjqWOWohFxYUpb5vlYM3QZL1MRYkMivMiZITeXUDmVrUpRouBMMbzJ5Xk
1r/zougqfq6qEzWk2LB7UvBpidy0Qa2mzg9FYdEW1O+g3pDkt5niTgkoT/1WG5ijSFwagUuUOSLS
voWBcEQxl+HIhGNYoxDgYaFhJcg5WCglLri3pmLG/Erhh4EdIBkP7Ox1DtaxTSkekYuEl0cDWzRE
UEb/5WGF3pcF66b81EG3vkMzzbdxdVJghbac9fsM/DzueJ82byC8OUG080m/Uui3axuFrd3CT97q
R8/pZrMSKpyIJSIlb6DymcSj0VVg37g7YvjUsMHoqEhicmiO3bZITIZAh0kkvQ6ffxmbn6uo0Efh
qiSX+721CFtGKvTe30ty3BmNIiCpx81HT42Y5+fwUS9fStUdYQ6dXNWQ0bpMUysTJ3UOpWFxc5xw
hAYJ00ccH9+wOUtKB+PtCR8xn8BSvJFslg2RtVjIjCdHwF13N4DBKdn9X3866eEZUWQpcDmfKop+
HkYyZR7hq7HM2DmROhL4X7/huUsqUK8kOvPVEg1oPHgNWIGizgdPA8X26ZmciJAFQ9TmvKY0lmHs
HbwtH3aHCC+Q9I+aZ5kGEZvQT8IxfYNJQmCATjN4HYxz6EorynCc+F58ZBN5eDOGMpGASjEaPCur
PZZCFo44W7MqmQmDZujcYIFTZ84WNoyyxl5sKJI6ziXDTB9y4H1Z2C4bJ5TzxTFxM4YLFRq9f2iE
5FdbKokT5cf3BDIBfvIlO8o5dkHbKuUufnKyxgFDovlxXUaRiKVeWnHcxkf9IEhucCYM12Jq2fkc
u6ZXxfYze47BRi336hY5RMWp4yj26vgqhoppGo5DtUBeOiJACp+37jdLz4Ifad5eBCCdTvZDAPs9
t0osJMxBbgCgeLxIiA6P8ARr9oxoZS3pS5Tz2tRAC+qiZG5bs42EA9JBUL5oTlKwQCUt/uESzppW
qKhS8CtMRF2wHFaPIiOkgUWr0Qb7rUk3TWVyv3vlTORSsINRuskmpblAvZDdRMJWSlLM217nDdR5
Yoz8hCpE8XRuFSg7yBXFHPQaBC321Ucka+wYd7aeCBJ+nVFFPLz1Kd2cvL0MLm8wyuxcwBwM+FuC
SmsONvCC0O/WAf3c0nnNMWca6KrHq7TbkWFQIIUCFo1GygAenc824rVyiX2BKnoY8X73A6lNPE7n
bEaEk+XNsL2SqaCWlEPTtOnSRawAK0NTsApZPp5hP9kTwIgSojpBzvAY2uGzr8Vs0zuN+WCZ7t/O
AObV8CFewiuUfB866QAHkseiKf2+Wj2w7q+6S5P+o7FISTGjwJl0O4BhtCxDK+Uui+uVdUEmSVUZ
/wx9AQMRaVw37z3SdYUIWbWroP3tMB2/XiGts7Zn+rEypD1g7Sk2sDong8kmUcu+Wq+hXF7kJfPT
eODgO4oiUCnaXP3qlYvTZroSU4AmvclsN3DyE7jeN4FUlbHLwmQdAWKvo4sq4i6cTtwFB2/ezdJg
XjQ13xDliXuXvx6gfNpu1aqU8MTspKbd887akiqUMiC83P/fiPLdG4borzcEpZ7z7sGaTVjOR/wE
6V0WtdbVK8nb/APmp6qs+QaJYuZjHqJI2guUaZ32C+ipEWQQezbUy5uLyYtSwVhsGWkEgLRwo8rw
mBBbydY2RaX4XH8S7DwpKCr6QXPeZZDygp9Z64uMGK90cEvHAgMvgKU0lc2A1w4IZ2vqB8ibQfRO
Uob9YsmUtS1RAAGgtNrMBzvBBhVyW3EGtUJpVUP10HveX3HQ0d1BbtQ39jfhlcKRi9EyEQW7SIL6
Tuc39gR/6xyxaJnP/k4QGcOPTCgLKvF069TQILN3jBI7Ky3zBbUZPV2e9jW27K3Yw5wNuj7WAvY+
eskYRMbO5s+9VtGVHBWoXpegusgzX3v98mQTl6Km1V+dhbwjkehYzzrHdy9oMpU+YonyjeAg5Oen
OjZMS/ZZs7QqkvXb+wf2g6t3xz4FerwRWzbxKVTFaljD/62d+/iK5WquwnLlQnEpJ7P5LitVDNVP
wgYlB/y1GnsuSjjMKAiyn/+ZiwSUg/5uF6kCq3wXC5tRMk/mL1sXguLJf1x4EXjiGXtEd+yTrd38
BnpjL4L/pWxCpbwLtFGN/p2tTc60ClN9e6dyXrS5BMTzeCtBgO66JJB4vAqFVKHSVqVGwBsgH72J
Ba11224mbwbqEcvlWqg+2FCOKEUxqFVjkmhMQGDv16EUXzQ2bFHx+50stx5jolZaboH7jzE7cS/O
Kzn4WE27eMY28sp0hEUQLZckCCDfWwxEu/wr3m62XJ/3558asf0O65UHFc6jWOV4H/vt4S1eftA9
j4SZb5xbyDLs01CP2QGF9jklb4UbZohScC/02KeOHijUJKTc9EpyE+xAGzODqX3Pm1jR/rQzm6CC
rdg77dMwMLYvtxzRrEoFEiDTFpS0c0J2eyd6GstEpsRrBROPLt3vHBzk9rTF/M10HIUMwXfF10L5
3gB1s7cLgC9+H/MHbPxosaGfVKyoPaHK+kfD0mnatTb7xTxKb4YV08xeIcdKhM4QbjQT/rbtrqij
wzCjUp6u40IC5jaueKnDj58JjdOHQRuKb2KrkfXRqyDASwYwfvDsldGlMf5SiEgvoKSGjYvEqGHm
po9QcQA9weH/fSpaonDUVeBXnKddPptS97M2YNOGxYaqza/5SUQcFuw3FPFC3RRK/WYlXYGY4uT+
JGMedCbVWAanf6YTP6oeC0CfpGGiXzWvEjAims+J92QdeuLk71Fl6aJfiBweAspt4VJE+0nHUlls
7v8ARLOcX9OpcFHs6U4F9ooQIoY+IILxu+yRc6TWbO27ASPdNtAY0/Z2jorgT9NWcCz0uUnH29TU
24/LvOKxUlNfa0z8Up0rePugO6LQKkVItYokBRhnAJGUIF8UV1eVcpbywS98VUFH+VMXsXy3YTXV
HNb19aDhUjcDWmMxz9ZC7XO7tYWTYD3se33BsAUbUcKEjpRBjt7es4zOlIvzNf4Ivl+Os71e6P1r
8AGOCGdyJt9LHnPAljJbs29wLXJpg3jZ2z5bME1Uk/jJ3McrtTKPiQ6ex63BHlZ6z+L7XM4tGasl
LhpK2EmS/SD6V3OD1WhZWsXajDro0u5NMSWebH4JoqVSp/dNDdFNhyutG6Og6eMwIty8Mx9pxuPx
vE43WJ0fdKa6LPaRN5W8w27krxkJIVocwYkwFn7vdpyXOqmCUPfI4aN5hbPPrjK8yNmw7xLnzUtN
Qru4WkwE1+bTxsnLXqrEE8nLDaYzmdPMLFN2TidJJ0Ptj3dO9AN7WJAD62PD/AH7unJF4ZMkZlql
2f0/diuvZNcfFWmlXpMxYVn8hMnXz+OBpn3DJe3aSiWWzQCxec8V5q1V5ry8GDxRHkcDwXLbxsxc
G6hn7jffJAWoh4XJuMj9ok0dYlPlU+qMs4s/ZNzNM+MWSFUyPsjzkP9GWH3t6ReTVIoBQrnfdbNh
VMw/8wh7Uv/GQbeKepH9EVT0LEWs211BxXD/xkkGRfEJOeQCpY5LGjkD9J4cVVaU4V5+8nykM9g/
m26222feb3XPJtYw4lDJg7/SsfxuyrbxwdUP0xKtdmqF51Fjy6GTtRqpQ2TAH3GHJ/vV3uWJ+NMV
QyA25G7iMbThEAgu8l1XE8CS7mQ1Sr30gxi9fhsC6rf1D0Jw+S7OHfkPHcj2X3exIimYNHePFK/O
SH/nMNWyBewIxP4FLwLe8U+/VdMxsOCYV6gAOYkeAUoQZOJtvSHt5Ysl+AJrJt5tx/m4wvZ9Z5Y7
3XnffDmZOoLmlNViyZjzmCaA6P3NttLh0UdaEjzgzoaY8JLN8sMSQY1xfCm0AWZUOUI1F66cHD1O
jGWonZf1ccy7j3RY9HwXDf+dcQakp8pT3d5l/wincyxQLSihBBZoumBeV/mwfxpB7RQrEmT/COJ+
ANTGKg7vDIZwKCf3VH3MWUWIV4QXiGDWD98Jl4/oUGVmHAH6yZYvGrhNydvmhix/HeLJp75QgZAw
RQtyDuqU2mQKkxVd9QwM4YK/drdtqJvnpI6eT4cG1T/xhnSwkvRwLdOTbzpFqSQ26TNvijwvyGDw
as0MfCZYzpcyN1cv7ZZjTv6Ea9tfEFGyOm67T/VFaeejnx/PZ+32mYXjPN0q+a8QVwsBa5q2iDoy
J1QFoKyI7tdif/umHsbgBOhLoOKHRn+FZXRrqJruILYJnmFKKyl643VBW1K/MbzXs551kL2fCiwh
JcvmDx1fYSmlAo1AoAgLEQstjlFgazKPQxw2OAHQV6s2dSWUvosaSo80OLKPUMOMJ57GQ0ZjdKBj
f4PNXL+y3i7xISOHkg13ZZY9hxZDJLychK3NHOs3ekQnLVc4g30nO8nQjvGM2uk/BdxbpLYJPcuB
BRNxZ4FF9cON7Ujz1eLZzpRUcHlOMQPqrXu2x4kLzEAron7hG/fB1KkubCB8OQozjlqtd6dbmg55
lnJN0h1+svFy72vlQqyA9om/bMILsTixLFaZsWRboVL6xJygA+HvcOpdnZJ1FggLOVocNaCS1Duv
eOR1eeHOCQBCxeWnxZ9rVk5EL/y8QMfUg0sOTGkPD83mRy90x3yqh71+l86AvBXgmea3jqsV9trv
ny0yI8WhLie0Q9wtGNfkwR4U9/nHvobOAeX5TO3CISPy9qKX9ojx5hpV0XkXJ+dg/bONnhmvNQSH
Ec54LiOvgMPV++oyHjEAkkKs0x921eR6tc5iX0NE3DkX/2VPVMHoxJTm+dW2ho6uTHS/T1MI5cMk
XjDnmiC15QFOyZeJ1q0NrmcwRRDLekYxFpmb12I+0bkIAo40yn0pI9l8nCBVfeBHY289SrBKfWt+
+8FyC6IpV+jMKPqDzOEGtvjhwe7vPVctRhB/YKAcjnZx88Nkz0diNSiwidpt1AuUqCYNAU9OY1nE
xiteuO8Lqj/avCA5GiuZkeeZtISC1esdFj7TwsGurwL2RZ37RM4cZvUtE4W9fLYtGwmH5hOSebWP
itnI71dOMgOphPovY/hE7XFigqLnNwDvIjCW6aULxEg8+j+O10cpZz53elu7TZrSk63KVSm8bAP+
duge2QBUCDafMLT46WpJgtd9ujn/3W17uelyW8n835z2NhpH/n08PR96t5MPDfwXiIYh1ZlWWehk
azizMxEa6tPdHDVPJn7F1sFP/ew+Hgfa2WpWd4W52uuBAUpgQdvZyOb4zbfixYYz8xLaqJA1KcnH
GBgvkBHyRBNQz5evPhIDHhBBZB/SXLJ+FnIW2kAgniACSN++Lvdm6s+lSKx2lNqBeMaCCi5HRZYE
3BleEbWlUOQUbvO5kHrDzH0Fqph9XoPgAVgMxPX9XblY0rI2kkKGmRK/NEuJo7yGItMVUo+RUL6j
G1RJNridlu9PGZ0dzZefvAXR5RpuzlZD9WcNWYdcPhKDn0XwjJZMhMV55HfGDrkuW/RjMEu9+WBy
8KpVDVOrVbj+PmxRwAafgFHZCCA1PLCDpv2jeZY1doZB4181zLWB4/NCAfDgJak0fxfG469d7YA4
DUmNephEn+exHzAd4TkuWrYMs6WUDGjt00TqOlJXqJeI9VMAgfo1s+I6dUyis0q79xGBnQU5y38i
QlCg2bvx/Nx0RdBvrlt6E4LW6Wq9B81z7yM7wRxDFYtvJsz3EQyi/Le9iXRdu9AmfjLPfpobygQC
ZvoTfLJYDmrOw4/K0uE/AoUnQMAWeWKIRQAYo6RWYcvpJ5dAh+oyCCvrUPfDYHoxM3InI0nAz25g
w6cs3UYsNrbyh+BRDC+oi1lwER7n4XsG1kmVggf5k3cVv98A+tlfJKHmeRxM/o7Ss1UYQyrKFavo
iMm6TyYpCbg7MUuSLg+nPoiNOSEjwtcra+Up7dwPELQ/v5SLiYiSd4mgpDusXzgWzbYE74dUeUw3
ydy6fwWP5uxNCFVVYNHySomUtYM5mAByP02lYKLtTnIXFJ6oNDUkUqvqr4l95ccBziQJQEpPQFE9
j6kLK84EqdxAeNfdeaa51T175biUCwRzguJwQX+Gmo3yRR/W/FfovXC6t8iG0KbHIZKhoeTshop9
9CaSe3j6NIDSLmLxQQMtGY60a3VsJ3rFgdXqxMN2LSP+GvFcXBIKBVcjOln/+CPKzGWofCMQHpv3
23SFj++FFb46c0oMJU1SAIi7HTjZG+3Y+rpLOVk1eCGkM+mTwlYuzn2wenPUHK8qK+RCXCXQs5Kj
7ZhJLfobWrIGqiXKjlcXPK8AVOpbQVQV1fY7xLl9BQlA20rjHcPzopUlKV5uIQHruah8zQyIbY3n
/5+KrFb5OssdZs6HSjcBNqdWvXzH8wHoAAhj9cWAGseV7y7us9XS7uGNiHZZFV1lYavnec1piMfk
Aa6XJAKzM3YZWQ+6yCiuOgQln+a/nfOavSLcAlTdd9TmCY8vZinmRZL/3T5DU387BPlD5RzDu5sJ
fc/c5xeuYUqAi35d50tn03Ce4gxzkN8dgcVs6tML61Lg5lsEmj+W1RcffN3JJsR8rqDGGEA47bGh
LUuYYrR1DlJOW+kGtWRGwIoYgr0He6iUpCiko+DJt87VJiDhbFoOJmP3cmSJl7C9H2wQlum7sImj
JmVUEi9Fu903HKTKA0FE+qmWgIjS3munGfpX8MDPuByPBvMmvg93uIuYu/uxgiOrcgGlMwG0505e
Nt4VRTUsJwdPC1dcJP/c7ieQzRzX7Th0QIv0XE1I0iSquE/mhYrPlm6BBZFLDEmsIADc7EHV+CNZ
9/gLG2Re3P1zmnEMqZadauyKx2BnRs2U3dVoPMxlxX9UIu3cDsqBrR29zLVsp3+mlsi4L797FO41
u9EhFG/U7Po2Gd31SPr8k+TQAPUE0J8P2rvhoqQ1Zid+62pZXvbnJN0idJKotMdLQRK06995i/QR
htzcL1ouRHu7jQNwF8ET2gWivZ2aZOFTaNWTUkCXEPVpPRzoXFG+Ahjotd2VI7x3na2ECKSP07m0
+hKwqsU4zbiHv01TG9nmeLdtK+OwH5AwjGrU9vO90doDH3Ngsdqz1dYNSHQNwItCh7+0LXT0TAYE
+O8al0q5qqQbHzNt4K7zyG0REjEheAIj4yRliHODoxxN5lw42Fg+L7aRv+M5a4Z/AzafzP78CL5U
uQ6o6K+s1iYuVzI7s5KVJh8zdimfZrkQpctqUwOqmQTC0VFWp7I2Hu+XxK9Hfk7mpiDZ+GM1EQNS
mtIeB4EZEGqvZbizLI3dusaAngp8bH8OyjTcMKCa6ejvS4vpSc8CbxNmHsW5CQOdUtaDkOSAwXWU
ANKrYYstbi7FqcKZGW9inHnbCZbmvOirsj+EPu6BXTmsTeLMPhALIiRsIK+G9ml4kkViQFvQ9RpY
MaTpb6tBtyAgznFuueKuBlxvTol5rykqv6j0icu1M462TLe9aAJID11k5+rB1LlrNVKCspZphlgv
tDVxNSVJ4HjqAHAnxb0+Lim3tNc4Zd9kmNLb971qoae0d2BDKW34LxgTn+uwhTah8otZcb8qkvQ9
qj9lhiGCwalhflXcwYZsfwHlf3+3TtGNq1hsJhaThu2rDZLd3cjZskck1H+gCfJQV8C1O4ueuBvV
kmE5e0NiECvBOatzge5OZjkG9u/v7qGITpSE5axo/FK12Jxhb8fUOkHsFnkVGMz/mVJArMwiEcDa
TpJJ/UpYtMua2uJyRee8K4maI+PFqNIHC92xXwDGI+NlPdFUU8jxzVnKZDDTaA8Rrkn4vuyxIv3q
n92BW+KpPHnccMKvnwsahHSdly17kfw/G1Xhqh46E3FotORq9+It7IsXBCpemqnWggaVEFar/KlP
Dd1G6vterUnSgyWHqnxsAEXL2yS+z6hFrmLo2CR7VzfJ8BwJr+K47sLuz9PbPE8KVVzVEDSyUfaJ
Lp5Mg6LEHKkOeSGg0CH7MsxFsqjWkfEKPKips7S2O8d91FzCuZnHnGEh5ZPFxIdDdMIj4j4RZJIc
cIf8NNMpMf77Fz8srUM4y8hfeQ79vMH79/S9yaTddiLmigZCJLOGRxJnfnt0ZSEE4OSThyIPouOg
hNJjpuAYTcR+ieJuKwQH96L9UreUm/y6dAq+8YUvT7TxBor1XI4OHibHSsTX64tenTkpWZIXApb0
Vdm43h1lL6jknZa14Mj/rD2xM30RI9feF4K1/YG8S1+34dLZ/CSFR5akBJMOYDm9RWkPKiTjqOvN
e4cAWHa6uA/qTWERwpV3SZrJwMya2ziSEsjtfj++lMGwpJIMv1opj8d+NNZ+PbqvbdyrXw/u5LgP
/7GmUDbpMVEEWZnabK+wSFwLIJd1ViOgRdV4+dJK265yKL2hcVM0GO2vzMaBigKTViSnOeKorUtF
/5FqDHu7MLAqWt8UjLteXtpN7UTV8E+U+Vf57271612FsDquHo/5sA8AGedxTDC4b7lFAIv7JFtF
2+NOIeESyOHBKWb97BVykv6IAjmAahiEk2QDtSD0HK1N/kSKro5Pwz5YmleKFyng9UNkmfvHWnV/
P8gde4Tv2jr0zyMjpwGld/w/pcERZ3enwK2hagXTrr9m1pt5DABaaE4up1QVKQh31f8LvbWfQIkn
0QVYgnfGU486ln9P8v/U7e5iOo+R30+k2uAddzEAAf5F3FIe7WpV8pk/SMBjBfTFzwSW7Y2UpUcd
inpO4c/NmdYYnkjQ352xmukxtCvUqOLOML1Y/B0We+2EfTmhaF10w+5as9c3048yvUmC+0inz9eM
4ct9ATCKriCnfuzL4b0ZYqdVwoLPRdcPsjXVhtl6IinNykcQJ83MAXFbIdi4HBm99EClguC+mpTP
/rJBQNVvZrkG/nQr55J1KHuIgDWrkqQJ2LxT7QZtcOo12nkmmOB5OQ0FCdalR4dzgFpf2snHwRLP
ppXMK+PvoVL6LFnIJQDkhl76dSq95WLvcQ5iDniS+Bg8gXXLx6vSV/sg1sWeg//UL1m2sxKaS0+d
OFs7uCKOXAje9jLrjqKSfKf5c1qRCKLpj6peNGBX0gsm555hw59TRo4lyB3wgXK2Cwab5wpSVni3
7ox9UMHXEQw7unGTvimURu2uGGqCTeqhkFRH8lbRZdLoyitj7MIl0OYWH5CrAISe55jhFQoS4JZh
cnD3rE+xtORlVRSEwAcRn2MHYt/nVQEkfkzL/xUc3D3PKvVK1Fk7fekixO5gvc6uOWKT66dzDgF3
uqrtqOnMY05119bhxWDI7SrPhE3RFrEw6a5eYnk7bOc/dJp8W8JKN7nlep7gfbl1/YUjzKdlOGAo
HTdo6rXp3csr7/1Z/C3XpI3hAG5FQ08bn+7Y6+Z+Yu/qzarxIUD+t8qnk5v8ryPriVcXgnHk5x6d
cZSN2PwCzLS1AvBM6hJnEHibXHFoCM5iZ8YEcRfLTarDNWAbdiGhogUnLCWP43DZTO/cjhLhh+Dh
AWw0HLJ3F5+GBl0rgEwE/P6GXjxUslziuPZRm1F1bTZBJB9j9WRqZu8QZbLjeTVlbqvGh/ZzCIN1
HccGFrySaeRjZQzJSnQOGcTjZe6qqaUj13pQpt4V4XcbjoNmsqtB60186m2e62F6WXQ+INY9PyWz
IdSqoFvLCtRZTQwpqSCMJt3+XWGQhikETkL0NK2g3Qi3hiDzaSltdgjGQrLC2ZhTdT5xs9DtLPom
7gS2NUxNXCSgM6JwMlvXibhKQqWM6nz+mWmhkMywN0akgDgAf8ajze2i2qS3XIQcRftXoUbxGGzq
Fcb6LXUXzHCJbE/AEDxFTbWZaVu4A8Wh92TW62y72KV0zvqUPAwjWjAvAYyp4mZj32U1q8XHCo+f
qoC3pch33+Ql/wMwb9FyNvBfIXX2S90TmY7Bxe+sShrzjBaQ584PiRhX9gIkAaqT8EoZOn4szYxl
q16Ld04COSVArF8S7kaLMmeojls6yWwVeb1UOyOQG44a3Cc7XIyqrwgSYlP9WlryXU1QGl5GZ3HN
XWdGVPpHrF/A8j2t2VDFiUoqyBKNMfe9K1/BXq6xYfG6dOjGQ/zQKlODYQOuT/ulcDs/IKeKnGqS
3o5EtoItMK4mLGE+4+0x/Labcbze9GU2QR671VXtI6zBH1Tadr4HvdhSDZ13AWw8yuNDPI35U1dw
5krARY58XbBDDgn2mDsi2wLWjddjeho7URcNPqqAruNNe9WCfvRHMY4fKW7mod7vHkYc8VPjIShE
uRO36QLK8GtxhzLNyDIajaT0677xtzkX1uKIs/ZK4vIK82ihZs5y7mSSfzolYSv5G3h/y3oBDLFN
nvaXxEsLxZuaeqJc910W7q+hodVSVPf6ihQuemEvlWjymotlm+9AG8JF1UhHHDLKYHHcU9NTLlmQ
bj2qYI5o8//5J6Lodtn1vqN8IJVwB42JQCi1L7pftZHP0QXSuVJiY6r8eA/vCwz6c1yYMwQgpzIi
jKECGC0nQs+By6BzNVqsMDXGAzQwFmgFGGfpXxirLUjTrXx958frSzXHcOnFCsPUoHByFJhNUUUE
17WXuAD3T3AdUQom2RZDxcFh9iP4iN7v/tRV65YEF4jyP9MNQHeT29FFssxoo2oxCOfC3ctmJnR+
51wVO9xe5bdOWlF1Eh29S5FqNbRqmitxf6IFhkufDms+aYS/iR7ZNElfABXlrncVLdqqBHoJ3F9R
O+uWtdGGfVp2K1/zUxrlw1XzKtZaNILjhPB2F5aRAWf767FPmr3Q6qC3YQ7zwRGj/T/KnqWg+PJp
UttWis5pKGhsgCVfd/zrYVzF+dejctYTJWi9SOXykZOZOyvYNxm3McrMMFY/KrEaWys/VBEG2/uM
sovGnHSOqjPwXLmFGc+6HRuD2RxotLMqbA7GFRbk3g986HcV/loORtS3m14QdvcvuQ0U/qVjuWfd
0C+m0HmlO8076SVzRbQG5fvFou01W0cxTxeBc0JLpc/8UIU7td4DRBKA5hi8IIFxvhiz7t5X/0Px
57W9gwWc5HroTOtYhwYTxppbesFJWGgjLoikiHSULIQiq/2w8m01T8jJKNugjdUCmVuiaSB8TnnG
QATjB6RbIKFUPvPbi7RIYQ4jesZyGQkzilqt/j1UH+3GWgTxV5BDhLFMT81IWrkWNb8FQYpgxw4r
1m/todKtS67n8VoK0NYuqfgsyES6kXvP7yi8MrwEuTXatNSPsRsbn+LfgWDMwKVw2DRTzIoeaNVa
H4THXPLAiWHKnlhbSCkAQOMhf44zHOC6/Ie6wKSRpjvVp1+lJryLl+db6qybjL3qNYdwRp/UL45a
FSoPPf7lwhpRFvrVWibRvg+ZkE0+I9XcfpC8msGEZnThqwqKAYo/5iJt3bU2HCNUiCCgiyOiowHe
KugCqsP+/L5aFubcBo5ahsY1V9hSfe2KvyHa/U0oxuJz3DtQsjk8DSX0TBaECt0RJm9mVU2reVSk
+oV3zj0dEhF1E5xPJQImWT2tERuW+eUrMVSWZHXo1l1v2Ak+rBRUwgChvYdfbYIt9BGMLhVHiNFE
KWwE3BoGS6OB45jg1DWugdu9imIgjEuzOXWdgRfzndd29xcuvhCRiqZROZ9z2W8Jo7UI7wO8GOCE
ZAqkH8CFb7N7MFHjI6Y4tIf+TcKV+2XQ+jBoDWtXi9bw3+t+Zi2xt+USIykD9nbSPlRP2rj023/y
QtZNF9Ez+VwsrlgfzVqx8J739GkjjEO4QOXtppynsXYywRDzFfBtS7vTHyIETIJ+HvswU9eXvd1f
f68gwaKeyfvVy3cophCXt3y8Gr6mIJLorZYU5PatHH3BW7CXmFjzVs6MeE0da9nNs3N6cjSx0hxH
asy01LDyFBMN7X0SlsxqF0PZElWK1iBXpqUYuMMubm6jJIhGMmUjYADhfvVe5l2j5cABqv3YDgj+
xfKuZMLYW+qAXUITJkZzbMi9d+7bW0ZK9Y2m/w+dDsGJxEneeF5fJnOqZVmbw4KVh3FzN6NDUQct
akLVt5kt8bELWUFDXoPV8eDOlmIh8kEQoNjD+Wg4vYFkUZSLUbn5E/9lp8TfwuKnXEBx0YXqeVpm
lN8PXHVmBR8lwRdokEXSA9xkj8NoalOTFRqsJ5Dx/Pr7dlX7jD1QgYdSpHCNJf1xfGv+loldJFEX
B5EEjejiJMd9p7bEoYf8+vdmM7kx62ebT0xTvTd+KUdwbHV4aDSMFNlDwKTA1dHVozFmO0k4Str2
3DF44RFzEGgdrq1ma4PtDw4InD2E7I1y8l8FPkIzJxenmDpm5IHdc5I3OoXouAz8/NsTEqi/6DUq
wi8BmGge8oNNRj7sibQqRbbNkuUEulsvDIzXgSoHzMfndmZo32Peyp/5bRNAUAXbJd8BvKN1Cypj
fuRmoPsfE3ez+OMWPRPM6SeGnlPOjGlIZ3tpr3mU9olPQClHsv5p4QMfUEOfinjV04Nslkv9zekG
ReW3HPQb5r/M2z7SB22ztlAyUDR2gAZIKWiA+D2j8EA0jA6WnRcY0jQIoksiwd9qYt70VWJhBvIB
K16bJlNMlz22v7q5OFxccYtDX6aON6ZBthWTRE6EBO/+7kcThwRw8VBc/uwmGLGPX6CoiMAndPIr
a1wCkmDSe+Q/V4QWTSr38qFs0bGLmCZBlhGprwnEIAnUPFjYj3ZQTp3XM2uB2cg2cS+834a0JWkc
Mf/sl8LkTXsHYmQ1a2wwMBNBWExF1kbA+iWodddMxx39xungbVIGEB71AuqTaXouWYNyj5Q+wS9H
frKAES3LfiLyFUViWntSFC/Th5hfZD4nGrna5NyKDi1CiXsBPqVhKYDgfef7uIARzEGF9ja295Eq
Ju02YiZ4iHuawQy6vDKeXYzJv0s5C9d4tmHoV1p/nMZhWT6Vc9UijBLhdQyQZELxX8IIbRmGSNLd
fWe3Xq2Ut2eZiNonVV4aLTwKUhzXLIOkOwJj0x0ClxXLjSO6O3fxrBFjxC0wN2lyLm5sNyEJCb6m
gR3FNYx98MQxu6kucVFSCY97ymYUfERm6AV6eBwxBo39MOECZMfd5s08l/SRmNuLGj/SPcvXB8Lm
wTaD6TxFLXG+lc9xJ+wjhIoycfRgrMzVnNSVeYpvUHTdilnd14Z/pUsUOWzqxWqNleuyzldH/0vJ
TT53KWYZhuASM4aaAE68l7mZ5NfmXSwdsOtg4D9WSdPjEhSYDcrK10hsAtyR6ZmRKmaww2hwLzuc
aqHzQeMIgXwC+gyiMwFS/eOM+MUoUmtRpmscQViGjSVPzkUydmfK/ZePhR+yGjJfJvoHwVd11HBN
wkVUBQsGqVf03gpe2rpEMOJrwQ0YXdGFMrVhtEMlFkvpmZC/TE9n3zEn3Pa6CKg9qfIlRS5qAI3i
2M7+ntRZiYi+f7/Bv3qR7BpPsPVuw0MOur4r9QnGFZWzhUOjwuyk9nEyhza+34/eaW4QUAobn6ir
wGbUktbsfbIB4AsE4a993UecGgYHKYYZcA/EgzD4Du9e+5TQzStZSX9oIlKMdFujBkLpbrrxWGfF
OTCHtnO7YBK9bgYwZ+HCUtLkQgb0xnzAffVfvrB8lJ17MBgKs+mL/xEukNzAQrln9XbAy2srpIqW
rl3BkIcuCG+8ea8HcRN8EVe6/wqd2RFBK8yRdHEAjI5W1BitsOKuPPPsH22UbELKen2JG+ZGVqp9
cwUlJa0evZKmIBzZVqF9zXmK6hYyQLaca0uh7m4kL1C8snAzBmqILRiThvNej0FtFCamqFYnxDc/
3tD1ANHk4avj0fkxOWcn39LBw+SR8+LIGaOnnBe/SJDJ07oJZJ4q3cABgZo3LvDOx8tFNoN5Bxot
X91cHJl7C0uBTKIwOOcJ3B6FtNEELpkK+NBBBkS6q3QJHsh4zboIIv6jsHAhdCKdHKfFxS0p7N5P
nQ/sBJazGTJki6oU48JYZig6aaXOEdxANMYGVR2ZwdHj6EQxJpIh4YihzbmfWi/CiKylihIs7bEg
6lmGQG9Ykic96M5EaLuEM8kCCY8QjjNwaxRtoumfCQ+C6flgz11VPtXUIYOQbnywUdhOTrP5YNc4
5ASj0SHk7+k2OVWzmlNcxqdoT/4s3z1kFcHFFNmGL2u6cbT4t3+gkpaHczAJXs0BMUVy69w+KkRq
IhWUYRb/la0UC4GKXrY6Vq2orw8mIvvsf4GkVGWNb5cu38Hm0VVh62tdHW0iiWzaPgelMzHrkdpq
DKt4sB08b3DiE9C+dU8vgw83MBtFRJrvfMQqtKDRHfWjkkW92ota6RhEfqzZSTCBX9L7nC9+yR2n
oboVRRir3tCQm5ZfSknV61720ng1ppdkVgr44D/9pDlJpG/899BQub6LJvJyzHcGQrhdXT8qGz8N
+pfC0ERP+c+kBbNSYef8cDSdQCIi/3+xY9pbkU4lH9DC65T0XLRwA48qUBHUvfj1dx9c+hjKFLFY
VwH52bwWalUnvpTTJrroKDMvkIknGmf+wli/OJTRdco4dfNZsB7ohtH3nU7Fwm8UBAfGuU8cxP2p
ThhReDZ3s19umk+6EBtrPXWhudtJtcjVf/AnFDi5HQKUyn5IjNhkEqLN+tLRy6V5BHu40sTRHqBa
YBniGkJt4ABgq1/UxzQEizXmGOgJD2o07Hnpm+Nl0x5OHrnUS27xGGfjNec6pM/U4x36QNDzfcxj
1CvHNWBJgEl62/7johkc8yT8jlMYVhT1uzQIHK5INbhb43Nm0sUR93yX6VWXOScsKrEuQhnBWdWN
JTMMRrH0JZQBY/lmZuZYE+jAIO3iatgnD4W7YcmVoK325wy0h/HmdiOJEde0j9n6ZpmQLssuolpz
wtiJGlDxj9DbOB5mqp1atBYnstrNBwm7ZIb5M7wLRUu5akc2vR7LEttVUFso3mDVLf8aDElbCvrD
KBQ9aEQKvYl/0UTn2okcI/8GlOIYdO1PJKY1QuJUtDj3xWB9y2qQ2+jdWzVLPalQ8SQ49+LTVBqq
vNyhc/cC+cmMTnf63pQ40pk4RPGhhcnEMy5nucMe3zK14ZGn+DDczWhx1Ecmuh1ZeAnzUot3TskP
2LhSy6fUhouz54Didah7GHQcSoLKk+xJM0k1rstlYDxoC4c4FPrDocQMzhNMbtumvGzxGz7kY7NQ
Y5Grt2leo6sI9qr0NUzxnbEAV/Tci/WDlvgNmb+bKh18YoSvEiVm+dFMc5LoI6JfrSfeA4DAJB4F
ctIBnChtZ1BuLL8y03YA1lRTvSVl1F4FsY8r2p10uo+sJPnwTrvIde9SnlD0fZWjcI49WzIggoy6
r9Wj9EgPvcs2OMoyRAqDLoQvmr+jQTE8cw6ShnsCGBsfH2ZwoWp667vFeJl/kJNNSmSYW5mXHxBw
qvgKxwn1bi+hZvFrXIkBRoPTNJ4gcqxRfLP1vpzLqq39dewppgIpzDb3qgSloFxWkB4Y56AvGXXZ
BxvgOCM1OuUX14dDBWU2cT1oEK7miriHMPlHPBRzDM2m9Ag/q0ODBjPR7uLu2hiPSBa2UrBKiQ8E
nwN7btkLhuulftqGGqmo2wAUBGnLUOJWwk7Ti0Tny0uJZuft2zCdISeR7GWXkj+zT8kSggw0zUqE
0K93ZJjHrz574WhRnNeCaGtr/+LJR9JIt/KJwF1r0d3Ha6FB8of5+0/NhPIypDfQ+R+gne8M1NS3
whkKdr3enz1TwIom6fqAbzNBpUK4OurSjtsUpZOA11jHtFphLUq8JQorgAF9lLCftao7rnOL+XPY
PinSP9KdYh4HZMq9p7GPgganK9DTfwPFoVqZiWYEMrBOVZzlXNOlfYaqp/pbVlYikhwV3cJB5Ud4
gAlyj7SufocOZrC1gHLcTAGNFYTYiiv2GPoH9yMijxes/Yg1S8h0e50MW+dFfbf6ma/4g/Asp6cq
IDECjGTPGMS4pHYLo4JoLWpieiWwDxJ6u4r8RmimtLoI/XwWMIf5y8QMWm7LxMwpCcIpaY3FSrHD
s7gJRu+NyHi/BbJsX1mbdMUwXkVqGgiVwTFdUwBxbZ6KBsMitLvD5qxsv0iNlIMiaAQS5QwoV3Tc
GzcG74ZCjY9bVXrjWOIFWg7FMlkXINFOkKlNCGbXfu6r6urrptwevLSv2/yOZ9oZh7n7U655BO2k
j2z9N+2jtnq2Anv1tHcMB6Nf9IqYcXjg7OvTvwpSZ1+gThmcNCbbNRXs6rR4H0i2bSxdFzLOgXJr
J9HA1ilfjso18pWLpEgC7i8jfkP1oXbw0aeO/UiqBGbz82bmU8AgL4/NRsSKgjvDV7zJdd/FLvfG
YuTg1aDifE/Ys1DbI63m9W7xDKh6+FEc8os30lJyflIIystnx/hByYw1jtkvuyFHq5Xfg+B432NQ
rb6DO7Ha8YA8rvzL7r1+yoOmVv+4ArW0Qiow6PHJ3y6plAJGCZu3aIsgnfrb4xnYUHpt2P+PKqEr
lwyLtd19HorgKXGpoN3dFIQEnQa0pEHXsfhD11Is/KKPWO3m3MbSyOQ6agiu6F8Km53WIbF1sZxg
+o18oD/cZqezi/Lskm/3Ysfcni0azNXZ9Jeu8HI3vaCqcv5dTomCH9gjoxNfhBwWL3E7Eu6a+0pW
OBZKlROxGPtyLIpHDwJdnnyMrcg9aDs80IxBrnYHELvP4M0sA7mMALwaju5lUkEkW60tb7I3ZwtF
Egam3cIlS2rk4CcQHYnhnATMU87TYSUayr6ONg6aqcmDVjkkJwfu/TNRLqFSxE2wnpVWjQLyjn4X
QsbtR3/zEtt1pwOLgeacyJcbChBlLqMeEGPDT6VyP1bwA5MSWYqXVQSXst+w6iTQoDlfSB1+ygYe
hwoS6rHnvozMdpi1/ZwC5vuf7+xU61TRDe3FEgucnAzuxZlljkwYRCltwUwGGOnfanYuw336xywl
MRAFvaKF6XToGOrGZR02opqBfy7UD518YEkBqatzzs0GulhJcohWFFbPf13HROMcd1d0GL+6fo3z
fB0t9wjxEa2+ur4B6GM9gjEtA4vdVI4HoM9Pwrizmz5S+gUrdTQm9XhpcLGEMsEA0tp3gQDB526f
H/ju0TRN6U7UIoIY/kfi6nXhgoguEWiIe0N5DT/Mjr6wn1PIxXHTogLB6/lz2CBxGQjrqTePgYPr
KVmvK++rRNI7JiWpJsh6nIiHf1tBloheUQAJQdXvE65bMX26Ao1VJI2rpySy7dhc5G9NHZsV6/nB
2bMYoexlE+s0ulHpcQRBKc/rVQ5h4SW68ODOjYyVvEwRXQIIQESip+gCdiXqal75rXrI5AWUv9kT
wy1BHXSdqmHYv3UK2rEz/MKJFyMjMAQ7wGvXaEaDw2vLPS3XlxzSzG4bjYTe3Tvl5gBrKw3ibB4b
8AW9FJ1qLBYPDmTey0Fk6kd+JT2a+qTmzfrCpYBVQ96qYnnC+X+Nd50m8kdnI4QE4st5FG9dlPmV
y53cMcAXuHXXYd9dF0v2ZFmGnWKBwFdnuZTCxgPiOfV1kAgnu1G3e1tk6HHGb2EedH+BQHFsy4u+
UkPH5cprJcGlJpb066KmH1UIabNS/5TWmuY4R9cSbrQVgruPUzpY+vdS9fdfN8GHLnQdCMsVaaDX
ed5ZY49WCZ6iqXIgu1zgSnR/1gGRz04BlGs/jtqtChGludA/kChsigQpCHvPhGkS8h7IdFLkOL7O
jWiT2D4+Vsi/y8io9h2mWPPttbSPGlESISvvT2LI6i4SO4GBwmtJGTLxJqd7sRZplAfftJijLv+z
xsju31mM4K1fGDQfIAtBuH2hDGy3vem2UuA4Js6X2sIepMiXJxl2wQgmIX1j3IEVxrWj7IjDRrE+
fQTZ8TZCSzNa7JG8JZSjmuAN6UmZuVV1OovBFKfqW2nM7svScEOkbjjl35otnyZQ7Jj1CFvBRezU
N39K7l+76SermRB88eOG6GmO5+Csxn2xobDsXSYmpbN69vd9e3EGUK7sO4IOSjvKU32ZWMArEOvG
WkdytsWmLkz8sGZnFDO6ZzzoOUxXAV0DkurWszxlbQxlY+naFPOJYHIfXnarAdpHNoYleFsutfi4
8ZxFKdcFXP56A5eeaFzOphZ5UmSLb4wYXj/fyc/2x+TQcNg6tCT8GWARArU4ShagBQkqnAK8AEw2
fIMm4ZHY9kw+cPSjTOOiccDsijWpAiZ5uj6fG+897ZBC1fL+sHv8kRIXa7sZvnr+3igLu05I60AW
G6FD2VnVfKj4fNdAZjVhHUti5whWxK1tW2fQ1JEo+WQfB76pAmb1jHsS7GbBgshJz8S0e/3mlsZB
+xRrly06ZN9nJP98OSIQJgUxYtiEBn7gXcl670rbulbmMdegHBgjmsU0W8g2QV9LzWyAyvEFjUIS
/evREgc1JiHlmg/Jc6Hhoqg87kgjcoAqn66nKi1dUNoG9SIuEAgHN3AfgiUcJavIYhatzph6uI7O
6hGWbDtdGXhKG2RHbMhgVxXdUwhd8A/SNSypFrEwbX5TbNCv5qwu4RHEUYHr5RdOIjbtt4PJyU3G
WNuotVZ6J/mpNLCET/czok2pI+B/cNDZCJgxAz9ZfeWH4QoYFQ0TC9ObOQyfhFyoGWBZMbW94OmX
W1mkgygm3GRmcDpALnI6icH4gQZyYV0j3s3yPa+gmyWT6FY5OMHMYN6eQLUOnXzIiN6N2e0F147s
BOmMypeIXXtH02eWoHC2OXm/ucfcHwckR4K1dGCeMxO8DZdBMLqzmcmE3OtVH9lzdL4EwemC/QwG
8qT+1KcINSMEow4oPJhcabHz81O7ZesONnYM0VIQ1y4cctOXzgACTHtg5tH4yomkXNXlQ4SgsQqi
4zCfo/nVfzeNRZSGEj8+Ay77XbrkLuGRAt7m6YYD1fGcPwMM8CId9zf4Y1KEqlbeIaj7P8N76iQS
J1oZzm4UfjBdnLyjbY9gxlZ99AdIREf6HWDiDZSoweiT+PC0LbuDw8h7UDwJjvgSn0wIYB+r1U4T
4tkL9JjJwmmLRXydw/Fv8Ykh3flkF4Im7PziBOGXApLx2hZhZMzd22TNQApE7+7HZEQi+8msL6fO
LpX7mqyemJbvLdV6WrGb4NbbqFcGjhtpt5pIJAZ4xKQmLJ6cp54U2kNJ+q/YqUk6TLRDYVK2cgOS
uhAd5Xkj2wpYt7qGP9wzeLalYTwnaqtWxJy7YyDxfUWB7yIdavmErrZ2IkuP+lBCIhNiy3fNx0HL
93VjMUoJa7WkcjAGMCwT8P9qD/909Qwu9JZWZ4jmZ9nX0FLXYWrO8J6J+nZ+7iMW6UTT7G3pOgr6
9Vrtp8pz7L+sDEgygdvRy5P3Mjjxc4j+L/ZSb6MB8AsD6t/KvR6tTQRp7KiiH+3gc0vzd8JAumXF
tlp3bxUpUCbisNYpG5vhk0VQK/5dDBPjkptZJXGNFYLewS24rSGZ4eGgY0UvHSbsDroHzsAoEw7p
vTfKN6QTlDoTrOD0DGy1nskLtwrz3Xa9BCMve6HZlU9iE8SIBK4yhkVcAIP78JrCRz/yl6ZuIjFa
ahizv3H51WAmS+7M3XEGNQIIqBxDrBcChTOXDfV0T+ML5pP66/0wvXw2FV1c/5VLDGcd9a7wuBfI
2LuC3YBHMxujNpSumYmnTugj1KG8zDyzyn+O+/kq6k3+/Gz2647+xsduDAKa2AZn4oReon7yGKS2
ogeWSz5t4WyWlJ7xOSQQtZCb8hyv8qCbyI8ormoF0gObdob2rZ957dp6FfvTayOQPQdJhL9QRde1
ocgxriI9Ai3PIbr0lKvIc50ZT80dsOx8aXdAyt0Yj9Uz70jqcGRnhrPLiKceBSx+ktlH8m1tmyd5
wIaZXw5jzH1oR/yqNbRLyinqsHx90MRNOfHfeNWHfNzl5kDTv4xk9N+9rnBkHHjQs+QILvd6E9NJ
/qp7mDybivIFWUsqve1huR83nIeEByNMJwmXGjjCW4mDngN4D+cFohTjPGfrltfwGGrTjE7izM1c
Ydi13+zU+Akn+qFAwZaeeUyKKzBk4miz7ltM91TYWj7T2yhZKcVpc+GGYQOebP1tkoUmScXwVBO0
JvUy4ZnX9cEMeUAbpNr5+ywNo1NSUE5vFdcBXCGW0VLAYx55PTVsWFgUqV82PHFO52kmDw6BxPM7
18SBj6nl7bQIt+6kKWf0UuVfYJPmZUFAdIVkHZ8wYLw3PrsoiymkUyJoVeXCaULu1epQ+YYRfXLU
gvuXAet2ZbgeXKDrzI8u6mEzir613cInCw1jQAY7I7mloXM8w0TjWCnuhcJqq/aUU8xUJulsBMbT
HSq6CzwitY3oP3g//TVJ5Wb4E0dS5X1gwOhKbLX4X+IjzZT24iY+1b2EMOi7o8fxyr55253k3Kvn
fwQj33FujcLM1hQmd9O4dLzxjjY4E0D5pXZALSXQIibiPDiGzR0lVsZ2v037SBuBMjqz7lMvqJkt
vGE27PnK5go2+gKiJhzzFXc/hJnVY2bP3xUGPMx+r3bBFUuOfuNyoehtS7X9HHLEs7WLT7RG9o2T
wR3F+yCTZgJP0hEKtKZJPqtidTyF+k60nwCa/yNt+V+LxyobMaVQ343pgJDrurXXTyeACVFfCCdn
s7Gu15rR40UWuGfdD3oHyVubkRQ53C7osBZgShMcaOMDGPTopx6XOAK1a5U9rcUFz0h7A45lDgif
zGFidoBgaflvpFjgHfSRbekSGhnOWafvDgNDoCdU1ztilai/PIiZOFFX/tygVbC3K2jqjrfpdbkR
tk5ee0J7RXTHnZti1Uqtg7kap1EERlrSP29WjafuTQuLh8tHr7j9YdXk6UPJ14CnlYeqtWdPdLuu
UKgkSqRHYaCEHBHmuVX0qgcoYc/7qOPqwk34O2oK0/8wYkoVkQYymY284RNjZ6HOHcefKJubFO1n
YeLCgxR7a4GaI/uquZsiv4N3mf/SdF7qORIlNRkQ7VfSi7SUnAHM80jyX++Kfb3xqIOlSPH3mqna
KRVwcRjXpXHLAQWhBSNh+olc1WhnLiis69oyoNUfRUqeTL2AaQ4oJuJsGEQXDsRtBtasrzt1r735
F4udN7g/I0sXHdCj7WgPF8qB2EoRCiw6B2aiYW7tHaVafDVDCOgF2DEXj2FSjBWH4SeU6YctOgx8
vtQxenxgvCGAFt1uV+EQU8HX9C/suF998/S05JP/SXqav/qLxk+r6gOj8k1/iv+7H0omANExTxV+
Rw13+kHPE76nJjqIVC8Arc/wVAFqDAQlrhoE20HitLYIahtEA6cOjpYGbrcQcXcqxNFSNETVDtOW
6d6QDHrRv1pg/h73u4b4sAompZ6NL3LLtOsyoTOBTG+lRFtmRyXPG1pD1NjrPTZSfCO0noPKs0/l
1n4SKRie/kPEHYNW0+WqG9+nxIWPKK1CbgkZ4URHvBXy+jR9xYn+sBkXMBiUTajFQ5IHX8jLGu7L
b/cjf7cfPXNdneQ/TWwfpAKYihW0W95yvc4tI9+y+8V/VOmf1xukBszOvGM31DeZxe8ZM44V8yuU
uAadWWl24neliVDdciknrUC6UddXEbluPAWhlqiUKuKjJhj64a+X+HkrL2MCn4UoTCgNdWnsGdHx
8kukoAn3MhBQUOyNQ+yzs92EPGItWncBmWLZYfWxSZ9CZys25O5AbAbKuh/jQqzzwZTLnU9QKehQ
UTKDSw12RmoPqGMsNCVXkjuI6zcCi7SLlGAq4awoNwk4WpwcFVwGi7VVZVLbVzWPFeJORa7EJv+H
y/Eq4Ty+2kHUakiQVmJ189oDbNQZrh4rzRkwgCtgYMXesdGQ/CB7gMAwcrXa0gsWn5WdZ6/CW6Oo
qxbRzlu+WUFJppC3YS2sjPzbLFJlWPmaF/p/pguqjFXyf9ku4hfBOPgKzo3WbOnniewumsGu3d8P
8FPRA40mrpU5Mj5SchfMTJVXXLXfwpI3Mk/BEzj46SwSNMOHYbGmyJBsb9u4aITa1CjkMP7WfgBc
OTxtZHbUt0mG9h2O55n7VEUSFpCYYOLBXL+cTlObhpq50SzXz2bv66KSWFedvJssBs2c75Ce9Zj+
XE8qcDyIrLU8aBveRqOPRUFc1oPj8Z2m/qFKqk/y3yvggicQ1FibBnKa765NjJztSvMjF6IONnEB
BGH+6rgNk9guTrwn4L4/vtk9ERJY6sqEQZamXTPd182UXl4qwxqT/TJk9I2TM6Rpv/HoplyFbxOU
LagfyXEKWRboLzFro6n0opeSTGk4LxNvJlD4HYJ+keNZqm3uFS+WOG7/Jmejvu6/H3fmKhJZLHKW
wBTuFVl22Nts+dJCg8IWAcpn1iWeEeeBxxPiFAKz1hfiomLPX9LvIlCVBpPwwqSfBuKt2bxe0zDG
SMamGxAn55fE7Y4KHpf0eC47eIGLqmdeHKNExX0ZwgRHoVXYffhJznl6li/aG9Afawrrp/AbYyCH
zRJ2hPv2JczHT67u75phlV6HLJrLpZ8sP7Y88YcLbfktSRndkREvEOfk0n9nkBeDIXKxZIEZai8V
t1nXhZsXF5Frij8j+drjvI3scTUIaNq3JGPJKLe8+FC3OkYmDl1HKys746Wj9zuc9G6rqX7pjpSh
cNPGnAfsxSqGwB7RzlQEwS3UECYtszyYcctcVTaT3yxYCkemC7Om2iwyp9n0I8y9c2qDSaRbQ647
DnI39xuOBrJSib4hATcwGDRxV6xwWfeAukMH+y2wJ0NHRGXWxzpETsFQ/YQL0LzV6MIBy3j6YCTf
69DuYqZ5TYML3DxZdWwW/p1kevycTahQm4LeBvmMjJ6HjcfsXHUH54ECiGdXFRiyMa5j0Zqszgtv
+1mk1U6gB6nnpIv2WEfokfhMGQ7avZcO/wlPFLuuXuJWLcP4RH284T+wrvp9SpDRmus4iqOZSuGZ
xOzg0lP4KTtfy+XdAGPe1/KYpZ9uTTmmBLhKLiz2C6v+EqPPlOBVHQ5gbYro2Hz53fz0Vqcat7fu
e+hzL3OlyIQXPBuoVlveMynTd/B+ug2Js6h0FhLYvLPQdUCcYodoABEST59CtYj4iUkvcUS0jGal
BBeISW4OiGOMoj34hMP+/52SHzKNqRX4qgyUpsBwDZiRMkz0pnG0SL+p51Y5oEmindgRVh8zHUjv
Pdwgi2lHFOMjypsTDUXWRlt6gNMU62s0bLBxLZW6xNUHbaVgSgdcTyOM1y90dk+kc3glB892v4Tg
im6rM2Fc2ieUKtjoZ9RE2D6mn3Z2ZBH6jkw1x3I8ZsTEh8qdpq6CCFaR6zi11X1mLNz3pY/dd9Rw
G9YMLcKDgstYv5Mqtip9s1QgE0hZQB2cAyaoESkGt24wGnWM2kvPP0ojpfgkFP7Hk+OUbyY+lHPj
ryjOVpE/55v+QN5j2whamELwWdlvYfKKbHJ5YRjXr+nyIiC+EXmKKeNE3ZW5/gljwOnO7fmX+BYq
KqQhYuP8ACK0/fZ6dGM8W+KUWg7OfVBv/ALMy+fK+IQDYkjfK7IAGU9V020dr1k5xhUzGHexVyes
fQ8PzYVNej9Tky6dIe5CshBmaRXTuse8RpUqhYcKKXTcgQNVoZ2ixVruq0XSVncmjiVUNCCNlkb2
2mkMeOeLlPRYO3BBy37i9oY8NtoUvwpFOlVG17KGgz+hDEsVd9SjQUf/u8d4BVK56Tj9yGdsJP5u
O8bkSSWdEDTa80QwBxshbeb49oFbWkV9aV8B4wQmGsmPIZSOlbNEHjr3pj/s7Rz0bxF1c1urlGpd
UcTRcQRw63oIdK0b3HnXjNUfgVd3lj7CRBwcO81JiVUlacoLm7bLp61k/LRHjBKOreDpc4CyznZ2
+3VOPNpFArvjdvy6RC9Rn4GbVSWMng+x5VoiHc8ItfgZfYhRm2y2SPOH5oMQDLtPA0y37TBHzmtj
Gcs8yjux/6+wels8jJXGw8pKGyxwRxS0zkL38ABrlqWSpHNfv6SfL2Q4/ufXJnXqYJH/bV9w6d6i
Od+AVle7F4x6WwVq33Zsc55F8GWgd5UNK9su/36xO6+P5dxBmMcvO6q8rLsSeSyTm4ocTCGK44JP
fDx6ewzsBi9uVLwhdGUfXKC31KFQ+bLW45itUcHrL40TGXF86+tc27aEKQgZOfFyEaILJXk9rt/S
SVG0ehrR5oDBiA30YnFo+lk2T5QMcY1jmHzQ4NT8oZ3hQL5y8Tu+e82wfID/x/Hbindd/1wWi7xx
XWCRlLBIDuCQ+fArusfi42adjOf425KuQXbjj4eiWOC9vbCa3tM4C71di6lLyt5TxgxKbY60z9zN
vqhLEp4vwrmwGoEaxUS557p3J3S8nMvhEGbjMYAk64HSVkU4mGy8y45DDZxNyh7JdnUZxfqi3Rtb
Y/X3/uDrY2Sn8WI7nEig9UYPpF4GOVyYsJBCdAgFfl+0+/mi5VM6KjScGB3C3gogeHImxoq174Id
LXgXaR99uEG70bK5jjsdrtLBhBsdoIjIE8wuVHgJ7VS4qseQvb7k9pqmxctnRZaZIc4eTSXcGTSY
nwmu2/XOw4CXS5RIa7qvuMhr8FAgD2nwTbH0qhCuKrJiHPj2OA2YSDX7VxYcxNzSugyZazBOUFa1
n38iWF8FAYXZfvb/1df3FF7HwErLiRhuxJKXooZ0yZeCA4NQI8OKkw9qDehtZ2eAz1OvorMwkCsZ
UWXfnVx7hgeYLm/oGjOVwGVZKcHyT8P8iXNn7rXj09HZW1/l5RLW2H4/Nz/6xHCRRcanZzOX0wxb
hM9iCDw7kbJ0FH2mI3Oq3APn31b21qlx8Qff8koXd1eVGJwzvEXhFHUSbdLQb5JqUMoEwMoNDD2V
imt6RDKs9cMCOQNXNZMJlrPTrX7eE9g1nrjuqUnhYnxGWuThlmKpOLCSkZSbOdQhwiw+aliOEBiX
xi1D92pyWeTLtHjPIMIE7pQanUJT0rGtKWcFfW2jCsvJFUKDmX1VdVJB0d4/Dkw6x3cVTk+IE3Od
Yn/Yer3ofUeLw5m991lrF2Gp2tOsn0/0kjniDnnwh5zqoK88d3jPsWzvx2pwclkNN0wMED60cEde
US1e/VhY7NhDgso6w374NfJdebmaI+eTtZ2hIcBQCSRu9RUR4k0TCX0PFLXhLohTFhzlm9P6mM54
c8puA56IRfPWOxCKVdMIWjKoyCLcnU3tHEIStfgT5r446D4+5LAMbdDMZHVgWrChPr74yZMd+VdJ
jK1cphe0YznX9cnbXR29SDjuIkgxUgPuF4XpyJxvI59ViX7GSl+xeE0yF2eBxBq/DuuggjtWwvnF
tA4xNrBhSTzIvZ+agJhQjp1u6ysqHuvZd2ikU21Vd6aWxSNjTcFhneQ88O1Opl+VTf3GSbGHsJPp
nII95feAjOolmGchlSDvPHYGeCJj1HIXRa3gGl4+rnwhKa8mo+TDL4evk04CPhWxb5jU1z4rgOxa
YL6ug48/xGG5kg7Wb342YZW67AC89USPmNv3CdGiK1z2Y8NBdlvpearA0864q65w5RMo5tKhwY0l
Jkts6mRQGwrKx+75jcABNwbGg5psVfkBvu+TR0BBN1VU13OVeyYKOy7lECVP2Mzdi5TI9l9k0pns
nXyq98B2mWgn8lMHTjhlyTUKoriBM41mN5Uj7MLuRW/oeZYoRQH8WWWSw5u62ZV8Pf94j8BJ5xPH
tW4mg/Q6+D+DTHuYLgBRrkCauCqqPlak8KwIpph8z/iOYlxObiyuLR128KcuD4qkSHsufoINQzvn
pZ0HOCuZ6YwL9fVypqyTW3PU5IDtEu0jGT6UeRXdC5DKzG/A50vr12QH0MVTY2CIqWp10NF49kKZ
lnLiZkDsgC4sjdS/+8JiKms1Yu4DvfrMqoWErT3k9aMWg/hXqRWusG4LSly7hXsx7cbQztTpGYpV
8Zqd4HQYIsBxmOFc/MXSM/gUqqxbYA/adiAV5CyePVr56k2iSPgW56vcFBamKjaCpF3DFjwVrqVW
PAlTvpvBmMOptYkLWogkdVm/Ux8ebpy1xh5yabR0jDvTYK4NunO36Q/ZL6aOkIFCzArXZ+qCRx2+
Z5I7Eke7J8rhHpE/wPH1Yjktb6dbewtGMp3dV95/xte34AwtV/ITqNbK6y4jExTAFbnGskdRJ7uT
IYUihgs8mb1h7Kw7ZRswMeqEnfrI5GEAzCKEb6QUmrek5ywn1biUUhDyE2qze1/b0N4sKJigaByu
pU4SS+QAuxlvneMZTCFkJC15yFjJ05NbkKN1Ufs679wPIEJk/WoNLEcTmh9SeGzUxpt/l8lKFxmg
s6drd2ESNATyx6t+/AznZwQo4CNDmjbmady4WH6BJ9a+E+AMEz8wFV3P5YEXoQ0XB8/BxnEHWjvG
ok0AELC9PuSWYE1Z9ScVvzNmDYjnxWaOW/yTaY1HvfkpXGqWCV0spgMoUgYPsznKhVMYq4VXL5Fi
bupKSLS2TAngxn356UyHkleQcRjm1sgF/gKZX1iLJjA0gMdWbCP0udbcZubpbIB7ikc0AtAw3E9i
wWEEYHU6KpDqoiMwHtlYm2xRt0KBUecdvdqemj3BO7gKELPO2CfSIa/IiMpFxNihFJVx0/MIXvsQ
gHltq6iPDT31RU01FLh9qCGCL68V7xHs9rlSlYqpXoLFbAC3j/Qd6zc9U4X0ca6cbMn5jmQY0uM5
nzBGQsPh+CIChpHrexTLhk1hEY6caTIsvy9o03r67cdK/a+H0kRMuuJhad+QV5k8t7k6bySC9Mjx
/GqFI1EQeIjCgf5HqJg8PGXg/BI4qXF6SwGuIjwI12oDfOlkV25p8hlALnSWtybEcrv8m9ZnCojw
Ppw4hcPJprlYKYDD9K97cAVFVt1seObXTVrWqp5dLvAW4rNlCrBrqblFWqIDzbQCWQJodmV6URDb
lSTczqB1AAvlnmB9cVqhMQdtIw/4aeHTf7NidjccxGT9DQh/+JPDO8tczB7uMr+uyUyO9AjxeDkR
Ceq5y7xCAhSIpd117uIsQCqeeRei47YAm5FTGA5ato5ErrHOu+Pn/MrzN74+2g+eMTpbDcf1LEWZ
eR3Oyvdql5uw//48aHdzh9k+/gnjJltUPIjrMl2E80vxX8kb42J3r9EVf3dwCVzHsSZxHkOY2xEr
++9Vp1wWvPYomqyAepE41Qh6kGiFh8m/Rg7u4WTK+utVBMwMuu9k1SlIIQD9mCj5WcvD4ZMi1GRw
Y5MoggrKi0e5C/UUz9+aq0FUVxkRQOIoU1wkv+UxD3LJ8b8Jwk5P7w0iKz6hybDxIA2bK6Hb1W3b
KOhYAuQakBAPeSl71XS6w38HvL7J91HoZfDAIa/aRKr8PAn6bp12eY2O3/UF+RuVgjC5rdROrYo7
GmeCQGhnqTCrrtSDts+iTsj/Mu8TS92f8XUkX66zdDAnnu5pJwSKHuWJS2uzf+83CppwEJHKTHaZ
Jd7w3CK5pXnK3zR80IBwOvNe5Cl2m8GgZhMTpp51nnOKnPBwrOvHZWBtIFbXLfTCKusV0si5gBvV
cFLeEeiVZteLfYufqr5nrK0UYXOMU+j/1AWPtjZnERr+wNF3jm0qBr3ms8GMjJZrInuIHFqHxe8r
JJgyVySSbL8lLuoRpQeJr2zQXR05uZsAvYgkK7waM+FihQhgFNDYelT6UsCrEV2yHFOaWKvKC9ov
tkOsfrrz1OsHfv5EXiSOOzCrylr2TdC2HD1OPjRYS+l8jNSTKcM4W/e3reIS99ukJKkYEXMEZBmB
D9XtrT6GKEL23+ecYzCPFIuQisv2e8cqp6nKUcN5N6d7o/4sBE2P9czsJ/qow8Avd3MJQeVHo3uz
dDqCYXc0ijPldxyY3I3eX8IFJSV/qFJoAmH6fXali12KMLGltJtNZKePksDLFPCqJ8ShzLgfTtIG
ANdykiSYnQ9VCe3cQSAhuS1mBpqoYohNMFHfZ6fXwXFTTxrsaK7qAIig9/A0wZkBpWGx802E+52h
061vtU0l6CosFMGGlrD5mXDBI88DmZ4u8U8I8dGMhs3gj4Sug6L5SWHrAyHvkorEnFkhQzDPe+rj
QaIcf5lyRJyrYyQsLgyxcYW5Uly1mtj474Pwsvmz9c/NX/S+rTS86WmJnzZ1tTUT88E54CUQ5QgI
dvE7XC82p+FsqTpxkGyaUBWT0mrEU6QMvBJAS7AatHN2UinSjAWAlr1LC9SMmdkMEm1l/Z2O2t2T
iEFVCD0rmy0UaNGhKqGdRdOLS04jC8lJ4gwb5oIQe/ipCCRg8e4NAMEZ+KscW9H7RmZUo6lvEltT
R+gW9MGChtwQq2RbbtLo9MiQwtxiBILhp6oQwbtQ+KH4fdEs8BXrzH3sdO7k00QbcZtnn4nTmG0q
7Bkg16nFlP1JThx7wQUSaJso9Ciq85id8o4Bcj2x/THnroHZck9d/9o43une31/A7EulhFlt3LTD
cgHNneHBZRQUG6y+M9f4gVgxfo9mBwTLsURitsXB+EH3327i+MZf1s9LukjQ6ujTEUPc4zt10GmT
oJ51MF7+Nz55aRBYNnxK7Eva8dLBNm9JCx+/C68p0aOyxdSZ/bpcLxKhqC4GyuoSTvIP4Ms+7Lky
h4/7tDSy60OVFBeRYYG+qED26R7/hkaQ8V99zm+gQZIMVP0pbSyD3M0O+VPEcf14VsB43jYQk7n4
7YPgACPjoMPEUJZC2sLtRDgWFvW6jjDbzW/U71i8kAdWPZRN6r8KjIBR9JxoHHA5uifXQihFFmiz
7IlEEn3nB1ar4tLNoII/eq96yW3niCtKIuzpV8FaWSPtvbfv/rXNlqhOutjKwKy5uaj51qmkzlP4
uIgdVVqjqYoPdP5doD2sFT8i374labiYVK1FerHO7tBPzoUhPmWcn0Xn9/86QyTQ2awvkftCakBo
Xupc+ZZaOn+UTahBmjUECizg6noB+DFvl86IxSv+HYbSQ+RP51rK26zNZXZAWUH/jmLmZiXZQH5C
qbLZxMQr50oSLZxj3n3vC4MkDwaJSrWudLzQ4H7B5p6DCsHdHv3Y9D0u8JLUmhn0/4oWclQYT8/B
x8ZfTqEgWnX2o6VB0V49YWz8vEgQ00wIkwLS9MIiAHaDYlStxbA7Y9k5RP9CVHixUAN/MSV6eG3E
67ztaHZGxjzhFoMF12++4BNzyfElHuUgYVo2Ckhp8iPzThOt+PULDaD8Buz3xb5bRkbNEBdQQxb5
vFLEmNdXEe6bBwUigGcbgUU/eVsj9lvqbhuOeEa2Wy5/tFMKslI/0qHQjO6hHsbZBV6OenD88yMz
XTwHalrQQi7G6liic6Mtin8UlV9aZPU62YJV6e7C4uJ7E/aezCCuPe9pp0dharKLi4N34j1LjNE2
ye8WbrAF+HyfTjFLdd/NpG/RT0y8KwgO7svfkTm8+AgCXkerioju8+YzQ+VQ04c38T8PVKG/R5tr
FEPgpbqGv9GjA7EJV7v4wLEUgOzw2qYCql9MWH8xjCIvk5VKA+vWF3y2uOKSAe3dhDOhOgK6d4Ap
+jUG9MkLS35G9F69ymu73flJqBfLi+NN8IGZvOKyQzJH+ewDpTkVeKa4dDPVMDvZUcUsrECaZerb
2XkhSorkWGRkP0YohGaCFwjU9z6TX+Ue1Ni6uq8+uU3IRBtsyCH8+GpAB0x4o0oymJsucAFKaFk4
Zjyrui4K78Z5++NIPOGxLlPmGvEgeCptzHqmShJwcl25Ju4vMdksXhFr8EE6icDfesvV0myxlm/E
KqYSuN1E+CO5S08G4wMhTpdp/URbg1cB6PnDKwr77vKpat8YYu+0BpELnI8ppg5SAu6IwdPPRTE0
JnvimaP8dryXB6F0GkyQcn+JKoAH9kO8F6cxO2940Y7UQX3VCnc04X48IQOGO8dn4VANHpY7jXIc
a+TJvir8d1WS/nZzIPGHijfM+5xYubeNOIkGSj1ZeQU2jB/TaUz0vCUNXrDl5hI8yL+qnTFlxXSz
atUTfsyc0K9Icdqld9KLmlVanvCZag+s7Mqs5YgA2MrEiBngIfNyh9c/3Cw1xAoEJv/2r/sS4ARE
r9X7iKBVLR2JIaPdcDwhkBZ1GMUjTWLtoGOwCSfkiSuxchO5PwCOzBoIjrLvs/PFHlEo5uz09D/j
VNuRPj9ycn+8W15NW0GDC/2i8VacZUIX/LIVmJUVgxJKzscOOZuJI7kWnUfcDkVoW53k+5hTLPUB
Urnfit+fVMftXoqZJKL+Cd+Joom7aeGckTYTbojJ4NAw9U/EajH+YS0ZAXT1N2Xxp66wZB0To4Xg
M8LpeCHKRtIdL9f0HJ+ZyIPmGbDqGxe8QnJMGnPKJegJ/4/zMMaTFOT7gZTUs7UGqg5/lADJZ9I+
uFMlot99hNQ3hOscFO66AmTeQxLs9uUSkq2lZk8wDNG5a5YmXzdypvmmtTxVec3qHrsaWI0vHVKP
SjcepzmP5MuK4y7ePr9CaBMbMyD1SP2g5A+KbmwLCxJjeApVaZ3EzzTrOQOEdaRAGWhpJ/ACTuiF
ugGjUdQLMM+3UHDfJ4SYq2ddtH8cDwZSm5kAzMc0Hb9vHmB2QA61lp08LH3+bJbxXPTbBSxbN5yd
eiNhFrFjyzWav5ZrQSREkn7GYxWN8T4BohIs3wPgjwCtvKnir53W2KQ3HQYRM6ToHxhyvMqmznNN
evU+0t+KIIfchc+lvQ8V64VyrqyCNZHXVBQrkRY9GMtEDb8Dw726EAuUtRIJNs+ZD2rgOmPgJ2fB
tZV1hMXBmeiIJdj7LfUvSf71b/kLYCAA51m4hcWfVyNpz/r89jcxkoFZylH4397a/nmQZ5V8arju
dnf8GiAA2d8hdgwtzoWDTgYrkPBDPZPhFL7tc8wp1O/7TQyHkSXpRw2rAPGqM2Yx6uIG4SZXqz1M
pgMF9+zvGLB7o3BwzMLA2rHpfZhClahpoocrUf9/+rovNrSV4XXzus589mAnkGqe1YZjedy5s9er
g0gDnDnYt7H2bC30fjXNEf7A2It7tiMnSGRKp+zbTV5jLVaBC7a82sJc5CC9bDu9HU843jkpRflI
rBXulPynVMClAfOufl7eLkkCVeEA9fMjnrPIaPpfGzZsI1LJPUsivQTg05fCeAup53OPIM5h56gk
dAxPXvFGhR5k3BSM3rWC4hB3Qgdb7gy/S+yAZCns8IrNK7K/cFNteytYBkIoFn3/skgqCl96wLQj
y814ikAyxb2E5eUuBPHPCVbJqpYsuSzTr4NcMmyNx9496X+5tZBtwQWYrZaY5UEYqDkxDi3FvmeY
tU4GDdvo9zOWJqvmhiNfiFOPyBokmVdPmS366kqTW2IKD6rGFdr8/uuOPerobUjBRsqihZhs9d8p
W6hVHrGIfnBjW1ZH232IpSCz+89cDkW8k6tMF/dW800ca+oWNAwLBxhQ9fARQP9tdJVqvF4dEycd
UEqKdtLyzqEBIyax4NgDGtA5RvdzgPpRSHqQbLjEjtQO5rb+Nm0ldbW83LkHmGfhEcCmUb4VLlvY
KJ+cmd27nZmXziIqbLLOmFRtZO8mUW98whp96nLuBH4mpdlNEAiZhJPDNn2adJRF2uluK9rQOnRl
2g0ruGo7XFDqm/F6QkJSemGzxP8/AmmgglnyS84wzKd3bRsVj5oowNfS/YytWCKZa/anvSLIGseK
RWNg7le9RrVisM0TtboBaQRZ9UOBOcp7RotGpuNP6p6mP97XFyZAXJjpXW7EItYPLvQZQ2XBTkNA
JxwkFNkwz8OSroP+M7yDKltI46WF6YcBaarA62jTp5T9ZchGWm+K/HLZCzzHjc0v8j4Q7ELnkp4J
U8HDDMjk0cbXf7gG+zujPrxBQ9tzk9OHXhOZV2ucTNlm2MdobHdYbWaHOYdStcmhcCWZxOFVm06I
BcIALMketRyS82jNjop7tQN36FYOEkQS86lXpX+y+OlGnYcpF88ZWv3yCFs7TXPFtyLv2pkTmpQ/
Yvi/lPzOg+PZhria9z7H+iV1D4YDXbb7UOiZNiOzOguty8VJ0zRXKc8ndwdwdh2iAgVnrq156zCe
7JhqX5zMBwgwrPQXACGXaJNeKhYF8xeOkN5iy1WlbPACyNp2Rd7jklJsJAdDM4PAfcXhUaZvR0gN
WrvZGpafSQhODRi+ibHYIiPNjgpVllpV4H4laGxJoDHJm1IozXcpWlCVPlIZV/KKGxXUuXL7jIdB
ws0ELWATuHBbYExLB8BMrdVOLqipF2Owf+TtthJoUx4bNJQ8rBXALQT3JNMgZlEL7GTRd++cshob
iROuwIoewOuiU06yARwGOBTS95DjSElI63HZJXcuSdqj8nHGj/xfR0FVITubEKx8oYxxMdae85en
re/nFmHhE/D+jD3hqgl631kVclx/1RLz/EEMUFKEnYYjHQon87ir69BP4Tjph5QGwksgacg7Fbwr
Tq9ipFNUMzWxhzJXTxZSysLXLXdzuI8EssvJPt2k4m/BUzxcPZF7zygtoI2T8MT7yE3veUo1oquQ
Wu6ANbm8QaHvJng2JflRXxBLlrABbBHb9DFWEcDAz3oTThd6mRY2FzdyMAowLfu20XGR3a7GmBAi
3QojU0WPr0kD0AIwES6S6vIxrkHyPSNB4Q0K8kFtuX2kmPwEgyf6cizq8r4lTSih9qDSawRByJ0f
lyT5MNLbhfhDWtgDHvVBUH7jJLiF3t74RLUKAML1ap5gc3FwxkfAMeajm2JM+wrwNlBa85lyecc/
SeRFLQUvzS4F4cEMISnigABOYGhqHjoA9cwYyYfv+gyoULEReTjY1wmjC9xZYaipcihOo59pgE0L
KqdQct+IeWz3DUOpb5y/1MsIStWrpwoVP9PkHIEP1Pb79zMc1aATRSZj5qnq7cJloG4IsL4X/Pxm
rcRnnm5kTAbs1QZ9uCSH7J+5NDlMrgw5liSf4ompdyW+7HMpsjze2CS4h85dgAuog546Wx49YdUB
CtSjWSiBByYaRgn+rEzG6I9Al00F3uJiVN7xA4XVDifkSrojBtIY5EAE+/armNLGO4nRi6ruAl/g
y6z38U0H2mHuhenY9v6V5M4iyHVD+4YlAHzP6DtFVxhx67x2bVT5zVoKC9Te5poF+KQojJVzbJDI
NTjoJzHzK2+0JZgsicXQCSs6+nkL5CxJBhoGXs8HFFOglwEZUpvY33cYifnv5v/wySyb7xVlBk7V
wEAqCPHsvqm29hXp9Tk+A2+TBNFHIyc9SaniS64PXi3s1moN3u4wtd7eyR25NIiu7brtYba5ue0P
xMAt1lW7up5dInkwF2fOdEiZs9O4YhHP23NnhiBB3epfwVzbP0b5P92yKH2VquykDtOshOmHRItp
jq/IqNuokIDfge8dN1h5Ja1zfOzq98faqrV4JDmlkMxNf3FXmCwjov3Wq4kv/XrfbzLih4XUc7JL
RkYg4F7hefCL4DXx+pkHxa7t1oZRCq4+ZlOqSsgvyGDp1CHYcmV+BTee8ybgH1pqdI/M5y2SXMhv
TFyaVoQaYR8MkRLz+MYx4O9wXCpq/K0ZfnF5smMAjdfZJfWCA/AaXEz4cXdsSJ+VWdmpagMafflh
XatG0LRMh+LwO58DN3klgh7jGw4FAx494QhftJ0YnFk9Ae7Fv53of1be6SJibU3dVlHJj+p+7ZPo
n4RptXUQL0GFPzBoKEs2lxU4gdC4nhgPkCFH1ia681bx83u4PUbxsNK1R013syFxyAg29/XnsSNE
t6VAqTKq1IUVj7R2ahi+WKfOb/BijSVRI+oZXbSpLuY7tjHjAAAbx/tuZEiuMCKN+nwBeSVpy3Zi
hPCo5jgQlAUY+ENOfA0wdOyz5yq1cRMt9ZiooIleRnOLfIHH0LwBOnAUud9zU2raftXmes1Kb+ec
rV4WXdwUFaemTPZxAWOSWyGbhJhv87+0WYM3exSmqeN7DQC7mspx3HA+Apptqegc3rVJDdQfFTrz
pKx7j7FIVMicRSYGpAryVjUOwRrwGPNAysY/BzD/535SK5HFhrutcAjRA+7XXPXRidO3FNq4Z2/7
fbvvhwWdPs2EUHchyYfNdUsBDTC1Lu3jZy/PKwLLzm8WUd8LgwUHtA23ByhbsuFXkVla/E+j4ONH
y+vTWBupHZyIP83PrLNSd1MfXoSBDy0CZermsWnA7GRMj/ACm1qbABwtfFUn0lBXICwndYKQPWBx
6vXu1Uzw4+DN0ZQUxzmX7P32jUY8Dt0xEGOaPiCVHOdxtVqwldK1goUg8JzTrgWmwBzyYaXsQ+lb
E1OhXAC466Dyq1HdTYmC8S4H46U3+q7dMaVfFvzv1mmieRp4T/tx7bG28ZHcuIbkd4K0qqSVbKrh
mKFksXqUsbIfYDUMuQxb3ajwPP1fHhdLBmrvRrrFxP1xM+HVz7xrNx0tOuli9Zz+DNt5z1PczWS4
d9fjJ2eFOAgX3ISTmfTO/LpxwqArn+n2bfdanoVuu/QvQQOlBtgOqCIJyKZUHno9e6G9x32hQEoG
KSfxFxxsJJ2TODzYSEfVh1ddBtBJGBG9BI1QPDuZG/dFF4VpiUCyDvNKoQHJqG16zs2JJUh5Yrqc
YiVnYF760bDBrPRZQLlhdHgStIy60nQkvYkJybVnhun9mIdjOT/POSlkGKpO9E86W/8c6JBNypNU
5LE+YLMhG0iV4nPUxps+oZY4/GzrXe0pkLhNniO112Z1xIVLrRPRUvaDmPyElayqollI5lbpmB9u
gkBXor5uvRSgf6I0hkiC8Jp22sWZMxwhOVGQbpm+tFZHybFSiomn6e44v6mnCI4vH3fu+wkELrqN
UaiomnsufPvrLNvzC6Vqq4W4t+fm1Pucrxqs7Rn3RuX5R0nCcwM7ZcdKFRNuBLpalm3yYgHZEKTd
mPSYWnnmEfnIxrhW1UWKiKCUy0uGNFRy8fmW/a2d1SYs1s3bsVrS/Wy3KQrHJmTfSAS5vksmAnXc
wqgk7xNhnqcVZDQhOn9R+hIkj8rDQHW0HCU3Hvo3UmoYW1weozCkSNYcLVoAFpja7r55HPxBtaW2
9GBx48yHiMm3crG1YLteYfWrNeVdT1eZFf3CyjUl4WtaR1olmyi9kgKkKh1Kdtq/uEpH5Z4rHWaM
Dr3/fZCr88XRU+I57SyeStXZOajZbRf2obbxyxq5dtpNoPVW0t3zTLdLg9UidUBWt33DRB5QF0qQ
s0ylCOHTwD/Vm34EdAwhdomLtQ9JQZ2ATYVJtoRVk0reyOOxvCa9eVkIeVG6Sio0slSJbZr8ZYps
ua46K/w2/ngzHf6JvDHeLwBiipGYIQyaFo5jK9WuRAzeTlP1GBHJTDRatRwoVcOOqdhNgsfsEQFv
SzJLamu2LVqQgz37iY0wEAAu2PY3GmDcwqJaCuDF7LJtNG2swBh6s32B8fNX4w3o6sosqEi+dnPf
w8A48Ce1FOEurEdGjJvah+CIQX3jwYmA8xxDDNpJIwUXrMQZO5EcO40jL3eeY14+8UYYE2QkeZLF
0zO0LBDKSsqNq2vZ46UrMc06zKWJpn/821PjLtRiuK/GfZxhUSgfevbRSpo4JVhGKByESKo4aS4A
p75BN0WRfK68R/6q+kjM7JpVVmFRt8J9rd3AuCapjXOvtjyRb2tnl/nanZ0ZN7zEsCWlI9xwARFP
i6ashKvaxwa5eoRY3j+rXzr2Rz+Zr9CqzSph019Da4+uRguO9XiIfSJQ9z9b2ITszm2Kox2rljvh
CKBxHHsbtQz63NZ8KFDAZinptGVndjAmI/sN3LKdnQ2+Fu5ZTUnwGJDKGD+MUrowUp5TazkFj9CJ
YSUSXGfVinarrgygc5+L7zGrOaoX4JnAJ+vsJtjYPfZvA3pcHUjJXmJbPtXvBU/cZRA/9sCQ9wuA
IOFxcEId2qPV6xTs/BA9TXGLZ0+mjKoNQt3lufpLDPVA0OIEg28XdhTOxVq3m/l3UwiaLXCSqb55
HY4ff4MhVZcQ/x47rP/MXFkXjGcHrIla0tE3dEhXvpxhscYlWWhFEJJvi5kf24whZdfJGq5iqmRL
39SGhxTP5vt68XVCCBSgCN1KgFkcqHBWx1VGkbM3Wamt4qaPk+a1jLxZNCW2lCMWVsckFU16yXxL
6YlL7MdixsuazwnEgUuZiyfI/PhMLaN4z0eyJp1ze0BAAFqRy1SKQXCazohqpI+fVjVR9fIrl2Dv
pmrNWD6WVJgqpzfvPkhKmXnXjGp6Du5upmLj1eCo+zCa5JEZM+HnchqKYs115Pnrcmquwz9UwaO8
oAefSsel52u1mckg97ZmT3VfqpaLca+gaqMepAKU65H6X/K4SzxIm7a4NI39urR5XPtDy6lNCKGT
E5yyKmyTW7brFbZFY4Mxclvr2W0hHeiknfUeFnJbwKaUQAEeXbd9qPqRmCo6dmRq1aG9R2ma8f4U
xAhHgQQFPc09oP2JmxtSy8cBvVmPi6Hu6fHITe3ScTmJr07k7YKmPU/67RqlkWllXMenTv4RFqc5
y6kAykK4a2Zg4+S9PfFnXvJd0oCRaPjSWt90wnLnpuouLi2JP1S+CCNTX1TTr5366opN06au59Ao
D3T27agjx1Y/DLD02LTn1t4ov3Eydf3TiaJmKnMxBXTOvFVxK5HwuzCsIOKRTj3R3uXIexJ6+M+/
M6OrDI2eRyYBLRRmqo7QzVI/Q6e9ld9cH9Ll/fcZtwxRYx5cyHkQsydkoA1xUeVcFeoZzK5e7yw7
kFs+//vKpsAPbh+txour4uvvn3Bny455qvANT3/zDiHtd0o3mybuZ1f6vMkhSJgoSMCCu9qQhLXf
pDFLSWU9oRAvtDTDDn73dhTiKk+YxF2pUyeFJd+eYGayuj7ywJ4dSLEPp6jDe9cm9kKc0fAIsH3x
zKRYAEXzt+jMdU37GDOW5gMgZj/BIgS7IB++c9bmFnGdP2WkpI0vRULhBa/hgJOwX7kFM/1cLbWg
3Zb6zveHqpjXCWxHF2woNT0B0pI+Vndn3FmxTp9mwneW7ym3mCv8sn+m3m0oeqeNLrsZsknSxD5O
CArubFyTBHxl6L1XInmw7XTuKjVOoUopkpa2/XF2bYc8nCTvkGOtABDiCx/sfC+ImvlP3Xop4BOn
Q6opNhv+m6QFCFJatIiTPQ0IjaNLRfEUDgls4ncae/YaYCqUwxMTQdLpW1ElucX0t8GPNBhuiJw+
YQkB4DOpKBvmraKbA2Xys7DED3Z6cgT4FPtpeZNyhdfMS8Mlig1mHeLsd3+nSgIbWN2cz00JtkXN
2L+PVz8veRbXZs88WRJc/EEZDVG0SW8pO4oFyVixVWyKvCSrA3pNxcejhruaD/BYVv1o5/fayN/A
XNtucZs8vLVHQGpsP2CbscBzLhW6nRqEb/7sE9yH7qW46cUAVJ7Tf4//LB3G+l83we576sZh3mp5
kpB58lBFOEHY1XEx4ZI6Sen+cmyCINVlwY+UxOsiys9hkIa6rlLPWasyPuJxtL7y6WgyU3kBGFVN
5JCliaYKRS2Whi2iiNtga7vl0+g1ZIpqt+wfN8DxtnyFL3S9jG5o1ODdwCNAm1EyeCTbkro9cBfM
JBwROZUqtw7BiAHvyRG1m1/mvWQ6D95+/KVgQGXmYtWfvFaOYRQtH07ADNW3aX+11lchAzTSkV7K
sCdU9ejJ3JX/oU3oJzlEIcekUi6Y2oviQ0yXHvodUVeNTiwihRWUB3ukko4kKXlKgt6LABo9LYFg
ObG6ySodZRzdU3D9XwMJnewN48UWJ3yFh17Z49irRbqfcD6oztR4P2Re7aHPqOZ5dMiOCa0DEeT1
s8macXgTwTYOduRRfSrZieyBhAF2wuzIxIIPTWBUULxobwnDkmO92OPr5NjSufkUorzjo17Kt0CJ
5lWmX2H7m2eOf+AguStn1CjyvR80w56cqi9VH5zARU1V78EMKNGY9W7xSrS4/UkJqDyIFanrzqkg
b1QkfuG8RV3N1aNDAhX2pzI2sjoVWA4xQE4OtFfkA+0yPgXjTA2YgPAX1x36tJ/e3IJmN36FKYY0
4CjXBg489J/zxWRFN4QFndTkJoQZQp9pzo5GO5sL5mC2E4ighC2GeaTSgX8ooPc69OzFGFq03WVN
mU2+PI+UYOgZD1Ri8CAsq2KkeAou/XLmK3y0noN8gPQh7lO5yeRPlrYeLv/hVl77iVtrlF1zygMK
qSi0KNbZ5oCImh+UgAdtrQuwPvVSGPn3Gfq2dBw3OxbTjW54tt5W0Dnlm5huPq4qEJshiGexpQOO
5mXEQAAXmmMFQx8wF/IhD4HuBtAJe7jcL1bxCBRhMW6sPdhX0/j3MDiE1AvzyPDSgUCDXxJ4eBuo
zgeP8rzXvQ9vsE34aQLdhUy60VGhGyCd4lSf40CUEQymKX+Lcumrq3mKA3zszFeId7tAakMGDOZk
yI6T6NKdEaNVc2vSzYaOqBBv/9EGQ8xoiaXn0dKxMjrW+EM50chXqKImm6IPx25ZitxALkqisAhe
Jofj+R830DCRftvaw9XUTWJQKH5ycdT3tPMH2W9fp+Dy7VGtxJVTpkx5YXMQkA+XlnuPRAAvVh0U
GnjiORYTU9QXNBZBqhje4myJylhqeIOb9fqhJsA3YogW32mxBue1Q+Fbx8b82T/c6QwPnMg+0VFz
SukxaxFvjaBiI/2RrEHOJlrxhwljfwMXW7E4iz7phMTNcr0yT/oFkDUxlpJDra/s0CTn9SgyJ7ye
IrD94oLoUy+pE0qjCZ81zDzSxcaWMx9+M2C6qhWVcTzxioT30geBhT0KVNCfB4B1jKkjxJypS31W
VV5JCMaSu9gZWS0mTdAVHKDrmCHYUlG42Fff1OUXNXAALEhG76gBK5vRpETP/H2aHNPg2LPkY5Ya
X/B9CsLWnPSwj2tVuFVw5tlGUH8bNG8ey+caCpETnbfY2736Elj7LDUOTjk6zLta11dG5NSNtNFx
5W8oHfmzrDQrVSvpnaGGjys6ot7jiZo19kqajpwtmTJUEt00dXot4sOoovC4/WmjwAiOANrszO76
k6hvAvwDYxjoMwcwiS6dEffEupMeaxnBqU6j5JWIcXBef/Bh/b4bVQVSOOx+O7MRKvQuPickd6e6
FgYwrMwfAS1hq5wF+Dg5TIUjC3lJVMYTXNl0B0hzJ/cVmi8++E2oImKWSS5A2dXE20TEQRZCrchX
x+X6CHfchs0ShYItjHvXaROAqJgP3hWS8ogeh2xegg2NtShXluDbTM6jy64/zn6jCvuLmhNAAmBx
OTGLXFq/YFfEfXfxHPJewEjwEoueol+pu93VbZQ8x5kwWNHEBOoe+hIedLBLWHkJqGcYy1oUO+R7
nbi8Ce9Dx2U4o5pXrWCNe2ZzOsHfW+0N4Ms929RuI5dVuWbk2lKXK2r2VlE2QAc8PZ8+0En9WpKu
lNDpaW7dCiLWRdGRQXRcT2ahPloXKUI5FURED/38PAclU2PUrgz/GpLE4uvJLc+3pbCNFDlWizgi
nxVcaEBhDhFWjj1szMtJ5ae1pEmijo4PmyJhSOVNF8NJ1EztW+r3yMhpTEUCZQ7D6a8QQWSN22jR
w98/YJwhG6gcVm+ASO0Kt+84i/a/W4m6rD8FpOV7SQWSuF6M4wOoOP65rI213CLDRKYWEpdunwHF
MqMaVCqOH7g9+OXQb6GznDFarC2+H5BBrTPOdiTOPokLaWudqfTinedDEOcY3qLajLnulpjYWIw4
HQKA2OlPVpXZ6iBAKBU6aCkRrQGItlvmG4Eui2Xc6yNtKliQtfPMBvCDq/fTxH2gEcdfswkj5s9/
FREXJemgAjZTf8VD+SRsVtMgIR2HmWOKkHkeWL3w90x15OZTaVq0QvcSI97Bx6Sfp69QNIQXM7B3
B646UUIOvxbw7ybfFTZ3HwBZ8xcSuWVBZWf9beBYCU6Z81Diazmsjn1ZHLPh0xtaXkqObsDHDx5G
ff1ejC5cyG5yynOkT6GsfkQuGTHicFrdpiHhwZ3JuV1LT8X8BFogHPZL8N+C1sjOWEIcMrpXT9Wz
WJ7ll/NONZT9ST/wbIxjKJqdwIu6X07MGbdU8teYvwL6W3xw7Ez2My0DcZK4lBnZmL/BBffgk0Vh
85dQO/3OdZa3RDxPEqKZU4jBfLWl6kVGEy4etByHVle7Its/aUdPtb0Y8pPqBmquJOcTIjAMNHXD
SKAtdfQtXrIdK/yhB6ugWFl0biau2SRZhT063EkOdU62mymyOqBs6k6xW+Aj4eIokuigUNAcPfkn
ebxVfyYogYUZJd02mFcheWzYKU5jLRKLKAYbIS8/Lvlmkglrxt8m+UwUl8sGD7eQJH5K7tYq97Q7
Hfs5J5CVrF8eXeLDyhGdYJ4NO/4T3HvQMB/ZgWOlZEx6wEyUDunr2/9pLcPpxqmIUrH2TmwmZad8
FlSFyCxh97NziLfVCx1KuEXxfXM9d7DM529IroIZMbLwokR3L1wrZNhdAjb101D56bS1Lhkgdn46
H+JM9q/uV1rQ94wkX62RShPKteRbOD2suHg/2DfREym0Rw0HJ/2t0k4gYA5HaXVKLd1RYdxSI8s2
gDnQSQJ3v1Ka/A9RHoCJ/gMlFgzlsFMxf4LqquKUBg4MaLcVLGGO/+oNGtZ6H2KtlQGe3ijerNsv
n3aaMiBz9KlReCnOFMy9dCR8MzekLjsaU4dkP02EhEQliZOIQrZ7U7VaxlNs/alQ7guSeWYWqtoV
GmxdqkG/b4l7cnTiL0WmN3ZYvx2egyTqQp8iu0rB+2CeZ7dJOypLylpKWk672wZBr2kekMiAI8fI
ZdjBOw/wF3IkAPsmXTPxl6JyqMOtneHwfkyHsuG1QJOpJjaRo7+OQb+LbO0VPkLayrl4mCPNFF/B
tJ0BW4bYMsMKjLC1o0AzY4WVI5PA2UgAPjqt9Sh2NuOI4dRgyatBcGQ/Ssqhc18vpL4xG1CDM3+k
kd3LHbQO755Z6pqz5AzdM8s1sLSoH59fB9F0TJ4Cchz8YVSrf8pZLyYhcZvX3njr0kmnHbiLSVpY
5WFEIlW01shcYUrbEzebCca8OoxXrUYH66bAJs9f04lUuWQMaKtLTLLCuZlc2i/nViyHPc4KSpLW
IVVyUSEgaK8OaFQpr+kHs9/rrbSX+WKFgFBa+J4dWrsdfZZW9as21qRubHzkllCSW6Ad7ID+ZHj+
LtIiWbbujjPRiSZ5BOXPYLbECGyxLCkvPpXR9hLExjPSjruUkUO1iC27UyIv2ko+WV46uL3kLVek
AqrLmaXVpT1HM49G3pWPd6U+Yg/03+LFi1PXd1JxYXS2i8kY50akSx68juxpiYauMYLcxGm2BX1e
+JnWifxqm3Z/1A/+Z7Dl7m4tJGdKobivF1l+t3IJE0VGFygdiT76LBBvsN4aucoYV7MI5OW/2IbZ
VoHdlXeyKCWgtqau/3g4hRItcKEn9AcxnGgqG+ZVl6Wz2MNEOgHtVutHCCVPi9tr8avhPcMw0Kqv
wU6jv8P0xfO2cgTJi3mzJ/1jgPHd9+R8eAIdb9nQhVMi+ZrhFcM60k+vYj5U5DZtk8UpzEkL2x/9
UnrqupxHv67Qumjq/1Ip4YNXrB7jj5LhVc5kJYDhI7/wCaaGkFjux9wQCX9ciUvCnAPfGwbRKBt9
G0ZyTf443KvNN++UqNP0Rdaduy5yqIGiGsu8cQEtNRAWF7JDu8NXH7ZybC2/DidjCL9m5mDYSllw
KA5urhAZ4oEY5stM0DPQ7cQo3Bk6pLqNzxwQSfCP11aNuT5I2rj6bJzURfo6aFnicFx5rQHuvo3e
d/Sk7zFJYQmtGQYshTJCvnlxlD+Qlh/urkIbzKAcvGSkO6B6fQmUAvxvjJKAmuev5X7WVU+w+1te
1v8lU8y09VrcLUY6PkhvAO+ix8MiBWMDlGo6KnKSqjt82icztFutJM89CXbq5U/BANR6OzANezyT
C1hhZJVKNMuc0eKqUymokp1ggjVJIbWfu4TB/vt0bFddRtzAAd6Uj8qwtemtsl6G0mRG/7MN5Way
5G3r48BPAXr/De1X8/w5daIWWc4pzV9NGrymV4OnuYR1ybD6eD/4N4UcYJkIUa42AtqWkw1Eo9Uf
kzlqTrDMRoYArJSTgq1qkDpAaTdhgJXLmHXhIECeEJAm0Je1NTC0aqKRfB3j5AJVRxARWVVg4/Ij
nAlzXdRcYlVpnihAj46MIR8ZfslRLWQM8KF78iNsM0uYtunFnD9F2q/xpUiNnkJOCbtb4CWD2q14
gIWshJxsSc4W8G49vacymXBcM2DoWH1hfsDbzzFoG9evuho5rDTQWSgbj/XKACyWi3P0AY/0f4le
Qr83EqvoivcpQotrxXkY7U+AkotkDvLTkExyK2d//qM9PTgwUnet3CG4HcGfB7J+YEdsucX7ppRS
rZqNVJshddQyKK9M8Tpsi/GJ1cU4EN+CXrIkWF9J3wSwU8tgA76Ewjuos92qY4KTQV9BNzwbBngX
qF8Sh5VZRQsLAv3N2Se5MOyjnNfFslbU317YjsM85jlKEVsCu78Es+V5i3jDPiLnlcY35xeRVDmI
1DvXLqdBRkUg6sCncJVChqWLztKmAQe+JbZKybtjQnIWoEF4zPTREhpMaiQLMrZ3X4qMnwvGN6N7
KEZso2f+MGicNgTvkLmAzAz1ICx1kQhkA9rWiEIFfusU6VjE5RUiXx5bQlDRBtjgwM1JXZnt8J54
3MuG4+MXzMFVY2LBJgwd+AnwFCNTy7UwHu4ZxyQzRxPTIkTbUfZssPrLB8Tc5MBYc8sQBXp8HG0Q
qeF3JvC2waFnXUfbqO8hVcNRWIxnZv4ZeQXu8GYVw5Q7Kth3VpfyPGMUtWhR4LVzmQLQ6HFt6vCm
4hf1/xxVQMrXiXaiF0emQaK9WnqGmNOBsHrR/ihsgf0kjgwwR5+belRYIfQcUdL36gKjk/yoPZs2
ue6zOQ3CSKwUy0PtzjkbUT7/0E5eiFLjJAABfzRwpXlGzgO3WmBqC+6tMLQWhPeUF/xSz92uTrBx
WLz/uXniqGeooVPsON9QYkMldVTFBicUvGFjHTtkEhcqTEgRJ0vJ9dm5PX9mES34Qk+aCmUc1kh1
YTwzwzS1hADZ8pdP3QE2JNW5Y87h7X/WvCsha5cy+y3lEJtoIVDuuynaxBCzdxPjFUVj1DH/otdy
iucrPZljPe0q2744mbLnwaSADonQ70JgxU9hmROGRNXe7XZTqR49w6RppctyoAPdj4y+JCY51sB8
bjmJxb6C5Q0uL9/Bkp6mOskMIzAhRtFqC7MQ5Gmjenepg+bgPuPpElO8Z8ohstiz+CDwMTBoDaRW
e3p/vhMUE2zudGMc/GKSYc3E8E5bAqGUTRUkr8ApRULzsGcbJI9R/UlTHBWoYa9rBCQothJTdi+Y
wTP7C8s01RTh7WEeFHXaCGsdjMInGve76HiuvDJdrl+ZaQg6BoilwyMPkKz140U7E3gQephugZ7U
yoPvG3hh4sJrciesvQQtjGNzaB/9FXp3fo6400UbNrZbjfqN3iaOSkGlhsQdr9XGVnodfnKmR9Nz
YDQNzCwa2KCEte8j7zEJAGY9aIpx/kDSra0T2coCBA1nXbsVMWSCZY5L09pUF39GASp9u1VJ2Na7
nbCrssYA0Jhjw0qm3Ywc35DgYtneT0BzgDxHTsq/gbgSYSCagU2mSOzW38g1icLP4aj8VrhirNQ2
/RB7N+GE88miAqo4fFQIjGKPZj6haWtDQGk5FnpuAIDYn/Ys0khjiZs8P/k+NWOU4zEc85hYVbLQ
K7X2aBU4osJ+dTa9XHDOYuJHxdBG8YCxSakhRx4P+SHeXTJcF8csgL52qtHw4KyMnAFtdiRneh3B
R7gD0cb0wTGZUrrMCjgmPzVkxpLvc5xkj32t1Q4JhXUp/hKvo7ptel4z6eg6hzKB6VGBMBFzapTM
MxwOlvySOprKaQy5wGQrT/2HPK2ht682QaqLp3xzCSk6YCgfji2CdqWlx594ojMsTkVP5zVZkM26
HTd0VizyBxPmUQv28zaxeIsctI6ncNhdhJANNVO+qr7PcxQdoevN5PB3hBUBEizW5XQTuPbtxcQJ
k6gb4/Bqc56NbAa8XdVNwHjp/Ywh4pfBiKv4Ig6GBYDvS+1Yhl6ONZrQMD24mfRKb9cfVOf00Dv6
F8L4vCHr2y0D+9nkNJosV1yJZkS0jG8seJuv+GSK79MbSZ/R0pK/QH2TCM9PBmK3qdhNMFLyCvZw
sS+LXXRUgEw3UgiWgx9H7A9KBQ7l4LqezxJ41ZY7ZGJOgT4g7TKU629CvXVGSStAdRLRXfuiu/IP
5lIlDVnHHjrcukohUs1dqt40fAlY5JjlsIB5p+7EWRXbm+xSCRRu2vg+GVesOVaKX09HFvlb2+nV
xAVWi3ApM7E8uazw+0PyMW3La3WrK+7lSgCdL5pmouCmGdUmpezXL5U7AFgQBYiq4YYne2U3WOiY
pZOuozIIj/3IDkwbfsj90q5RUd5s9CxyZNsHDR1LCce+AwI3MOh6eJyM4z4akukOS2YSXsnashfp
4zDuXeZC34ouOgkbo4CWzz5K9FZU8wf3Q+4pPi476aoT0M6XNP2VG7uE2+2e+RxY49aSYxi4dxBW
L3gaYivv5/4ioRnAvGW2BXFSFkPY+JOPCSCg+uaKlgfF0KyAREa13Dl1lH0KbQ4MS5rjh5eAaAxC
1AuoaqbXB7yHGnQZR1GhXFy0IxxVHFJ2ymJ41cds91Aezhf+q1ZhaYT26H3uSuoYfo7qyCp30sfX
JxVbkotQMvflF/ejBUE5ybW9cCvuv+JNL8WO5Tumjmjm0419zNtUhLVFWZ8bR2TKo/Xk4ZELb7d0
UBVMKS4RIBJjtUQ8HivKHLyiCGFODYqN/WYMS639YFhigEYqUpq3wX/XXKqnbgL4kbwcpy8SINhv
snCBQwKasoXOdyrqTvjulrcdKv0B9Ebu7tRVdiSgCMNYjhD1I61Vo0rQK9KAIlyIyDH3WrncuW8c
4CJaiGig+xtCmKjpAulQdqjmYYjS22IChgMfWJRqNCq2aDXbaw9XjjeIeVmBcZ/Gz7HBhH8bYpgB
1M6XbIai6n+VLggSkgSV2WsMsPASELoric00pwj6NyfzI4Hnh6g/njoLlwIgBQRyCkEbwLN5kbQ8
JhqAakItnavTRbyzZj/6Y65uut0+xI3RN/nZbbRPA2MiajrhZeCTShAINlC3a+Ig/IR9qA7uzj2i
W0jtcfQCEGu2Iy2RRflh+m/39lmOmvTFAnT8wlT3VxJJySevC6MF8QK10l6JfTGMhniDEX+OvhMu
WiGeuDTp2x/0gJve1/st+rbGQrtfHD2EAbrx7kQ485l0hMWfEIHExv37+b3uDsYP7vwTmlM2yX9U
2J9f0NYLHcmt9OBzFaqBHX+5WxoLJCSZAFW5Vlal9Vwtnu2mFdrE160NeJgv2mlW/gBztQqPQxpK
MNJqHluDRw2KWeezQANbmDIGSAI8mBNQYGG3/sOtckLRsvylSNGIig6a2LcNQR8huL14aOrsamgD
hFD+vKJkEeDhaLSgmdZ0EHaOce3rhiXkdGk83QVY5zNKvCGUOCEkkVcOwi6zkkOOa3JTGsCdqn8a
36+ru5Y2wkvKaTeDMBK3OZ89AbnDyk/9Ld3wuWi33TgBYR697BptB3uvkhdGmr7jEGpocugN+QIj
pex9kkwXFWdmNCY8FBAHGuFLOXcEYL+JIbJ1WCK74RX+mv9YcqQNXxJDj7PmzPua4zT+6304oW2f
EyBF+Dl83g8OdTsW1UeOpvkET8FLtOsaUf92pWKrEXewMy3pSZ2hOud2Hd9ix+JO6yHRRDvQkLEi
wmfURHyiJmtTGlTx7wcr7/RS3XlLwEDJuOUnf/0b7WsoBo7UsUM9t6TIm8QqW/Z3ISS28da3abYW
iQHKoVsH05iujkULfEkYk79ECMQpDYaZYJu2ibB6xdaAdsROiK4/KuGF7amUngcontyzrv5712Ct
H67eXxNaxQByWz526CuoP729XNMTku3EWhwBh/K2K2u43k21m9ZaPYDyktycU1gkqRXqIfLCxsSI
lmttZYVEQbepsL58MSAIz+H4oIZRMoBZkf7nV4+WNLM2qNGpMcz7AcpjgMLXeRbsurj4pOzGNU12
CnkOMBrxpydlihVZTUAK73X4+dLPkcUA6QPlOG7ZUBhxDvk5KRoVHWdNC+uZKhBkVavQL4Hx5KW/
hz8HfNoPhNbn4teaKCDAmvFxZCL1sYpHC9MOvk2BTEQ8E7IJ7jOW4MS/vWWZYobFToaZ6SAe1IJW
TTWxGPs5DzN5N32pN+7/rjXuEolQoDm9IyFDyZ39zgkNXQg4++/KOZfTr2yeUg5TlwVyeiuhXqHe
KOkrHUbyNlOJpruX0YYoD0vlddaAyJY5yW/M1MFjff6Ulz2rfqMLta2kodgOOjtVCyswWRCd7G5E
H20Af8Y7riT/dYmA3lZ3D1rAPdMuKVG8zXKN3XWPVkvAcQDqilrLmJKC32jPkuL8PuQaCeBVPY1E
5oaE2F/WyvHSHNhAXXD77xj1pi5PWDig7zBhFm3WejvKUM89GULp/ne/6JO2jXlFXuqeN7ZTNKft
v9WJUbp1gG6+7igHxLqtxS/3ocoYOAsJ5ihb4JPJdbs2MFzYwdATbLS4VrZFZ4GZwjJv5yz82tuT
fA8zwyo5YOZyRs7ixxTpRkh8b7FFEIhbeYb3QAhCWUIkG9UoWd9JFkvLzGSX2cEkW2L0ye0UIF/i
80keuo07LJPIQdFraSGES6YG5w95rxL+UBCn8WpDxdjYiGVnj8telrrNMjTMR0/ag3MX6MMZN+tq
lVwB1QEXZWeqdxkyG64/2hoTU2GIf3jw1d/kFv5Lh+BOHnNeLMA04U8W35+aQ1FDk6z67iMf/Dh/
X3/fdd5OemWcDrnrKYD13goTr3vLIgBz3yaXsMu6sV3O2vke0Ii+bJUPVPJx3oyVUvme2c88v3xp
jXqhxz56kPt+dqzQrbt6iglG4EbkapEBKtcAtR3VwF6oSM7BwfSxNlF77Xt1C8WCPCSyk/2dYuKH
fdqI0ONmWKjUrA/AZMgspmi2M7V4N4M760lH1ZeYYlWG0Z2ofz2hcaL0hNmEooaaTyy+7koHQ/0Q
/BXfJUWSCW0s9HT5wwcLvhQc/QkI9VjaeUH4JfjoE85BXCA36B2O4D9pibexn/Ro34dV+fcaIQZa
PY5JeOxWghw8eJrCrMmfzAFh9cYz+z3XEWrewPJiMccKZSLakHAh4Y4bTBOQEeokUsUneUPojPn3
WJFnJKe5o5siglUTH3N5ANPVP24YUxMPuuGcVHdWta5Y343rvCkWMFCxNaBTlOKKyZwtYTIsycOt
UW3vFHgXo4exEKANQTF0cGQEUFlcPJG76IsSLvORDWRW1RokwLINjHejh8/rubnu0jVm5qGXfxSy
qeYlnTpBmbvV28/J6YignkD/gI7FSKZQLFnbv3h4irsxyH6DIkvMoM7m9TOxSK4OMhIWkoEeboza
FfjAiGqe6/wQfhvxgYME713WjB0kP9A80a21yxB24rDWV7zNvMCq7R1LmWnY0Fd8s5mz5JCqHL0J
KIBWx07py6UkH3MEIGZ9eATp6Q0gdeL9+AEn4tnTmHnGcf45UBtURQ9cO/7MdL5V56v1JO8LTFMn
9qm31r7SXF+V+bQG1nd+fKTwW/vVTe9ps7i28s3N0H/NXSoHWH4DhI1KuTtJOfENS/QLvXSnFJnt
28vYRPfywtN5tCA9Ovm+XbbxLJaLCXs2W1DIx0HX0O6Wcg1PhFFnS8fcK+4qp+9egiUhsGd6JeKu
O2UPfvAGe08frWEZ0lmjTVrODbzeDhqBZVBD2rWIWqZ0GLO1Y+x8YFIiNrjH+TMqmFx1c6quqVTD
b/Ol9xroqEN+tsU+StAt9+GAqk/BZPdOx0jWTggQTJXr6d0vyqhRnjbx+sz4a1Bomu9ifHqhjnyI
RVQ6laGsn9eiF6UoGhC83r5wzeb/QmnzIs7gr+QOiew2t2I2McBSRTpeLkjy6FcnUbyM60g9O6Y1
oJj4uBvkryrz1oakJcj2dqeWfy1LBNoBbeKHYTr0Sj6au7TLQc8xb+vORhpgIgH9TXOnRLuQAdqj
Vm1aC2NNyQsahsHEu99M+ecNcdK+asbRNiw2HStKVLK91hy5/UeQFPa2kt52gZ4fX9KA8hIFn0pk
9Btoc83axINq2YpLfYwYxNA6DQ994UGW8P8kmNp3SXQe7Z5b/b0g9kTZRgOHjaUnmpa79lEDNGv7
/8YDvZtpXUqLfGXI24ONC7/g/vfG385M71/LF7/eSs4tnWoGvYND1tLXQv5URQtSmt7K/vk1+MsE
LT8GqxzQ2BvbZhddgJ638fO0TpgaR9OACt8t7F3ohGnHRQyk6Qmdgm558dX061OVNbjrqx2aZIGG
JfNj8vS3kljuQz6ooarN0zrIiKnfJcEkajuzWIOLSncoWcKNx9aWx31H+rtqDskhVJlBbFk93g9e
0g08uWu0TZx2gGfL7uNnrJpDBliHSpFVz8f4nHO+8bWnNMsDcOWwpD2FaGE4aRlwBBDr3Bwueb2P
55qLREBS6y9MojwO6e44f5fZ1sNTXZ0oHaJs+dzeUOFi4jdcu75X1i2yr8RKBXiofpKdDYwO0NZt
fDD4H6PfCklDaxAqnNtRujVeJp1rXmwrqJbmEVMFfgzyn2N7ZvBmkIG2miQIInQ8k3v6Atu/LNP0
3qhtzc82wjAF65+tlmZFWWBBejq/DVFAbBzbAsQkpAVHRCFa7qGQ+sjmbUaxuelaH/HEb0GoeJ/w
oVOnqugaq/V+ONCCEsZQF2bkhJNs6PH9CkhpNGVXuyW9BSg+Ty3Uw8mff0JabxmiogVXtA3q7bpw
DEsxl6VxZ99c3CeafbFTFHxE0BdWqioMhb0XJXZKhYLmvYDuSrjf4WukyTkUHjMk/7Kst9rZc/5Q
nIBMOvBI1oKFp9ztfxMnb5iaM/SuSOtO1R00orKufM8EtgVLj395TVzHk3T6pp3yoYK3BwVwIH8V
8luNAaD1CwRoCmhp3G71hTIZvAK4/PEaW5vzcspoJgoudXS7CmCEu9blgRwjpoW1vZ5+rV204zAC
EpAO4+6QNJwt/6y0zFXngFop3eC1SS5KpsyBVEqrBG0QzFn32R93YcPxmK9ArkkNVWcjk96rCpoO
hNC3Bbj0tp09AfcQAigHLM6LpP7D2bu46vAGBGkiEyncdUAU9IXf/VS2czUvm0ICYep/hGyr8zP+
ryT337tX0hu3Pa1gdr+1HGADe7wmWi7Vf5PxyKzURnsRHUKV9p9ba2q4Ce5M4WtOVXv4K8TcSin0
enPmkDyNSwiAq8sgl/adk/N0uo3Q/GsFKURuKLVoEu8Boetzfzs3jFyjhXAWlbgflHQI2/Z41z/M
/AZEtzafAV9yKU5NL5+tykm9Bqesu9r1IBaaDxNSTC5UXXKdFlc91yqvDJR+el8AgMsOFwH+5eT7
Vr19uO5Wmm3tRHtzHgm7x+T7thKidwzZ8gfZSbFH292TX1fgAgoGBgJRx5a4B/tKmyVA04ewgyzx
JkHz4UoEJz9XsWhfboFQDMQRyGIobG9Z2EJBdFUwvq4HP+w2thS/J+dfRbh42yrwcDWERpOxUx5D
hJSjvOJWWAE24aInu6VzcBCV96ZXjb3yvkQwnSKon3vuk5MuUZUjbx9YlyVKQon7EZ0oib482Gje
qNY6+BU/5RsQaRY5JOMKEGAAQch025HKHmg6nUGM2l84PCQ2HqTrFgjghb64PexdiuabBjgLO+IN
b94E33FnpofS52AAJsUsX3nBZ54X1ICuMJmmx7S0HP7vyaxmXhWqaPmRTV1FgNuyYJc9FfrbILMK
XAHvCfuX2ZQnQqEFVa7kduzx0jBdFZxgrzHdO4pw+Q6jZABj4gZQxkZHRPtZLiA6ck5KSmRSIP4S
zKUCGOwaMnsDDJaTtdUTBZde51Bvxfgb6qJu3dJ4TZc5CpI/NpwB3uCSr/lBYFkl3SbgGC3OB1g5
Gmegq7r2/iaEYRW7fxni/x+eG+l6Gc3/kBXeAwPVDdEYVY6jDRnsVGlOC0lgmc4K7nHfRuSPF5O3
PWzXhUqkU0c7b9uwcK9OZjH8ViizAN3iarSbUcRIgRg8h6j/bVNfm3s08w6x7cl879hF8pF+u2rS
7jRRa4yO5W0zqfn7/HIDqFRERKQv1zGPvXq2xwhZYPb8uwt5oRJeiX2sGngIZscuE4hLFKlwN8yb
7AqG5QKVlzmOoUtKNPrXUfMxPJjp3X3e/4YZ2zrZ1acdIv6PYcVFjgjx9VHB+ud25MaIMqqsTTf3
PpeDl+X5ZMx0I+1sEoypPzfkWb5GttMqUHXecDcN2zrAwSdYoTf+jR3s4L3u9Et+ePULht8K2QKV
Tkk5to4RGP6o0p+GJXGQXigUEebiAl4fTorNHNsN0q4OYNkeutNUdJBJuU3DETkGX9nXw1BxpVsh
bZwixuX0z6TUJV9TA71x0wRulivvMnV3FUGA0RXkGTZfpagfXEDD2f0aMVMNYt2SrwBW82xfGIYp
wCIMSHdwrvG1AtpJHT0EcaQZ9c3De7yfV8UQmP4rMNIFCgSI41LRS6qnPXF32k8hdDqyH8CYOy8z
wYwok4CZShZe0HT2mWSzdolV/ZR5dJ9DdocRZ/4wBv+WEwBCFJZz36keah6G7jfjR+8YKbZ6sByT
eIwXhcvDj5GYO0QjruPWb8VGLB1XmS/IfnEKiv9Vd9s/a68WTYkKoMoEQB0sauU1Cw9sGvYez90P
869s1hchQrE79I0MNUM4kcjeYg9uyGv+nXA7WSTZOs24i+b6cgS125n92nEgry/y9bpsQ2bG4Lu8
j7sKwtfpGG/aAybuGSkXNeVcnCLGTZSg2uSjPP8nDJPABSuEe/eSuipW2U4rLOztg5OO0BjmqckI
/sgiak7Gqo/kIJlw/FjcUhGU8XmlEuJKMcQQj2SEpC13Iwp1d18hNytVX+3VE3AAl0NkBtoOV/lh
ddoMEAEbgl1buMcNpC+wXHN8TDjpvb87PUpMbwaeAAj/9n4egCiRsKnprIuxjaQ8IKZKtsghk2CV
ovGzThPnSJu2XOBoyKSTveEPxXY30prI/9upp9HgcWFL1npUMMCMMkYSL0jZLj/+tDkaQf5IRp4D
NsnqZtvDTD6bizyzafOOW47b71a5vziMRuX1OwKOG1IyMFRI3pjG+gpV9Cb8bPrhf32PBTl6wzjR
lHM2Jud8hAKST5wDMhUL7WAVUTiK7lPuVQiEi3rNvZBzbBimVHAfJeVBqM8kUaM3pgKSb9auNcgz
pQ3J4Nh92N2JXUtP/esu4gTapXfgbj+SxhK65RMg4kvGov3SpR9A4HPEYpReqLfl8sU/Ywr00ooq
BhszCfZWfaxZjc4ovklEGxXFtYHeXWvpMHB0IzfXSBhOsE6noVzDKDpyjqguDV8CPkBDBcodKsrU
OV2cIvnqjOwliz0ZPJph6scaLfN83QzhP4BAGFzxvLREoZuZgouPFgNYEVuC8KgfkoA5Uad351mN
KVEancz3nQlOIZJ+F5bcPdxMzS0sEQKlLHxrsAK5w4lc/zuCvfdDpQsEbDCyLXHVQDuBNsGmMn4p
JUp6qq3Sf3JudORX84EMfLroNkDjtRvxzoc2GltXSLogzEUFOEuKG6iFQmpVfIj4MI3ajjpA/ick
sOK83rdCm5vNAZIPXD0wiZXr5jGLgU1an0HAdaBhBrm3ZrTddWl0kflRjdJN53rZ0/GqeMFnQ2tO
leVFS8g9KFBG3X4PnR7xqtSt3Ahw2gOUD1Kglsqv7FaqeLcr+GA3qDaCg/tCuurQ9Rsxe9013xDx
gJ6vN2/KpMBe3hOsidJElXqLHM+BZBuBtyzBVT0S+F55UMpEpQ9pTHMfBXmjnlqy2U7QB6VVp2X3
eu3PvXXa5Yw9CKQWFNE9GpQfzuWySLWY47cYpFsPYViQUfdyxSQV6PcMl8r7aDVMlfU2j8M2KUa8
bEBZMmvY6o7+fTVBDLISXSCwcEeilf+3j3s+mwXHlWvI5xLUTZszaj+bnKRmIhDp1Uh69OxvYNO3
wY0+hsIqhfA33EY9y+KZxLIjHMdJvmFmJgQ1MbL4Lus5jQW/PvH1KG5GrTsuZr94Mpv0L/C+F7qs
FNzETFQTAuhu9bZRYDXmGhz9+c/4f1GF21VK6tiNVmfyrxRDn4RXk+Rj6Y04LNC4OR4umjFZqfrg
0CjfXkIhvRc3vSm53PHk/1kNUGnvIeU6z5ED50wg1hrpnAuUXsfLF8pJz0ZppBgrBK12m2O0u7z/
aIYZGjrK50Sad2BuDXlnFPJnsIYb7HzRlzYru9i9SnkPODJCBr1CqjAwnr3QagkbDoxJAhfkOqQ4
I51eO83J2xDAzSc0dgkiub5/d5dIzhgu6lvdDJk3ZXLqG2npAckLfd7mh/EKJEHbzs4BWgCjKQjr
ncr3RkjaYiv18gAvXrNfy9Bv3Sn/ug2sZDTGDasZmeIQZCas7EEyd7dfVJbmv7z0gv4MhOC6dPSW
CIJIgZOxI493oekMoBUq53hxL12EqEfc5ah3YQ66OaPLSM+NdwyEJIWRAwwi1M4/+SVHkEZByKaW
9WQ+CocsVEAk7ROzVmsHHQataDSzNRhTYFDGJ49Y+dlwzW5hz6hhi+S4NNZISz+9dl8NSkdgbKfA
YCxKzWH6mTK5Z5JOZDmw9Ly1SBWQyCbG5wWtgEninPphOYrMhSErm/uJ+QGhN0SYLimuZ3FC2U0T
+b1JvhDD2ns+fu4XIsg700Am4E62VmxUcejbnjnyBMVhD54wokTRxJeVvaAPkYO0A2W8wD1i/4O5
0A2tr7R2QVDRgwdRnu60n/OOMW++dozQ3zoN5WIKgShd+aK7J4e8dBgtdybWeqzXCoXpMGn8ZbQI
AiR49ri0s4RtPumwzMOs4kXxKCF+ymL8BN4li3neVkJRUL0HjcRc/UCMTKA1i36JsoVOB0UZ0uqa
wKgqKGDv3YksxMNxKzPQgOMHrbXaRrV4OLbnyoqwBI9KbRmD48+FJDvQEaKgmSqs/BjbZycTG66l
RaYyWNMYlMxTZX6j1zd2mOH+eCRgXitRw/H5zoxSJ+0H6Ma6MyVmROSxIRlEmHwY8fLbvEcoI6MH
FhvCinQ+mGAgrfp5SoTgpbgcREqOI1F++buBM0V+WhP1lPY9pphbfOITZU77g5d50u28fShteKpA
ro55BpB7+Phr5EcR/KIfX+zPN8jIUoBQkox6FRWobr0FqygFaBZKpV/JJMei5jL4uC5zQvp3lN94
r7jmO+UU/FWTdhJcn/4/aG3KuGZMi81sGOnmBIm4Yb67gA0KRuFvJRyjiDNQORTk9XfzP1fdjlIy
MpiTu623GJcVGao2Zt1g4Ld95OXVD6G5sdQQHHa5dFZFBtbj47nNhp6p1hdhzIbuK6SLlp/h/I2T
4/U8WyhkIfrJXriCnfSmjMslF4gpu3MX1klhDERckRpNIZch3ECjHTOri8deoeDjnoAYNlYqLWDT
I2JRMNCi+PAtvgCW7YlH7xhMNObUt1h5uPUa8yr2Yqjuz1X190FFJoaHVrh4oYoMeJAYwjTwKsLk
i9l09/oTDvuL916Pw0dH7sSYvXEOIaTpGkuN2X9cXpdvkSoKOi5fuNH6XPVTpMxvdYTBnZ5OnMFn
99uKByueIXVfST1xrecZQR4LJtjPDXVpKbNryVkJCYOiOU/996liCAe4ax4tDLS+e2zSvNGaTavl
TcAxSl/yd42tyv/R6U/XciKicPbN2m9xwWfxZpd0dEHbtt0XN1c3rTN454pflh6Rj5anovK1nYuL
zWSsZvxC620+0dm5OdMYU2RorZaiQwvMbTfR23V1iGz9f5vpvWGFV4/b8cKdbQQvL/q16dqAQiJj
IbpUwAmOTlo4+dCIh5fDBnXQLij65xL5ezcWDPTAta+W6Ia5OdbzNiQd6TBQX3290vYE4LrtxP8t
yqBmx7VX9ZrlefO8UWnVg/mJleBm/RZhUMf4drPMBwDqFb23vtCDgSCcQ1pWUN+7kfdaxwEg+DFK
6s25jCVYQ0hUbRUGM3k1YpJNRtvXZDPIw5nrYK2aC5JpPMx3hQaHfBniiiuktEClGTzSglO/LRs5
HjRStiGDfNfwnDqKd2mtMZhpI6MsdncZ+cR0/qkInYZWpOWYDX+J1T6ghGqY+l+moTUGH84S+aon
RtRJ4h7XBHLQGLooac3SL3B5okGluOgsnatmFo3IgdABsJh0mjT4/iSPxVfYt5RE+OR2Z2vj+8l9
jLnxgTtHMOU/l1JKhT1oHlb/zk3eyrpL2c1gDhg4Oc6kZPBVh0NapL/27b7E6vMW3HNC8MyFmeMh
Kp14yXg/oP/elbXqB1VavHWR/Yso1CpplHhLJyk6tR76O5U1K5wZn0aAV9xwdZeSMCodYT3foYPh
/x1yJcJIujkZTv0IUM791jwqaSxZcVQj9Pkd6qEwkH8cetNkL7mTiaCZk7nikqvG5YrBmntOXAuc
IQ3Xtk/JRKMQjZFEFqeLQwoKe8de+Qn9dBJd19m7/R2gnj45Q0gzFacxLEFjRJlxnbgLgrMRi87O
Ni0t4tlyUivP4CtjrCcFWAXwXTpEyqlz8K2DNmPGS7pbmSPu4UXnYjcekb6d92fGKBXHnoN3Caik
vkUWCB6bZtxIgKxmZHZJ+ifmJ16HLlRjVkA+HaW+9qGWPTp3nyCyQ6cjO+s1AwNO41ocUaxPZtKX
F9DWtlSMGr/knTkOnUUXG4pQGUGOaTHHf54X/eem0QPBJ6SHWrj087F5fDI17ZqoeuUXLjWBi14Z
DqmO5PO4HnO8wwru5z5KFL78+D0/Arr2kwyH9IArlVydKCiiHdUJ6Shch/L8JTuYZ2fDi6qAkI/F
Nx+QfzEHjYW4SDIx1Ur4HahnlzKlP6nufDTQ19RXxM8d5Q1VjdhkzYrSkOtbusc5RziE4NaHGhH5
b9kddoD8LqrvXMgJkMdGgBhjUgaWTvqnkelkTSajtYu5FjzTjBm8WDBaglSZnsaef0rtdW/RIGII
vWFutjsaJUy3381CAUPIHHqogDwFp1wKX3zP3fAuVg31ZEaVzxvI1czTQd9d70FPd/q9SMR8oj46
caYNkBxI6UIOuatyYTXHohSOvj/DZMu/OZZSuRkgce2BLvsJ07S3Lw5qmq/GaVkEEpFkVlrIZCSa
1FI1vb6sbO0yoqpPPMJnqMhhh6avWR72BdM6if4XFNM+E7/hl3f9OWin4aIUIQP4+3JGy75ks7xp
kDxImf4dCobp88apjbC4BENqgcZlE9dmp8vOojgQ9QAwMdt0FWh22w6NYdFmH4AvR3IjuxLnjK17
J5MlI7exAK7s+ttjRwsQUrGRBy0ENkXlxwZvkwJPN/frIp1wT7cIL4dJv5IFM98yIbCp1XNsgckh
QbLa/SKj7zYmxqVFzSXEXJKTx4G27MGBFTOdTN0+5jMkwwQj0a5yuB9ykTWDN3deT4RTbAnQEYEL
cMdHj60Dr/xTGllT6zlfqei4rKbz40XEc2aaMimPjhr/vsW9q+v4LDRaboktUYahBf8tfGmSmUSt
8asxpiKEnecyt2LSxYQee2RxEbILhof6VXCjHg30rDb9dqNX7cbc6iaj6vBIbJvWrmhjCeKEfQSy
4v6psCaIHvEBBJMeNDjYqtJSFuSDkrqhYRdmN0//YHKwfmP9W2Vpm/+UkFfdOl5s2tub/K4cUhpJ
EK9dWioFwI0/eYxDyAYrcvHly5mSHiCpID3IGWcspNUBNc9YwrGG8QQelMKU6dYERhK1srzvLv+C
pTSLCVzIvcrBsXBitayVbikM97sr8YVS2hn+5iAbcK/kpS9hXTlJVLb3EYCpdQGPhhaYJ8kGAifk
WXptwg/uRGsTpWy0mPP39+3dya4rib6kmV/PJ/dWSdWErptDXu6o/JOAO4VXWsVV84Km4LqU90v9
i0FbIQy5bGa2LtfpdFC3GRxENXerAU/Ci36btbMPHUjfAtMsoaq5x2A7+M4Hrni7WdEgo6rz12I3
/ar5mOTCLOex2opig74Il//8bYd+RfhsWwGf1IQ1iA3zgBPTaGraG5NAc2+/fUe2Q0YJwg2uOj7H
tjBEjwoORysXHrrDhV9IS3BKPSnvMieek3aYxkDDHayjKyp0kqNV70Y8CpItW4a7zPr3pRWpC4wi
6HwgOMaRzT2Ts9cYja+HItJHSTQIGQ8P4u8PR/89Lr3QMZ5Z5bTTpU/qrhrzOpofG68d85wzLVnJ
KakfKF4z80YMCcwP6uN51gGHPUFrt2yPZKdQ4VOHm98HGUCWlwWabAPHbeAprurjJ2N5AjRv7sEW
qcKwxXJhigZHjmZCsbsQuxtoZBoIAEMXPap24Vw97bE520q266zjrPL+Xr9chewxGtPFtXlAXhKj
s+jk23Ddsu86mzsOGKseBZ4CB+DuF120/bA/QrCkRTG2iXTHqEyIsxx7negf6lM7WhGNWvwIOeMt
YeZNbhYQ4WwEp4I6E6xYButqZFMsvTBW9lmfLOmfbVDoH+sRIZKglegcnz10nhbOU37ZFcQIXncW
n5+Kl4Cpvtk7AKUMayN6qqJi65Vm9SGVx/adVLd87tw1Dt8nrzy++L+IUWv+gCSTE6MFuXjA4I/R
JG1e+ykSdMIfKeK/cI0q/dAbblJYNcwSoVnySUiYWK5M3W1xXQx5YU+8+VzuagmA3m0lhmH/zCTE
Qwzkg8FsMHT3AlsveyNsCl9qpldX2jSjaYE9GnYcSKsImJwKDKIOkyeCyeVLzu8SBzvgkvNJC+oy
U5FSLLaktqCRQmpCCpxnkRxsff1k/KPTP8q4ZLjVpiZzRSFYUFU/JGXuUIc9Nvc2wwQUbMdqSrYA
t0+TfDPwZyD3IdBO5owRSpqHK/bol2u4XMy5o/qGtP29lP/28H2qiFyztB+fRoZXmef8gC23nGwH
Ir+9w/95hg47mQnyh2D7OMYI9YXMsXwPLxd6o5zRv1o6RdJWB/tfBDFPf2DpyL4lmWEWIeJYRaMJ
FQxNbzNU/5cMe2sZCfAUKsCFCi50H5UbMh9O9avL2HBy/mK7uekukEdXuDLTP8B2/fgs8sfxnD4e
hUNLydGyDutprJi4CBljP5p4OoD02SNJpev1SSPbsH8Z/LwXcvNJ9/Gid8Z83v0HledFUw0d5LuH
zLMtpeSagbjAZOaiiwZGmkmNWUxw7YKdZaG05AhUTLORPjEdC15etxelaxobpTw4dFBeXmG0XEvG
ZIm30bjAKxhv37uhBN+ZXec8UoEd6cz1X2or16DyuU6OmtGXgQ/R+3/2U5x7BfIVD/mA/h1tE8Fo
FcPO6WZtTscaKGjxDxnpUwnXgWHVXnG+FibIhovkX26+r2hwArPT6G7kHs5yB+KaG7s97L6opBe4
EaP8KW2aOKqcpaIF66iznvhh0xAwQYzcYXqYAtuBQmgflFL9pEHonPt8bgGtcaXlmfS/EnpYtn6A
FzPApTJelVsfAG3Fsbvn8erVpv8bcf5VB+nK6yVpjW7/LYNC3HzNHAtV6f28Qcc0r3YL8JUM5WqP
0rJ7H6PZiWAxetIoTMkzJ9N47qvBOROB65zYkmdsxTbQrhCN51rl6105sUg3D13jpZBwdLZyrTWO
5lSTb3g30HA/ekVuKfJ1AebvHF6l5vP5STgjwMfNXQ1MkfOCe1q131j42UaVmSHLYnrBeYB1wnEN
GCt2Mm5MoBsXU51r/r6rCVSBCsEF6GIhbzSk0oLjAnhxNcSYvDMylFTw6iBPekJSQoyikNq75Fp4
f/fsXCnN/iglD2D+vSYb7njL77NUMQZaUHLDLJRNQpQDc10UtcqrtIgtCa1AKONj2EsxlZObebmC
V3aelEUnWbgIJ+6Vy7fS+lRSxVFBjyZ3nO5MXQ/mT2aeHwchysOTcymcMQMaeZ3jMMf06TiL8LSH
VaBdosm3iJjSMeMOebRlyb7QiKv/oE5+HcN83Q2I5u4lImLv/IWh+/NP9JLt9I/xz8T671F8FSX0
9tDiVoblICKiqXwTUDiDnUcoi0PYBsN9G8AxQ/7la/9EnxfFB8/L60MLVOzKLMYGKAwtfD/+4p92
iIuR3KfoMOnSKgfvUjZVBzUya1U+ZAQaS96XNIfzLN3xqNyyV8sarDEobdAchbMflC/lmVUkJD1z
j7toSLgF1xpC+j5Ao0A0cI24WpVX3TEd1O7qhlNCbrwPa8FF1X30/uNj3fYeI9LAWJNvL9wx7zWQ
f4LI7afMH+S9Lwcs2RNFDP1W4gBO+9+soOzQ32NYH9cIo0FqC11rRS2ivjflIiJE69zUHbyqQ69w
KfQnh+azbRIm0uRoX7pgoesB80zBkFqwG1JpggB77N9hu0WuJHOcDKkB4/0E2Z+97wgmzhKKdTgG
+oifcaaFa7fbKCtI+cy/MP/VtUzsV+CqucvTSiMpm+8LFgEBOf1zY3bSMJDp3RFU9q4rl9T2mg+U
oV1XhzBeNQtnqxY7xqPWora/XyP+dpUe6dpHd1b35YmPa25Yqgo8UiRFTcWH9wcaVZhtYPMQBdGd
Fu8bJiHffvK3GFINLuRwnd7T5ciKnLSAusNByIAJzFgLn789DS7eu9KtXK6y+96ia5Iq/E2E58IV
Of4xvgiHH/yt0o+NJYKEL5RrVdNv4YlRHf1ISFdyut0gT1F+pcdqyEUHSHfAyGRuX4vbzw0PO1OB
dHbWqi1vRCEBBH9CNwnxwnRi2E28lcbCsWYx5ngaLtb+fnG9zBgvuB7zc9YZfQoelMZDypR/fwTX
1OjpegWQPbd8Ey4m0P5SO/jbi3WOcTkf0iLzJ50vNGhLdvbnpBWfTm2fSJTL47mJdPZ1Ign0Tp4Q
ur0oE4PfChVTzXJirQTc6Ks6M0Sxf8xwoHsx7nkMOuuiSwEeWsR1XgHSLMI9ZTsItpcduVIApYtL
O+zvYnuXgsx+EL6t9VJyQ766/ZMTMYimT7DQAzP+7cx5QyXw/0ymbH4lhFs5RnSwr29bVt45OLJn
ZpMWPwpjj8fTDlEGiEjs/lhjfxeajpOUa/2T8OrgxSuLzCRdGChZa5sFt/PwOBqP0AL6/uPWMxUq
QEFRCewqC7rr6XWVnrZ3RJ6EXgNZWk6Cr1A8LrbKAQIpxVh1P82O2iESHtHsuM6CwUk5y1ZqtEXg
fGIsU0icw6vuZnpxirUvxI8PB9Ypt9BhlMt1eP2Und83T8lNGnsjMlpY7zGLPShvz1kg0SLej775
Ajp85bbrUVnB7kOea2K60aDMUdYOAQD9SMuNuATfLmY1cedk5ndSWHuHOsD/IoGzK2c81szkjq7O
U0dH2hr/Ucyojny543tZ5lumoNt+RjKhlzVu8Myk7f0nIddtWLyHcDENqknIE8x5818nOlCiqhBj
JMpfUijrrYeZNvQsYJ49hvMbVdkccDwBAL/62bPy01+bKrlIXoPorpSquPeb7pSfLT2rB4s6HJWy
NSq+QS6I/wyTsL0g4DCnkYg/qDKXrLr1f+2UeALe2SpQ2wTIDwuuHVL0c06VMrnfa7PlVb9Xugfs
a0xRbLXwQBXO11xYQLKt1AFk7Yao8Tktx+DjUkqR4aW5QUnOTkwlYlnaK9iE4jxBOqY62g1VOWV2
geC9UpOD1FpqROUWZGBk+q86IRd/W+eSYOMThvNY0J2LjDHV+eTnwP+2fdp2ytHlXMXWkU9DxzZ3
VlWO+sEPc8zuNt8Xay/7/iiIWqsXa1rO2g9LyKC2iAkO+tJwumlZI8C5BKhSr+8w0aKdjXTZ6wDA
HQqg25vQQlglq4PcUhmVOC0ytjULowSua7sQBmHbWCQePb/75mzjBiRSd1++8Ktomhe/3yPxfogh
MBLglrAxeUL6sf9IEDF1vWmjk8YtKPQVFLcIbFD/4WFdPGcZyIQ+3JJJH8+DU5I4YXy55zRMe53L
eVXRL30/btZvrSLTImyTfgg6zymRP3HtE3eBZrze+JkCADAue8JFnLoQb2nEZADQy1KngVpph4ZQ
+CHfg9mDdkqczF0Ul1A0QFLXySe0VMV/kGjZVlWSqof9ErTpCUFCIs2g2p/3PdDW13lfT5sWKP9d
V9ECH6mwUY0rrS3VEVkaDBz9QrhhOKBHkesJibcvNRZOwN9JwNry6rcTdsW6XiyzCRtQYVlppvJE
IVXlRbCNKaBUm934Wj3r0krTtq54g3j49t8/0DlETxsQqiGhtHx7mf2N5NMSVdaHSdaQNpMrqu+J
r6MAG/EIyJKg+6e6SSW5BYngg6m4GRg3oDEe5a7nwQ9bAUzlJjyci77OWH91kZcKQrWDpxdaICLI
U8B6c2V/kv2TpCn+vpkfPazXqek2oAQyQ36WTckG7ueCTtlR6x09A7XwIEel4Mcn+1BqQubOjIdh
WfCG2MYZ0UFDh+wFtgwTydCnZd1xhR9WdYvn9Jwh1SOIuTwExAIJTi3Xt+6k6XmNHJ4GS3clQunw
rrDWHWnQ3nGcQyQiGDfSlgdd/TFxHoT/FYUvCo4sEZCZJGcHskt3iQ8wdUBvyhal4a5syQdGGYSn
01DJHwd4ri5YqPgWCiYVvB70j+0L0APztvLt9k0PlyO9m45HcyvpJ3OvcrRDWWeBJQXA0V4qPxta
AJuVNmzjRPhXq8rVrGy72sdD5Uw5Vth13P00+oopRlUpd23/lBdkilO5Ivb0zoqxAa6Il/Z8rHvH
xmVQ3CMOgAVRkHuqlnKHLgb6elmuduXwVEfKpt85FzIa/dnkfUhbrnwHjtEv8sxRApbqUu7F/Keh
qNDYrZoWM5jM8/VxjdKRkoXCX1AfOVwVER05ccgaKt1Csmne54QTom7JWRXG5IhbP+PQSqiY8ZCa
8GIiSFViGI48Q4UryUFdS1evHzOr7fptIFngJQVnnuhCbRKNPezV+tAL3DI7tZvSrIXbLTnPIURk
E5qo8rEiHCcVYWTWBpvza543Ks2EtFhrBTzarFXJ4dmvVb4BplfO/Pzlp0iIs9QDOD8CvAH59LbX
BsClXVuDeGYyLuqHnLicdj9lZDwxxbw5jmfkI1eImsdHncVwsdU+odIYGyvxWuduGmPDM2F+Ni07
3I+UbgzF9QomLB+Qmw9v+z3uQNccrIffcClQXbZH/bUhd4Pr/FMu5axndwOwkJjFfLAmOwdSst3/
nFNAUuiHd3vqxh5r2Sy0XyuVN1iFYb1joQaMDOP5AIWwQw8Y+U8ErZnuDaw1msbYy2ejEDKwz24g
n/gfIWWn3HJRHC26d/m2FZT/FSotQqsJzwCwR7hm/VNh/RG3sKynyJDa3TDF7tWxkNkq3DigwNqy
5+RflUodQi0d34XOI04xtXsUXo+AL7IjLv4mvRNYreW8BEiLLO3K/taoDrVC4QteWQvgUqe40Rcn
JCAmRUrbvnZvykoXT/DInb/En2x6mIoKvBTTTMJEK6f02+vskedpKIMuF+/biEE1//l6gap0JO7V
dGJUKPBikBcgopt346SAhvz/53lf78Tx8/LAV3gp5W0HrtNqCM3QXHySluy3PtQ/hX9lsqBe/Ztg
CoEutnMiPlucwqKbFdta8gXp5gFgaVeRTgvBxCCjpj/4DmfjqxgtlfRc1tLDqk/uC6GDU+N8GQei
9QL4XZS97YM+tEIp6ZhULxtw2eey1I1YH8B23dm8jy3ppP5Gu2Yf1oFSlCXtCuttNu8xb6JbJxFz
rkZB5eqxe+fslRWUXeTwkop8Y/a8QuzHXl0n+Q+fXqrFlHuUaUPLgdjm8Pl1sW4oeCBohkFxBgBg
cfWXJHClSkjpynjJdcSEi2dcpbnaofwQJMtrAGbtsjM/k2mJzWt/K4GRCQ0Q67ApkqiMz/Y72t3e
EgdwarWF/xgPiCol+dBJUgJbqFXnZ0NIlCU+p51lARfFHFLPr/zaRHAsEKxMjqSqd387b1n+tJQT
OE8VJ3ymJQGucCX8g30YqF8r6EX3hCSpL+OVBXz/b6kfYfzyvW+6DK/oxkgUkCO+ae4enM8gPLvC
JMJR879z0bF4hFFle+7R5k2fJfp89X7nDRhzlnNsVbiwOS9FKbtmfEJ0sBMAasWgp+tX1od9MUXr
DTJFWHFCTn9D7QExiyJ5N1m2fX762LQ6gV39+0nQ7GE/7xcpk3HkQPU6XfIrWF4kgAVYwIvRlxrI
o1MDDVlwAzBy9+WnG+/j1EzGjezJSRSp36ZxoaT9QHuSJd2aHlLxCxyVdecYmXbtRtljdaFNFUpw
MYLrsGGceJMK/dhbebocTCUk7ymxQ469NKP0xbTPkibU7JKF4L9YG+hua8lhRx1xw9JC+QuxvfEh
D5muj8WGYSW5ktaBZCEfXHofh9XnkUuoYDWMpjDJf4TLDDxd0GIziWBIBUpVqUJuJYCYu15Z8wY4
R9swVu4uL4ywOyGdPUzRW2cujG8RUwjUhLAfMaqS++4BZCePHHlAoLFrOMg/UUsKjYj+9uh9n8Xj
QgseeOrroFGhkkqolC57WNMhkcaTnPSbrAlRvhQy/8pXX48J+6+49X+/N//8PMxz3pwuz1Y8OpT9
ayZEZBXk6cwUItD1vcdM1kuX36pl6j+HHzqheS5IcdD0lZtlAAvgrp+sPHTrTLpeCPRHKcZ08YjY
ni7+LqcSUBF2cb6QQ6EFsBwKgaDCRC5iGAI14wGG3lfzB+uZyhGpzm6g9bdm6lTbNaM/AZ4ZHWr4
uLQbnqTgvh/1fw1b5Ji6RTojRrut17e02fY22MOBMPPEoeLfRTdGelDcMiyTBUQlqcmAPfDv/o3e
/x0wptD8kD7yq8gNTOLywbEZQwXrxzbVLTMJ3wwp/YPCFki2KVY0cQbiAfOQ7pEKt7bj5ZVb6b2z
oS1d2DmhCr7VE5XS6rctOAYRXDGARHGYQ+a9Djfiet65UVX2TkNWmrmRBmU+vwrhizSQYvnrS4Vz
XRleC51aUTzU9RJL/lyRrz2o7LTnoqQoFwCKY7AQy6uf7TR15jRfipkKKMe++EyXsOtZUCdoQ61Y
UF8XZlOqIkYwg/qU5V30ctww5IqzgLoWdmigYuVCVRrhCxbWk14Py7GyJPunS1GrLx68SJs84WIr
WswSy72otVEXLTdAmJ2mzQZ28FvCm21xBvTTVeXffHf0S7qz0S9J125qTCNfhrhwHFSau68WHxtY
H3X3nvJ0YiU/9juem/cEAnGJhK9QVlosZs2xrCtMpmjwsnrJg4D0ZDxGitr8Vpsq8o5wRtt36x9M
oEEqG7cYKofhxfDsBDUGSAH9iEqT6DsdqMH6/u09JWO7d7pWNyXQ/oMNQXwmHP92d/GsvEJUEVNc
KPjedVC9lpDNunguWg3eZ68S8D6ug9Gk9MjzPhpvh8o+PpjljLys5JzS6ZxWlG50AJziC9cFP6Eq
mrEaTczYdrzHJ5LRRsOshqlEyzGz44uZxjWt7zrkc1LULfRsko9EYO2kOmd2MOXS+qH9JSPJVzvU
qyO9u2pwBOVd/aIqiQlassw0oK56bTQcEEx2tO/FJi/88Emx9dmQhOu8n8pyF8hC6Fd4HiTCGNPl
WyhjuH4YykMsFto98IhF9sptMLKSJpfARUgiX9/Dwoyp39CCF6JDExRn7T6eA/8Q7V9EJRL5bSyJ
/tsAKezSQaQ7/auTgRH2S+KtAJdZLC6n7EIgbbWUr58+tFodORb1GA1MGm0GYf5NcrxSAoCtoWsd
9TEXHxMkFC1vNClxH8w7dOZnZJMflHXHi+gGEvaQxfSLj64ozxbgF2ciTq5Vcin7xriBoU5XTpWi
uqlngfDM+gmMbFbWrNclKoJuEHbAcN7wNhEvhJgH7ZWx03xpr+q3DKmFWzvv4mpXdqoribTApvhS
FLuHldxoQVZkSD9RgLa6DlnobwtmoFHyZz+i5muNR04pGvpXxXQxYkIA9Md7Q3+QAFXshZZDjg0m
kb2cqJ5hE9JXXeFjj0muFpzGlZaaahOHGig9OnDGbvKtwv6Rw2c+OzPHqukoTmk5nRjSvvEKU1eb
AXcIw+CrQ3d7Lz9Bwnr4zoczRQitR+/dcguLeJIDrXz0kwQBkS/68GRBkuseDWGBzAAjTQ4fW3lA
FgboUvFx2WOTJxOqeQ7dYMPYZqzczdx0FX9jTw6mq2lzBb3TAI2dzIYe4gN3+7g1oSr1dBB9dHUW
Qyc1ukAq0bPxxk6P0MtHP7ptV/00EQOppLmm5AxtckeK2QQBftFM6OIPZfPfPm2fjib/SAgQOV2O
iGg/9M9yGuKylo0a54TypKlZhbHU7fIRYcSGN9uJltVM3lxm6jtQQnEiL026x+5HRcZ8g5t/Cln3
aX9Lv4FjdOnDTlRG6vRVLccLGUrRQj0RSrSwqE3xTP+Li525veywGOzguj72XciHj3tuuVmQ1W6T
ENNnBrLQcO8dLVntKsFm3jUUuH92QwfiHfBsbWNtlMI/GuosT4/S33tqssWpJRBAwAi7TSLB0wR3
/t9Elg3Qk1+U5wYpiHXOmVjDYd8Hq+8GSHS9+X0FXv5o1/u/3D54e9yYjZFuiLMutbRZfkaQNXZi
xUmaLfEJmKg1wCdTPJ4SPP04xs1+IqLbe3l+FVPlp71OG2rnuddK5ptQG4rott/aUcPC7MdSZTJW
sxcMFE18cKZeKTNuLhBfl1ViuL4a7pRMVK+I16gICjb48O+qdSqivPbpZYZztPXriAE0K7d6cA5Q
JEpEa4CUyNKYH+1gTQeghCVPCUNSmd88YNrO+4M+/aMdYxh52carcXDTuMVSuqZ1Wzz0IxYUaYyX
QwB3kijXD2Y7SbmqhO7s8lmSQ/tChwcWuz9+J4XitF5SS4RlVr5PC7H8iLIhD8bhKnM2ubJfDCT9
etU4Q9k33vLnUJLp0O9IIQXcrMZ1lSWBWYl1QEyXRtPkjjqdNS8U4R/oQsS4j5xHhd18I0gFRw2g
A/O07Eta/SBJcOub9MOxBmUYz+/0A1spx87lI9cd28uRCTQZJTskUGDaG04GRj1lwFAqOwsrt85V
PkxprVedhFlN15FazK4eUDo0//85V+0Bo4T886TiLMiQI3s5Y1QcvnsftKMftq+isf51VPIhedrk
jSKMsAydlVS+0RfY1janMjYxgKpUgwNhf215Vgatal4BKYKiJ6iFvbNDOcyIP1relrInEawDwQxv
81pyWgFHRFfbZHioX4dgsWon/gmegQkd5zQ59z+B1TaVKcBw0SS6Ld8/2VSTnyCv1VQuX8qGikk3
kjAKuJLT6AHqZ1wJYNyhO7WV+XeQzv3yX+Z8sZy4RZBhTNwrDS4DortN5xS+7v5+TnkeZ+vW8sTM
IBOGFPcJH7WnE/L0iWKOTjfXmuE4vbmJj3Un+gYEMGWl4TmxYbyrBn05mwfhZxQHeQ+Zub0Juyik
7QenxCzfRkEB39QNLm75KdP8SVvzBdoqCy+/Iw7z00M+Zm0itrHGRZRGR0FqDQghrLkOzDx/D/JA
EngFxCRvwSaGrRRegEnXMw991MUjliAbWHLGVtcnJ6exb9BKMwxIOCa3RJBd7pupigEgpBh6yztl
bBBSIKANjL7Rw97uS9EjdEiUsowJ8/gKk2k5dep3nr2K2qAzhWVIdMfGY5Pa4LNFFi5MMNM7ksun
JF7YQ+4jUTcAltINQ7bczeT0RDN4ClArshR4BvKWTaj8qv6jBXx0s7OsOf87JpY8bm1xUrDqOe7F
IoHQkGfmSzCkVzdjxN29TvR2y/cRiaaG8ApE7VVoUnTLS55MdsuxPaqLb/PcO4EkcvYYiU3criIO
xeesLvZAkvSIUZdmKzAH/axH7m8lSOIV1d16aUbkAUHfiPcDr7KCqeDXkBgw56N+ytHCB9GrdT0j
WBLi3wZcqhCmVsg7IYA2QiFkS5oS+VZTTIrjdF5pp0gQ+yeYytuW7ZpdQ1Z2VzqxXoT8lZIOyyMO
6u1kc0oXyJb9L2ik4saUz9RPtx8zqCDiYdKLZ0fkFEKplXH5J12r9dD3OexG0XZXtfCVZjLUk1x4
ps8nsxhHb7gvkn290Sl6A2fA0ht9oQ6xmnloyJrG2F68YUvpLwa4nvXWyoa0Qpt3nqdg5r9PB8ar
UIHfwT0pE8IAM1Ld7p/Gs+lKAbTJBTWgyDy5zk9hv0jdWaIWYoroiPrjk2Du1LNBtK4jE61aNAI9
oyuKsWr2mb5VijDqGpmV3RBhoQkIfIuTa9F6YIqV47+sAer8pQoRpMndUL51rheO92LjDQouHyOC
JcyyjnJV3XkW2cTWcEkZHlVupf30+R6oRsBpxaa+lOGaamrqYclCtZ/ENF+fRb2ANpJAbkqeUCCA
w1gKI2eR5AKgGfCfykj7WhIAhcaBJHNFa6L3F7gyg9atj7YaAtCLkzvi8enach/fC5B8Hftdoopr
zJ+k67BBeKT9shECFKu5+45WlFe5l8tc7W8ZMtJOPf3K3/hchucRHirxMeLW8Uugls/5lcGrF5WC
IzE/cQt5kWBIlABj8iyKKpoSvvVQyEbwcksFNaCLq3vUS/2l+yDCzrV9KzEPvyYsD81jlCfsFDS/
+lqJxWQ3vZ8vEL2lUQILDdL/reDCUxMzBibL1fNQFk+FNXDs5EWA4edqPV6rDLln8tjkDvqcAbqk
obcHTfqn//mGBQmR9NiebKnLr6HM/AuOEQTNJSy4x4c47+ZvUtlEVF0o1ytG3q9NykIwZFP6BFC/
szxbCLZHrACkznQ9YdXsTCVEtg66cKi/WfLc1X6V2E92FXEcG98mTd8c4es8RyooR67q9TQXwOBV
rit15qb7hhy/5r8s6keYfatW+qfc8j39QW0E7vfM7Ys3z8Lv5NZe8bCnTGlX1HiQLAzL8NbOnzqr
dq5gTgdtnfce25uQnF7TV4JPI5vAfRJ2UhLaGTmZxQVdFxkJOSo0nx4ymDaAPokQf8cZGf7f5uPw
qPI4h9w6L+qxJ22nrRaLrlXrJTiXBm/0fJeFBnSUZjZiF8v9DH6/Li4tD+F/Hfnj3NMOq9Vr+qZ+
3RWgiw9jFTsQzSy4gDNX5uKSFewmj1/9T5IyHaAv6p+0ba5lXMH0rqOjNFNEeMzC6qow4dUB2WMz
kwCGuNlDJ++vlDAzw60vlWOOAs56BJ042Xaj5nU8I6g49aYBwh3UsqmmghNoEQ5DoHAkAdfXasEE
C3MXXdFMJZ4l1k+b2fdzbEVG0x+FPOPbtvl6STdv//q+0HcjffGsAYDqdp+b9dahpc8BwmmIGma8
lh95wkwwsS5nasnls7UyQqBJZj5yulv46Vc8YvLI8Gzfx8pRG6ZdLIHkIJsQVBKV6FIPRptiuqJx
EI6iigKYSzQ4jfMxwuB9erP9uvBQ0WvWZ7cWtDEKSQIJG1l2yVx/ykUTj2mszXn7obMumIdppLes
rgSOoR9K/0AlhDqHOrpHPhepFE6XlDlUOn4l9M4JdUPC0IJUgp9I2UoIDNRFsgVy2JApAZoQpPbr
WZpqeBCTVXa0S9zR+a/wLu8c8Px5PmopDqPuqAuBeNs5KUPCRW0unjVxrzuwV+xP53/lMZPNbNx7
BqEpHXpxFCoyLCE/XfTSxPwsMV6hOftu+Ay/wPBqsTblc8glvUV7Sr5sNg2FyfJcXxH4YKAVOdcU
iijI6zxHSFmJLzBrOXDMyz5XT+kuq41bHCIrXnyr8loQOycoifkJVi9h4Nx1MptTaTcMxiaBAbZM
fGAcL0BYd1quXZwgaFPCRd7czvKdHKxsJy8FMxNRXz1SnJpD+foSMLndEeeh9GipdvoBfN9/dXwM
xSTR7ObbNXJQ5Ntc7y8pfMFOzhznbj2tWHpLQwZC9tth+sJ6fQoAkB9KSGpVBVanPT5AGrFngeaU
wFUOO+bMThIkP5VxHFTYSmvvyO2G4UAPO2sZjkFH/UZroTEdr3+xS/erQ49nx0sdgHbmrUiB4LZZ
bYWybU9kgNTrLwPJrEmSSGRUKMEZfWSqDVSteBuD9tV6xflrPjlkaB/ORpQVUPHnjHOLSP01CxS/
z0Iqp/L4uxdq0glFY0CFZvfliPlFF6imhlxvuJu6QzMR67otm45PJBvAX7eHPCIxLTdTOAgTgTiy
S091YDQox0Al7lejLqtTCPsC4EzdedKdrxfDJTxF04cmYTkdo/eFv8mArFIf1qYRe+FXP9Jx9kkl
9QmtHSC8mjvnurT5AJfTHVr5IZcZ4fpgS2nAPGx7oepNP+UNdZ5PhNM8rzs6PO1jc1swliBmkNHZ
7zxMxVJw89dV73oJr5RyoxPUEHNC73Cv+6DJFYYbJYYHjr1U/cuh80jQ3Ifgrsd3gfU56AXIRjAw
yXLsiALyG+kYB6nrScx93BxRDzaL69oXAXmbK60p/nfp8PIEnZfb87YffYOwsuledNmAusbf2OGL
Mul6GFFQLOUmvYEetEWYM8+XM3FWHyu1KjQjrpLNvzOz9TxizDGf83U81l3WPt3sxffLhU+I0bKq
ijoiz8FodMAJ8ZacgWWVdi9XhrXUH2AWGnNOeGcxG5vsxwGuMHlkRXrBgfk3ITCDwbYloi+BrmG/
pXEEdcVOJqrbdEtbEhbOmMF1hxFS25AjTG9Um63owkUg6ZPiYyUyYD510wZBj80IbHiki6aNjZso
XFVIgIHC5dXvCQ3UHaLmdXGiXUwevI87KV9N00RMnrmOWvgxGa0ZDaxi2LxAZSKgzAiHyLzoyRA6
Nte5XwDYXjtqfbx5a/jdtr5KZEuzgSHdb25I19eQi9LI2PesJR6g4CdD8d7fR8yPj9Bu3S5+RGM/
d/NRv+PBvIL2wK/vhQG4QylnVoWuUm/+zD2ZvdJGzhe8197M0ZCbhVQL+jXNnPduLRa1dLOaUqRD
2qF9LLvIUivOYkqOfSjnH1I6SpuRRx+6Ks78dF82clzT7BwtPpgDrAbZSaWwjv3rhpDMUG/sf+t4
zu/LUk20lQDHkLxbEJxxrcf0w8TGZ6Zr/dn8Lku6aarBX1cgqL/In4fIlM6PTH0VMlWFDDAt47El
+YGz9jin+Vt3sgOXj+eWkjwkAqb90fpdHfld6MuREYOS51CWKqZwWia3h7VgQf97jli86QYSl8ue
VSfh5OW61an9ECM4LQrtf927FuPdEFEXeMzrHtl6KFVjnau9riDwzEb9IlR5sxDYsEDIhbyV84G7
IT17kYHXUM5O+gvYCO1biswYz/iIIOxNywyVJ7V8OAHin4DKVm2ts/dtBx1z8nUDxoWsJkNL0D88
mwfTEk6szSXKVvTF/kTpWCMCrlibO63XAJrifoJMgTvbfhL+a1LxkGnrMQNLErtPFtJWMEjmF76a
qBJyR82FmasVIF1Beg1tcBldS0k9hsuLLTZD7L4ZCHXMb83wNEfApt650VMUT7mbBSQnuDHqG11X
/EBbRIP9leQ7qKWGLM/ye28doDdeGBRwDpDvj/str9Ct1FniTnM8MRk7LHLALNIza4O7uDNDE8MN
tgFE06h3evOBGfkYrSi+e7add1aoOM/ULGYbGZN+L+BBXfDpnC95n/RgDrD+szqjzTT3aqhVzzra
rApbINKUWshrfCG1DkmSboL3Vvbo8dFUnjBQlZAbMvF0xdFNQNnrrfnXFXFwyKbTlVtCbSfCArJ6
5kjogoPRHliwWRw0Ro6P7MXkXR0FLAZXl6NvCgxrjWaksNDo8KjFcTTzPikXxzQYwdoTgwT074cA
En00UBAzFZhM2oOf+pN9M9xCM9B6KdvyKS7UE54E52boqhRT0I6dAPZn4l1tLBLZp8mm5/kXrFnY
fTAl6AMwi0dXPyCQDY8OK7yWNIa3h4tM3NuomOmo6dniHnYB0w+/ABgzdjcT3IgdDE8WUZM1D41k
xFzDJuELfwEe6R4WP1+sxTz5QKXtGxvoESzERGeXSgY34BbS1lmbldzSp1KyxWPHOQpw0/gQ+boi
MgIZBFKdmPoDQQWF8M+n1OFKWtMT/DxD7pGN5vP51RlvdB+oMS0VycDly/Ju27jUWW42Gfk+9wkn
BNthTfJ4ucKaxRW0uipwrR0XjUU3CsPHea3RoRr+MWwkfQSNmCyCsofYPvWCOfkLNP8z+ysHAkGF
9uOyJk3rr7BIWNKf7HyyeLbFn45dupnAoq0I/cD29jWAA6mF7UqeCQk4EGWK+eEZOEFJFdKvfzjt
kGncr+A9dBHAPo5DJTZ4pr75FGAf9a0jq+VQi+k3WBZ2r1Y2YRZT5aN3b8+MOD/l2zcIP984Y4TH
pOGEUSDOxGqR6VP9cNK+9Ioo2a0Pb4bBHzclNGp5rYQQ4gknas3dfGxCFc/d+T+7QlbVIILNYjYs
uH4zbdsoZxeqEGDOdVzBVel5nKBcptOHJpBst8dkol5u7xNSuoZDRwXKfm8B9X2L5f3iBMiZZOxF
13yX3UWuzGPPa08QVjdJ/XQFUwwNCIELdaYFp7ZQNfo53LSvqbK1PkcU0SdQFmwFCwJUczzfT+IX
0T8f9VFtfVkp8MaAczAX9aAdfG/074oV2sz6dbhZRpzoZwkpKrPgTbRCcZ5FiWMfdRhX6m1wR9/r
ballxSeAO8oU+Xta1ILofzBErkggaiom0gnw85DWVJSHbmUUp8vd4lSs7XeyQ5M34Fbw8ohDCU81
UCQ6DRm0kSxNiBswa9302VsEKrsiDKkX+yLuz068yx3YcWiWiRcJ4cCVvY26pgE11LLANHaAqIs+
EXjvBSKg0R0lbnaIEgTGJZMy5dO8BsK8nOuluB+emGKl+LlilfjUmVPjJTGschKuNzzSQoHVzob3
KiYI91U4oDsOvbTnLKMLaaP7o8rK/pyiorqt04Nggna9b9DYoCqae6Subuhj0C7nvrKHrdyP9zf5
sPRcemzhS18ovtTIGL7fgriEeISMiGKCRFZnJV+CxNaajSNeDKQosUwYqK6vokZltqjkTinTxRaQ
MPDMyA4aJHw0Iz8w8dwN+6IuCO9ii/YzmPXL828ItneHKhbrQGmkCDGaP9y0rooz0+J49Lon/3Ts
MwuN2Y5zPam/nwcUGNltppFO1Uc/U24MHd9M71fObJLaZLtw2JSu7RluGolm0vK4RmSCEicwQC76
957RYAw0luTGZ7bHabl+9qIQ3IPK+RKswetDWxvjk95JLVm2KWYgl7Ppi6qquLZthRazybjbgKiN
GF9HG4nydiBrzSD7DnRyPnW0k+Yb5laWMIIklHEU96lYWwPfv5eMoObAUeXCGh6iQ63wpA5qYk8Z
igUI9kg4If+tGsbQg0XLlNxWfsEwofzsdaFYkUJZfR8bJKKQrB5ESYD9Wj5qrCFEYKSk1B+OIz3/
jgA8t86Y14E7LldGeyNj8V1rqVykodpEHtM13oN9DXRRbAAiH35C5tr49I5McTbv5YzVNSgVTRfG
OebzMgawUoqK8vuDuWgDkJ/pJ13mygDmGpHLasfkuyUEjC28MihUpG59dRFGaRGbLbV06jeijsyV
wiExvbq//zGdlYpjXfxx4C92oskACw4vPRwiv8e4z5mfhLnHKl4QW5RTwOq8EOCAHVUfhB0kWON6
LdKKHldgzi/XQ0jKSeG4gKjWU2+L/KQfyF0BNUln8GaWYtF6ckqwV3izomwvv+t+z4iCyM2ivIdt
bUTeWU6jjnwj9CncMPiNQ7bLdn1Nhg7AFvn6uvERFDsFMex8K27w1srdutBs4cyyt+m+wtQzoTAR
jDX2SqupGljfJEbFKvOqCZ+IPW913YV3lBeuz1HMpzNzF1lb8A2o4aDo+oxp87yLpVE/tA7HfbyN
WzlauvSd56weFv5Gr+EK3XE96rQXA1HInAqm8s45pJ32Lr0yFBAd5NPoxQoszu8sTsDmB8r8Fouo
EXtAxGiE2quzm5OHYFWULaLoOlbUFY2o6mHpPfR1x0g/PA+wIVdEh9tfVZAMw+uXoENBlem/K275
VmOi/zmZdir01OBrnin8Cxkn7mbNwXtYDxLLhI6ypy3hMV8x6mGbOcVUCuWhCYEShGHlL2/foGTw
LhJ3wuO+WTnp8WEYXTL5IHFz2Or1O/r5+rEvcIiOigTgyq3LY7uTrRetkbsvsNJxLi2X1Vo/J1gj
d3o1/LxOoxv2gBNVefuHCLpp90HwKXSX9Rvisy63DO896rSu7ToXEJ9VpckgMCukzRZh1E4jJLsz
c3QyyIELd9V+m5LSsP9Vop/HLzu0yY6hF61ZUv5UDZQRBM+z6BFdk1Iz4THuPAG/1R8hUFWpqseb
qimWBKZLlrSpPUd8VA2rlpV5W5MwhTlx3+51H6xVztlR5kfqaGlaZHrdiCQcA+OQ+kaNtu35QbRy
jwCCT0i6YXZ9Z+pCg0jIY5yC0CDHwlovKwpiWeaqRxmFXR4fGjj8+UDmWXyhO9ux4uEe14xSoCyX
wmQmk3n/QnPaCMO1dH9zi1VEVo0mP2hIAEx+vx7JTR0ttCXg6ew/h60EYMTv2cSZC/8gOiK3seRe
UqTWoP8wVy/c5rLm+qzDAI5UWM7viVnVDeX0qy7Omrv4GJZ2frjbE+Kh5l3eg1oSvdDDOeHUWAJL
dCKhe/Fp215VBoU7sOGkvRpuUbRIR4++KLFLQ2YPYbpSXqDu8lRj3lnXdT5yaTuX19Zp+lQUa6Dr
Vmbb1HPbCd9ffaGUdit36i3uE1TPXWiFbNi3FDribvRDRm20K4XLc3N5cqkjwOrS4bVWRy19h8Sr
7eU1jk4ArjFNvYMA7NXKdFQX4ZgW2islojr5mIEIYvhyhJm2xxQOqd02e4WDf/DhDwgre1SoSyga
4YzrEuRi6BJPOv+z+m1tCOWGPHJMVX9akwr+deqCiwDcz4EADtcwAhCwK04dWG8gnLfojJKOUCtG
5iB3mBV1pqQMLYsyQVArFMz1IeeyKI8YI2HEcfdUzkAeSJ9P4hAqZudyMD2CLIOWvuFoI+/PW1VV
BXDOBuk1jbmVgZXAiihcWTgeCzRERh1yPsloF9Buz9IVjVflT0UViCtOMZA1bwag4WPMdzlXvyh8
C/cMdhKlx96wKIgoytgH2pT05dj3FqOZmHSfLoH8+yJtHn2/FQdlsvi/TimzF62/nJAQSMtM8nlT
416ibFshjro5+c6pUvCMQ6JRPWlflj6i9UgM6dKnKyl95wAoraqN9Stj1LjrrDsOhdb5T2h9Fxdv
egjjkOhsqCrTcLum/IxgjL5dyXJZiwAbtdREatKLtlqUv6/2SU79g/TcNOfYH7K4snnVLAMAaGdD
3XkbqG7A5bBNcDQjR9lDp+nQtKoljoiEOFayL5sP/15YRZIairYcJnmK/Tp7NSbGAQPtG9rPlPB2
N9Mns1ORIDoYZK1vOx7f4/8qvfcHMj/uLCh0ssus6YCqNDqiNc8KrYFKVaoe/JP/uKmzs5pKG5zu
/ReThgzGalJx9HtyN+xkmSjIQfuD/V+0X0wSv47bNswE188/0/Fae6aJpjR1RQhwM7v9L+Wi/Uch
woTMAr40emu1I0Qk5EKhCZF4iOvzPqfwjWI4/dLKA1Cd1IVvN3LtQKav+ZQ+0P/osWPIqfIO0OPJ
ttipI2OQhoXEh+OP/2F7FRGTwFF8f/96QUaYOcluxB7y5v0k6inmi4upznnfU8LupLt3gZkWxics
Dc7xwBgytoiDvGE1smBFSzgvtqXSz+mWJpwiH0SZNCt37c9B5RaI9w6kt4K3HbkMhUVSzBUCToAd
fEI6odjzd6nHgzD4wyA9ykvn/gZJqxYbHM7okOgs2i16qELSrljTw7CY+En4I5BM8adRlB2ScEcE
BKRW1UxMklRDe11FRksMrHpiMGF+0N53uwO/iAvBVkj6Mo4ZtNACObR9MSAsuoPfzW1bdQky7QBU
0m/N8E83v87H3cqBnPAGXyr1XkazuuI14q4Re1H2bqzZIQM7cnNhFhdjrr9mkJsiQJCLyJRBqNh8
IZGwZ3GJsyEhCxk5rlkrGDu43IPdiYHQ+hYebjkfJRncJZbWEdqSihyRNPMVqGb3UeiKebjvPSoR
SlVD2z8Ocp8LIAm/KRa38LeFJWEeddyMD0+Wy4WL1JnpRfWwnZFxqJuMVs20dAWWYCDIkbpB6UZL
J8IqRP9MtOlSVnrXFpPdsVL/y8nFTtG+qKOzMcjZFzf4o6pHSchaDT1d/soGAkB0mpgU5VjE0vhp
dVIU0MIreB8n2EE5LmjnHf4oqFTvBrs2CWdQFQSEaTdDmrpNHSJECAmsXteZXjeN0RWNpdw9VjSZ
zVChdOpFye/Y+Dd1rsyGr4wosh2okLLQUUz1Cn3l6gIV1J3M3AxoRpFjBmbU6KQhcOQ9JzTuAqGT
Sobyi46dqopH3p94eK69PwJ8a+t80A9pptEJ8HGQc8HtEIgOealoG6rECF6nUHGiP/Qctym32ToO
sJm9xnFuN5aspj4LuE9bgeRfTMdSzDW+HzazgfEM6xU/YjxmZdwnsqofxTJdnYbmD1OA64cF8J4o
zFJatHwvoZJDyMNOSlVINii2BxhllZvA8PmUMAKuHWQqVfA+H4S3mciM7EpriKIzSwiKOBdz/6LQ
VMZ7zs1C5zo9Sxihu0LRHW8PUNtunyM2xEUX5NhsDrrES7J8rX2uYpoIC4TwlzlB/rC5Rvx+4cAj
mFc8lk1WmbrNdzrPo8jHeQRfybADj7ShjCJCNSUE3vDOCIy8+co+0RhUhqKiv2YZ26orIx/mkacR
RXt6It7LDfegBPsHlJrTVuPjSlQ8nIrc5VKMfkA/kRYx3mwoRWW6+0B76AsXJE49Cq7tW/Fjhhdj
v2sGg653/rU1u+Ev6TBzHPGe+yBHcD0C7Ci9W2Bvb0vqAnvO3iVcEoEviewmubsLWw8TgWqhfC6U
Rv+fDL/+yIg4kwY3yo7sm7eNoPo4Kmvv2EpHAOElLIxOndqoNldYvkY6HRGjOcC03L0dKJZhhpJW
koDDDu3eifRm1GCv6gkJpa56cr74gZZPJf0mxQhge46wBOIx/dxPT+6QEloEQX/QvDkCiTBqqztJ
/jP6FvIaym+pYjskMZGDiEbYvj4niH9LmIRAHJ5rJvJMJ37GTMZO8k6PlSGhoObJ4kq0goVLhPeu
2waGS5ECEUnyXidjtgP7B3L5iUL4uEOVAZ8Llnbm+NAUtA9gesQEWyNpNnNMosHdq6cEy6XL6xR+
GuXaFoJhBP02AEqH/ZrbOTrwfRd/Ygj0LFKmoeIYtCr7aUMd7I+aLSj9mlBqi4osciPy563uLzCi
qwOseIpxiavk/kkqMPuXqRL4NfyeusMRo0et+RlHsQpQQHAHjySM1MJdDCWkFxvcSh/GHpZrB6zu
NLgzetjssH4+mwfEQ2gdvcOIM1LdxlNWNDwm1v0z4FBl3tngN6v8lmJncSxzpBCVHcNnNVeXHIu3
tbf01JOZwF6cE0PrHg151KVut0CzU+Bm/StPe/fhK+Pa78SYlmXGF4A89D8nQEU5db9wWmbCOV2d
8PDZUjRSHrFLFg4qpH9aOwUbspUhkp2VLRY6FdX1zpV75E3Uq4hWKMFHTsfbjfYjzegHEmHZ7m9x
AD78CTP65x71G6OBE9tW4ZCcjIeJ9xPLF6c3YZS3EPKkGyekRFx9bhnl2WlFj6n+MUk5sq0oVxMb
QjkzJPSf3cbgT2Z9kndgOt/RZcIlGyQyHD+u/4cSBVNEaxzcPqGZQih0vHfwxKsKwo5HqrD7BZ3H
bB2E2i8NZpGxxnuS+qitdz6tXZDW7XC4v2vQVaCPGOHHUn171KHZlJuTTLBmV3AM89IBHA1pZPf4
FCpoiBqH2Yf7Hicskxm/Icm6rUowKBmgwtaawNqnZy1BZdWUMyofnZBMKlTBOU0K1pYuktra3/8U
phStQkeioCaFW7wCakVv1GjCNYMM7exfyY/v+NQhuN7zlPH61WYHgt/zGIwQIDYlh4j78XN7VU7s
NrAsvCJNBssTnj5Je4iW0dcHQVesXG/HZsKYsAv4QbyeQByZOq1Fgst2Wi/HvDVCkdggCMx4Y5gg
Irl22+IAuSp8iBxgN0Mj6x8Z4ZvROjuZ21Jcmezl5JG+CIIy5uTaMNXFSXbh/qInn9ArTpwasofw
K6oS19evjIZi9zdSjZ4z/DqqCA6EQNtiarxjKtQnMOPGYcnURSUB7xIZbT9gdPxvxCZZCOFsuv0w
Aj6VYxteTq9m4dxLqGCLFqanKZdnoteqIHZY2QxD+oclxlXX8qe02XdMAp8CrT1TTbKfry63YPlZ
RVIUUp00ZK02aaFqpBK/WVKOTgpKZaFmfdiknV1Xf3VlkYADb6cCl7V1NhA2x4o7nCDtQCaswT6d
rPogXCYFF92YQNQX+F7euIUl19c+1qv9PJCfxrv+ISa7VXAsZDlBMXLAXFwWi0kRzLH49JBxqEnz
gKbE/+7wMw8obG1YfHW2sNa/cpB+l5JVHLhbGGtnKjb1jcV5icWPVetTqVnFCyVobbC19UfbNros
r5p0gERpVM7fem+NOpI/QVyet9Nn3VZpVtP2kdugefoSTHsX/XRkJ9+n1WId67HfLspODDrFiGwU
aqHPZzkLVoDfsrEZWvQMI5+MM+uaYxYp2y10BeeBYQMX4sPe6zi5Qn5XqlFs39aY84Tukwn1LpXw
mD0ws0mKFZaRow07B/DPiZjW7qxRcxQkbDcKjhLo8D+CtI5/+boaeMNNsIKYhvd9mT+xfdMjna4Z
SPjZnf35JtSpsWy9ZBRaRJ+dDVpBmApIIKgToCYb5gguorFPVNfxJPi8MvwDwhWFHF82KS97UL1p
3g/H9xLCUUbPVokTLyD8o5cluA8sWMRPRQT7twEPL7BoZI8dPnHhfLN1aCA+k9reBkVOGs9gcnVI
O0OzM6Z2VxOK7miFglZZ5ZAykwNzCgNAdMQFllNDPw2Iv9KCs/LOq8TODEhnH+Wvg40Kr/lUeOM2
FUoTmIehlplV/noJbGbKpbWVAEPgAee3rPWOw+2Isk4IIyDfdfjXqRIPKfaSmqqKIr9CgLIMt6Ca
NtQX2W/N0h3tQA7s4t1x06D0Ca3zKjpaHfHbZr+P/+CxB19kCxpnOlx4gnKDNcCIDJ8k5sfpjxUC
gLZS9U5LBUEmj8YZqAmLm/oxLsvo+j4CmObCfxXT4uG7bIeYggtxP3RAg+YNHqPPmeAF1IejIpiX
cw8lGjJOvsuOzV5x9sy+hpL/rQSci2M66FcThe0DAQRkc/EhxvOWYJxf9D+b1Qj56M2bubeSyjax
fHakOAPKmA9u6dn16W9YXSFifr1hB4ahOwcRRS5DzX1UAg2MJEVF+00XpW95ZV5c74VUlEPeU9nI
nLCEpUiu9ZzP60vyMA45dqh+Z0BkrwkOjS24GW6BJO04MOEzhMILnGCyEEgpuJbanuAvkclKjG1G
jroB9L9dX1J0K0LEx5rrxwjJKKyy67V2Td8rJQEdC72Sr0MQf2z4R1c2S7vWjeVKDVBDUU3bfgXA
rfzvQGzTM1PUJkpoO2sEtg8zXLWW0dwQmgdcIe1EU7uNjLBlEDBIvxLzv7fs0S+92x6Vnf8VIl2v
zvb4P34Ly3UV89VREepHB40hhzokQo8ed1J3nv29Xh+IAypzB+QCwjXduoDezQMroWSfGqLzc3Ro
iTpkiP2i8PTSz+DJNfKyAkyQvyHYDFSZ95/Jk6DEhH6x78Ompq9SF3kOZu8f32YteK6qrxNX7y/P
M0ucu9NdmXPwEFtEfanyJN0bs6B5s8sVr7z2hOCMKTUWqt/wV1k5HJGt269i2K3M1kb6oNoI4+bz
RCN6djQHy+z2W0oKr+TpgHVThp7flVRpedVZSe7YBiy/v3oKLMTOpUwNkKy3QGm0o81S14jBGYvc
h/14Y3nRLYEz5DhpjT1j94+/CSH1L+uNxRoNOr+JQDPRHWm55QO4B2wjXPEUDnWOchlgYaast6gw
jUOSjINttrr+mJ0HHeJAurh8+hXvXfIZbZP0i9N21H1E6ALTGXYUZy9TclfCTxQI8/0YIu9xO1ln
CEGOPMYUe5xm+i90eTvKUvgRkXOZ4A7qOoGm+tSGKI8AB4QYlFdJ9NC1TZyrnR3KDUguQkQttnro
e+Wp4MDVKJhmk9vGkZqjSW2gVSStBhX6cvQ5pBNlU/jzGy73gdHGaSZk+oWwMZ2CYxuvVohArEJu
SFT+a2MWc2Ad9OxKmQP6MJsU2ObEf4kIZ6ZRDFiSMcoRT8JosgjggCAVYBF7hp3ZoJaxWcPkedRI
uuhyMHcp/qlP0fBVnxNHLQ44iKasR9iTtrVb9WWEzbXtDaLgg6fYh7/7bNI1ibHSxKh//wZugOSn
rgRghQ9mYHXDYT6xTIp0CA8cTKCWzgVh4RJ1EW0lJRhwlqK0HD9aw88nHrDf4ZyiSEFeDxnF97yt
nSTm/flS1bhUzg5m5T2ShiJGoYPeru4+JAWW7g1AyigBevZNbi11xWAmml6HLXpuyKVVsJawFyZu
yUcuL2muBsDYUVYI5qSh4QzxBrcaW3Q1gEDjbZrPSXV5UHCLYvw46Kdd8IJPa3Q9yaTMeo0n6WZy
X5ucJWKVYvd0iLFvdNA6ZMqtQNR2EdywIQ6Z39vkJZCpN67Im7mGUn4jwJlpXGEHZvmSvf/yCERw
HJQlkqcerLICBwVplo61Yay77hdF9XSS4vhmJWe6dzjKsT763zI6oTv0uu+EBFcCnEAIBDgzBBzY
sNKCS4AVYCHWJ1Y+TgmYvM2sygNUXrjbDMG6JJotiFS5DWhNCABDP5sN8oCDXQ57X5RvmP4SxVWB
Vqk1Mu07jM5n6ScjJoWRztpKbkVz7+K1+nYidJMsdCOfNb788ZZckOGncM/1/kIeGY3V2kE+pEZI
p2Vd2WqLZWhksSXQc5Sjvs0dHODNtI90DfxZwS2RxO+RY+Y2AW+K4CJVUUBvcx6yBZE4sjESw6x4
waGmabPRPYhhf4CXVmfuY6tW2gU7fGvysrlp1DZH34OpbzJsoGZ43/2D62+lYPI4pgue6hSKO80d
QrWFU3IzZ0FYrvW3qo6K97Al+H2J2s3WX75gjC7goBZJISM2aAQU4VOjGt/v2PWYE4ukPgK9l0y0
7YTwTrutOkizSB+iIJNX9NpcFzRWZ2byNwgrJD+oRrFrKkteV5cU34TCyoYJTzlM0zl2T6DWWYVS
Y0o8jXG/Kr6bs7bs9ySmH6WUS9mcZ39xssyhnmFlp3KyMOrSuH+rs4B3HlbzwjdxwnQI/qzC7pP7
VMDe1o6vIAA37w67TrzSihxeW2G4FNkxvg1w+pqdR/jUVBllxDI57dgHh0LdjRO5U4VGvljIGjQh
TcFgvrLF8SHbTaIMCCHkHBMdX2auR0rtDDGMSmaJuhqEV9Bhgk3hT0jeagfLM/OlGwNIJgAx0gM0
PpJK70gpQ3b/7Ag1i0OlFo0Ur0Yqqah52ajUCzPZXg4HsN5FnZmqAoA2ACytwSYaVg+FpaVXeBOj
irzsa+Be6W5uALJdaXAKWGS0mIifIU8/ZwOQO3IZb67uuJiLVHpTUjoIuT7smQBc48VNPpRj1uGy
u0pZ5sHFQPIqC+YaRT0iihxKbFliaVlzAscU1B55UTPvXk0Bt5+Q+GUuYddZK+mbx10xd3tlyyF+
bisYyHRxYiFm+8uZOA6dy83CzosHml5Fam/mZUiPupqalgrTqLSch8YNjzZUqZCS7N96QDP5ixUW
VYagVybmo6dikEDhIeG4/AVEcKX3SXOnohd6eXfP0udWHGDSpXC9eY3mj5zb5DbbXnRD6g4SRyQ2
YGM0/ImYlN70zCiSNVnbzMecgESbFkWa2mgFvPh3ZZdmAZQy2Wwu8Bee+a/5WzWlQK4ylAIk9DNJ
puPXsKP/6PjYlCG7+vheA4ca24ZMPaOvSDinpUj8CumQIY6RKyJZzrzJcEN8U9Ysn7gB0fNcF9TE
4k3XwcOULk38dcTF4IZ95I2lXRpm4gHIFCCXArIUU+q10fDijfwF6PpeSWsOBpm+vztHhIoY77ke
4naa1CrFZV7aNHQJ8WUy0pw0tGsxq0aG5dLltv9vc/nqCAZfwE7FBgQ7+MCNJscZ034On5cVlMo/
RK/e8KRr4BF6XIR2tJsYCveFUe8Lb/uAFwdC3ciGiO4E44Vn6cXubmI008kpVUZIVbtD9OxkJ7C7
D1i81LqpQ8xUd30k1EYMlVxxEQpUNCz/YXuaz4KCA26GA+TRYZqhBErJbUfhVjCYaMOYuQ4mjy1R
vnn6axvHJgUpMvEDOyucw08333okb+p1ZioE0OPFKno7JGQlvh8h9ybCDztqwKMl9PcfPRuIWo4l
DpP1yGkMH25X7AwpLKE22wEdtwIcMbnseXRtseCic18ONzWpHl514EmUjhpjAQm9FwNNwHPicYAW
SMVjYzyjuaj5klSjBxqKkv9vSH+h8pZ7aQeIJ/pGFHKgFw0Lr+L3yNV8a4r0eF7Of3vk6BcHitAN
YrP/H1K6SiHQ6cUpeA6QbCI5qDKYvn49Y4Vc2NPtFY+d/qhrpApCRXXLpktMSHnyCL7LrIRjEuGJ
zr/VwHi82Tp5f453oDAG/3a4TzuyzxECOY4hFcRwmi3g4HYw8rWqAzmX8JV/WRjpMpWbt16aKGH9
xcHz102Atn6gPm4uiYZcxlbJeT4HbCuX+77Ns7d9T2zq4FI5jXHl6YZsjuZ4rYyIW63m68WTkIVP
/eNUaSqpa7BBUVh7wGSYQTteIShAqv8ENd7IiNH/lhh9RCxxP/7JmphVG3wSaX4tBCnJ1CQA2MaE
Q+30cNWSoHToTWp4jU2k/o398BehjDw+6wDpspil8KXELKxmoZMqE9aE3UMBm4DNjex9/GmaJceD
ojhHXB5bWuOqKYvKskwLKnnDmg58x5Ppiec7rlcwUmZ4J9ySkWqq+IV9LlmZJjngBnAIvS5XlpeK
UtcUu25+Rn83sOsDGHuraO7wqqtjvEDQZpeeez/hVEU5m2KdrHAYSLTFTXx4BiwZJiCf9Ql3YMwV
rvMOtDaoiA1VxAqH9XDeSJo3X5RtxGBEAxjmWwZKKK2HeKEYIo3k36O8a3fOOThW3gcXdNHVyzkD
cXojK/GHlCWnsz/wIe4GErq1k4MZ6BGtFUJqwQxNSHYyPaszL8fEQiYd8wQ+IlkcFVxYS4h7h7eL
4eWUoG4CYYtnHbiyzU5fuMVv66M+0tQ+GG3DIw2zXFd0nW8i1II1MglUCBpvZp5OQgtw5QQvnbCS
2hOXleVqvRa8t0CCBxGaF/v0GuilXQyGzCFHmnioxJknTV5H3UxnuGnmsPk/Fzbx4jR/sFakiVqo
bDMvImT0GfgCRjM4y7yx1gwhEpILtXzHjtmX+ulICIEfvs+SRI7b/FnqLkDNSw7qJwM4/sdBRzlr
hm4GLPPJ/LayqNNUmRYe0DAenoh5J6b+BdtrcYN9Yp+hoHMh5vFAp0/WatP3Jq+CCo+hsrye11qk
Cwxf7I7hoQ9qmk8MzpbB1H9mJph+jLv2zx/fvGZNCUu4A6fpR0W43UC+oQy8vVOxeJE11eD5RLuq
H+ozOY+rbC+19QIqSxRAY/9HN5f6n5f1qxLeDiSWZFQijoDs49QwdhcprvX6Mg0NICI4LljUcDPE
f+tT1ikj1/7LMOopXAEQ5orlCeAWGIAm2JrJnGSxoZJ+Z+PzwcHlXbCpQNyPGyEp6qJBQwycmDYq
VpQqLGjVifjC82AdwYQ69kF8lhMKErlmPKtSwHpyJ0djbJ7sJom4xfNU0HTmrfNiygLoieSw7+ay
nt/FXz6fmVAkWwyqfh5ZijmtaOuGgIgs9th1jgtZKZgAQGM/9qVNlT04gZNwj3XgSVlbvf7KtR53
A+yHKVJ9tba8Zaaf/+VmN/OT/2qHEA174X0RYrQIM6qy0MahubCM2H/7/69QeN0ncLMaTty5QzsF
yprZXexam/sXqsnWhqPm18dc4AIVK3x2kHDSb8ots9CmGLqpxNgOvVIoTGxlGEetJz9QQLSPWgH/
kllyyFl6sOAtVIFTB2auWsItOmlYplcCfA2p5cN/dRcN2EH+uBrGTm4yEQ8j4ewd7x4R9Z/+ZSUz
Aqbk174IJ0D47Ce14MS8b+lAu0O4BjTwsF4nO91fLu2A9c/aFhM9OV51B+OFec9Rmcp/IBXz8XUo
rEg4gF+DHzQjPg+R+yFnl3ElCYo4ty9NYxh+/kvtF7PJgt4o/o0dSM8Y4vZKHAs7eLUFawoQdCJO
ZiSFrFTDsTTq+kpHvibugoqJd+X0lCzi0rhQ2O92WkvJaOyQdqSpC3BgU2v2f5TFytBFIJ3FwHDy
HCIE/aKbo5YBsGErNP1sSHArf7ou8D9VrJM5ESKbLRbBYLlf8FOCPRjZVXIckLySnOzCOigk3DH1
2S1HKeqAjivHQp0J3MhfifQQnQPDQDz6/XzGlwT2SpmSDEbQjisAGXwx9Uxq/N+ob6KWOnIQQ4SP
v5EKS4/527rCF4wimlfxoOtsAyy1yLvqsgdwpTmhOoKZu61mtr+qmSx/urLMsk1LofTG5I4OEZ2G
CE5dVlsI8qjzjSVeY4io0OO02dFW3H6cn1BSa09qKfFHedITK1eQIl9T74sj8tq+SG1wKOpZDUy7
9Apb8oWaxo0ZywijmuqvAEqPkT9dZ336UwuUHpOuus8gSQoZUJXeHbEf44J7rm0C4hkeyR+2b4AE
oyk3b3FWa99aOrfEjRfJzsfZtSVpRThO85DKol/Gd5bHCBFSJWaF0NuM22AFuABNfGeAfCvmdmBz
WQtL2RbUH8cEBahQndC8eiLzlqN/5dEXMDRdGOYE9Q6K4C8fcR/azazDhWh8OtGsU+WkRM2FWy/7
zQiP105ixyiy0HRls6v+gIZ4L2Iw9U5MRkunPzUtWoAT+TorBP4VjFk/tIlqxANSP6x8gkmbx/3u
hA306sNeTzuWfTApNoalag0BrE5SaMsHSqnqKeuNjBazeLpFEdUQOJDsoK/CJ20zgcReNahAytJW
GU76wCsBacv7qEVBPmXhGHhiJIvDdfejVtfr2xerzhEbHuOQG0FB1j5SOcefUKeCRsIlSEXf/Z9r
Zi/yI9DE7Ec0crbkvPAbe/eMzq2yVVoG4W/yDihyRCTZ0gxuAM1kd2I6FZwduhp7hyHcqrJA5Ovw
+u2XiyTAUKSkvzZ6tvBa9GcV4AFCTuXlVXy/YWvbctJ3n9ewEiPt3d+Efj6dwylwrRmkBROdTbbP
uaCstSSR5zl62QXg6GpDr58uvADE/TkBzTsJDvLDyVjcDUQOv8e/Ycf76/jFkcs/7Gog/M2p2Kmi
RVGqq94hiSiKTLDDljRhjusxdVAZo73zaiZMswi9qyYuWjofFmReMRURrI8KMxKnfwTMbOXgIPlV
uxEIUExzTNYgAjA/bgiOsNfYx7aLbv1TkuVeuPlHK0WE7rFzwyKeIOPhfU7lfc90oUPchRXRjbDe
cxZIlwZ5pVUkt+g3ZrrvrMUFtMw7qFb22xcq4JDX95sklBVumcSBHZdivnPM0T+WsBYw2Gkxvdz7
qy23a6V3WclX3frWkyRLRBeKI+/0zOYwO5NRJ0RiSbv8X9i0tOS0a1uQqQ30c60SoLR88fU5827Y
QnsZFrQTJ5kuwQ+qem+z7uogyK8j8VEvujRCWwRfqF4YnjWHSdVTda6Qdmtuz8qnMz89fbu9AczG
sxs40YhuTnX6ZjXCqPe9kLavm9E5QxC87cSEilRoNmvnmoc7onkOG+HRCDoVPEVvjtqovpvxGXdJ
gQ0UWDE28hc6kn7vFvHI3Bihbu0iqzdm9LxwGdCq+g8qsK52wLxo333IWHBMRYQMy5/GXrDHZ2P/
hztTRe3uqos7msGlCbfqicrYNhCcxN2fHUZw96AWnueq97gjIgo2+Sw9tinIbAUVn61lhLr39DYi
Zgw48cSmRvzONpWDDNBKnUNrJ8KQIRx1g3RrBVTpGIVOKrKgMnMibw0mF/x6C481+4VchggBYy1B
YJoRX3Cd1LsslFWALV0Br/3RjlomiSyDIfBn1naqas3C38WkyyfDBlgB+R1UpuB6qsHC9EAo8RGm
jtiNfpWv0BuVRrjLqMDKyjOdU1rlF7s7pj+z3Z4IWbRlelB2NQL/v4Sjjy6nX39dkAB+Ltgn1OLs
oOjqf/aghcvWTGXEgZUjkxEgiSPgD6CPqNRt3i8MPTiMyAIFrqVIbLFJ4wIKdFLF+UkyRuE/jkYz
jNFe4NWhZBERPBvfnJrVvIyVhK/QJEwclFRiV8lQEPjBUUFfojQWOos9rmanLEasBWLrciSflBwC
3O9k3KhME9mJVl6JpE/iHha8mKW1Cj0qKvAQJNNGKw+CeFok7rKjlTtC0mX0zX8CoLmLERiksiSY
eKpug6AKezaVltXkGx/qYjzElHGWdy5oF1oLznq13flTdx1ecz4lxaqo9ULeEUYYW/tpqBxcldDc
OKENG+9Fi2uXOIYWSM/HBxpyUxCvoU5O+vuGZVEjCSeKRgGrZ2SyirJKPlJjZwROTuie9cXrUSeP
hWHk/xh1gqbuBHr7Ehds7d8mBhyy6DnsTxDRtnmEwLtpiwmK/z0nfBfN2Rbl3bGCuFjweGcIsySv
oV80DH6KH0L9b5VzUojrAeCqGRaOAA7bJsxeKQKM0HKXSC7FrhZ9oP9uD86msHv1ynnu9bA9jFw6
n2t2YDEvQDWIg72F55nYg9OP+4EtbeATsEZwMXIOtAvGbi1GeMGP3nxr27KF2vD+7ZQC5j+7dWZA
P7WQu3HEt3jfYnQ8KZXfN0Fs6Z4i6IEggDYm1/g4nHYZNGLbfop8/PQumoBPtKdY0vGDfJqMTUgQ
e2bouOL0ShrI1Jk5AMbFzNlkJL+MzS1r2fMxJj/B8p8c5RF2w2KUtjkNsb4dFdrvU0UrUyW4bYm/
tNebk9lnzu1Puu2+/ckFBXKr7ZZzvPADzMu3sH9VkorE6s+I/WsS/l2X3jOT3Mp6G577V++ApnR6
sUXxd4753OE7CaEprVKNdIj0lxHrxvV+W/Y84lB+adQ707scgZRNF336leA8QaBAuFynVJOsdYbz
mnf2n6XqIsSI51BFSFyLXoZvl9hlw8802gkLUYI/Sz2JaIbP5fCdu5A2chUU/PYqPOEKM+Q7GsMu
oVQ5P/KPCaSkOugDjNRfLxLytG/gnkPPqB8AyR8YABuH5qa1TivPaFvevz5L+2FfSFyIRfnnvQ7V
alNNMM3tzXEiDXS4o6NfFFgxW9VY7c3l46CYyrWRNadzIOcsW6B0S+dIM7zY3/3zS9hXB6Zjpe5P
uh6IGB9OgeWDK83tsdg8TiTeVWUYkc2iZ+DrLNt/YUmv1DlitZNQ+E+0rvgEIdtvMFVFQAF0VDtS
/EtJPuzH/IfnlUUXj0ew36GhnXf60nVAK3P913QhD0xuwfqq7aZTLyFeh+aK1b8StMtJeDUYZpDW
aGMHxadqHYo959NFmGq/Ivwi6snkracvjwqkmYcN0fyDVKiqTjoxbKYQaN8qwVPh6FpYQYGlhCU3
g7h8y4x/KBMsQDF7xL6MqoLsrGI1iNkuSDMZHRUpKHP+0LUTFKBj545owzd4oMir1HQkL8rmqeTa
XOjoYatKPaYNCyN41zurpZdxkAHGbDooj3JuPW1QkisqAicNlUTQI2l0dXxtj96P2wcLAEuJbjR8
CtHThAhCeSCiqJz8hcO8aLyuq3rsfv86tsoljTjTQtPkmj19l0NTrO+LOw66pP/NhdJYPGwF7ifR
EKJrq/XK0jUd2v7Km3d9+mMiKJh2TyV2GvZHnFAYOh/mpLe3LyxJ5t0PlgYtDRAQEd7IZiTiu4CB
9a+beKr2fZEL/AQ3M2rH8malNWngdQvMMKe+RUOjH0MozgV5JT67JuVeBjpxroMPOBaPXXFQx0AY
lFI3pTbHa1xHvXMNws1rYVPpJDb/5BjCQVFP3JEPal+DPzmVWv4xykMMOtHenAIIWttwD2caNY1a
HCn49N7bKMqbUItG8hTQiX0lnqBbxj74tM0n8JqupqNO31u/mVF0Z4+ZG1oYcFb3CyJhCKDm8J2Z
LIE9YbteqHAPKcNvyyYdcmopPShaDU1d3hDRfcyy9kjE/Gtw5llUP2nqRyx7sYoUUtkseH+uU322
1JFEBgsw2DrwHUh2b1CPwa7FwbbZEyFkIWHQqQ/zPTWkbhqP7tgsNVFMUaRNPzhBhwPGggEa6/kG
yP1Djx8HFEeWZNSmPnRdkqhHY1ybM6rOZot8lWX2EeOpmrP7gSBy3enekLhCO7qK6mEG0vzFc1xa
/8WD4xcl5Xnkqa8mzB7ccwBw6o3UtxQliF2LRaF893ASYv85Q3pB03ZURTaVRMm4aJd4Iw7eiqna
oRUkCC1u8CjVG8qiNK0qK3wp4uCxBhMQDksYBs3FPiJ+ZuSoqNXjpqmkop71aZtlSu3KDvFr1K72
z0alLtBz7W8UOFgZZZLz5osult6y5bp5Y4ltkGjreakO2UbFOfhJQ+K9An1X/IshYucO2KywWV2Q
8t41ORfCLwyDoOpkcp4jIWcm7LIJjnL1y0kdw/bbi6X1y1KxtNEu1DnLQ0WzzM5InPX0jsY339gU
hmpLuNfnnJaRP4aHFJndPBNU0t5sUHZgR6dlVYr8wAtUV/YhnvcQbc4OcxX17POooltuOh2/nmoA
E9q15lyrGRC0rpUGgV/1WrNtD7qIgwO323S04MkJvrCRmwUpIm8qJJhom7bNMMAkESRpgUf8hN7j
FkQtUA/uK1xOo/6+mSN6AqHBIeqFDeaHPXCRTYawlYd8bc7hAHvjQ0nzxYYcn/FW72ECT4nK2Etv
ygQ03l2iAwfpm2JyETG+u6hdIRfcD+VlHzqnrVXDAqjsAZK/G5aYCkaVc+ykHw32ARunekiSsT72
wvYME4eXGmxfOb0NAVBEEvX8OH3C9lxW+dmAIHSKqm5Of2b6L4Kzrb2m/Msi6ZT/dmPE1mwfu9jA
M/6+D9eyAa4sgL5+igiv/w6RGFBSk3vqXbPzKNZYF5mW5Wuq5iCs/RPUXpF/cyPuKTF1ooN8cfrU
5u0sAHSyuPQZL6CliVQ14uE3wiW8k+OLACE7KjC2qPEXzi676FmFLo3H1o6Rtj14hhdKLEV5L6Ri
AVq5vjCLANeDe1q7ReMSLzHuzyU+kGWgoUnhY3tHs1P1wl+MnreBFTm4BKDPdz201O2Qy2jchhvj
UbQ/3fPnvHKjlzEWm5N12Q2kzITspL3WFMfYHhle8KP5dJlzRRFJwQnE8MpgUZAOFJeZUl9L8e3r
d2dn/xjHPkAcru6cMxfOaStkEgM22/BSPtepEMILPvGeyuCYPY4ma9AHenN2vvupLuzEDl6S9Cnz
r1DQMf4kruY7tJQBlCXrUjpNBpKxuNYZrgZEPm9xjnMgn+jOeMgxbeMSl5x/8EQHvwELfVjXz6OE
uEGe4ju/zMFXs2uHIAEVeCZ0bE5jPV9TaSd8tSN80jDTf6TEbQIpdKDUMDiOA9iC0U4K6af26X1Q
rLzL53rn1B3k8K1hCpXayLzwFfeY20Ea0yrC24+TE4XB9zZcR1Mu/j1xukLdcw9NO3qP29Q7M0nS
nv6dqzY4sPWaEA8K7GiAmoFaNAOl0raYad4OAD6/4Bf9iWP2H7Jv8/clWkFl9DFA090KqmxoBr1c
ebPDfxsXv+Vz1R/DCobPwxLzNdgraYFp3f6J9PjGKxjkutignMjHpyycGQI4LaSYgNlmc65CFEKl
18GP2o2C6ueCMpIr2NdxMP4swNpyjr+ome+2kMpuEDJoyToCjaFvjZZFi2Bp3xcaZKXuB2/DhreY
YyNBgfOSWfBkfOHENoNqBWGROzZMvmTPYDn12TMMilo6t8a2kqSB4kHFo6uKsQg9sdr1tcZ7bpGU
ZWxSZ0pZlD4ZTafEQ7V18KGl8GDuVthleiBx2NiDjPEGliSNoHiL4uJzfi/eSAM4w/yAky6Jmprf
wPdcxt0hlBwNDcxEz4smJW05ZiANz6C+NH6nqhvcvUNvC05nD6kuAhbwLuPkc3j1evnNDcNUO0QS
2v2baVM0NdQWBTbMIqOX1orkn3YEKzKgPh2aiMPazEyK32scTPzcbsSaWM1wT5Frfz8M3Xe/y+wa
v4lbJBz2gnPK4QmZ5TICk2F+ikSJie3DvqKgT4HBP07Hh8Hx10RRPB2XM66nHUqLolfEcN7+awmm
ZZNut1seiWxSP7CCj0AZTj16VVPDt1tHp0CuLKU7EamqKQxCvOjLe2WjXtNGaGvKvFK5Un+phnCi
QqZ8HV2ZB6Oh5IV7Myns/zMhZfuPibThcG4iFyUT/Ue77FBSN1WV+H904Ni4izzrj71ZesxIGd7o
cVG+eqHsy67E1d5MpqWz7DE9MvrTN0XmkEt7ecfNcZq0gnfLsnnSA6St5zNf+zrybOjD9CuGdkwx
EYz/tvC2hY9ycIFGYRLtCywESd9jCIOoAisJ5rSFwUZSYrWZcFAalGzL14mXwDMj2W2CuP4XAKdY
8Wc+2jEMSXYWtoAp4zcPyDgbq//IvPzcUByaKg9/wxHju4MhaB5DXLWhuwmaoB4KQZsbbctv+CRF
/YIi/RITUlNPb8GBdLzhhty0BtNp3p9U62oSo1Z+KqhsuUzQPGIW1QSzcf0/0KmC3vgr7Q4ljG82
wGmAkY/F05mttxyC439eBnKdWNOKmo6yZrIzqwaEUMo2S8qaB/cwADUZk5ewN3qe/ibFViRdDa5n
DZ7L4MgDVf1Hxb0PSYCR0NS6FLf/EtkK5/jO4Jsx22nbssqyDGlC3pm6L70ODHB9Ft9jTMumssvE
5yfQABqLri/6BUQFo7F2sey9p7YW5fZ0Au40vxhticdpW/whU+jWNc/ZsYPICoEeMB2hiD94jf61
XWl0eUMHIPHATtSS9PLLBz+DwSLf9WrVjjpXwWS9zuDFg/AbKFrDO84WQerUpdILBEUZDhVn8h8b
ijXuCNlvyS4UWLPbBTE06CcLGDimXpnxYOWLyfyO2s7yXMD2IJXeeWaZhbO3baDdXh6yA1stl9O8
a9Y8+06+j4hU7jC07Hj7I68bANlXbF3GpzlNSYSwauQbWMov3dQ+OU7KwttwAUO8oB40bZ/dRiXX
LSaZT7YxpkqCDPVyl+RtqPk9KYTYX2OQxsT8ycrF0rzwrRELViSstMePEMFJGLDFDPWmHDKo25AC
3FT4NRBe2PpQwDC8blgPNGNzAzvGwfKk3dZb5snsAbbdLY3qc/k8wSt7idZAp3TUueMsdZ0d7UkO
8Uj0xJ7S7d2DdvYODegdZoz7oA33fi7wAJUIIAuHxN4TMx4zd/2Fl1Qf94vfWeZCZkvVypUb2bXK
tJqA79qbEtIDSbLjPrCYbF0q2lZ3dPAIGjnYXVFN8t/3ztzF/Xedik7MqWZkz+aDc6FaYFicxy+g
ljrWM22dzsjrV/7pdmCKeqddOPgWTc2r4WcAd+mWxeU6lzKXswJYQvvJjSl/cyjxsUE/5UZHC8a5
sXXRURc909KBakLfpRNyr1XqvTvlB5PFjFJNi8zh/MTc03kEdVmAFToREOiLsPjpaKOI+7xAU0wc
FMD36y4xHZpecy5gRhLoF89m1on5mTzcJ1eETqnghvmXs0naQgLYyz5A7yGVQKBQbMGjZWEOxKSj
iuxsDT1+if8vZEqiRI747xxl1FivWp8vFmtSxDfrdYy4A8l1eUABRHt1cDqR0FbbwEe0xAfpaSqv
BPrppME2CosS6xi6CDivS7boWEJpzEWs49LwCi7HeAC+JEOEHBllf2szQ9s8GemuC91ewSeYvRJ8
yxbsv5cKzZ2kTkCovVSK0R5+mNoNcrkWH8GfaJoIKIaJ901Zq5jjlHMQs0JoJwZVFyAwkzpR8Umf
ujHFedyem3qWSh5mD6Sp2ObFUaYzyAeNadX1bUgPDw6p3u9ApHmn8NubgzEWDF5KlNBbWjxVvr2a
yhJoZ6NNtzz1RJb8l9WBrqPnrAuRHj0uHdSZvxRxWb4/qmL5GeGQrsyCbAnZU47EsJJHPFPiuvIc
cdc8OI5Mtb81ngssVoqVlB08QIh4qLJIP1DotAfJ/qUzPUlVWSEc9MK5UkWIboesq76NRthC2hRO
zlbWF96oD6+ItoMcrkybPdS1x3bTZWxUmf25tLJp77asNjZoNEVCkm2x0BGHJZw2ev+t0cdyj5GK
QvSalztiwPj34aJzOS5xUUAzKRnuAxXf8ZH8qeomtCmjn1D6+OqI338T8pYbfwu763e6WzAVusYC
JUpUEpmbbz38Iw3MOKnA39IBO79dMbkpDYg+VQBRCBesiEsyGvqenpxOlW36InPT+I11dChXFcfu
ynb49On9lWBjRNMvwZaWsfBDNoNim5//WG537t81A9AxR5w410uZf2k/kUCBQk5kNrs/NLPUIoLO
g5Wq4RK6RHmg337skxMYAEJnGWX6bFZypLzTIEhobkgkmi04nC1iogVZvvy1KRmobVF37hTJB8Pi
A+ePUnSFZkh1664Xa81AAokRttmHXHMIJ0c5Jb3V5xGJKOkqA8CFxRYKnD35Ax/izCsIe28DyXL3
7SPJyR3FMmAb0jePT0qIJOthpU/e072ouwtgVaAj08S7iH6KCkT3M+sJxuF1OLYk7m2+Fsxxi9MC
DErRIMpKv2Fv4FsU0Ef4a9Yia2A3XoiO8Jr23TFJda7KN0ZGoUWAgMVxRq+d39IDIK2ExUFl/eCa
dU0okNI3KJeNfXwhhdrV11n8IOdzAt4lCFP79KkGAienLDT1mWeDkvNb0IE7GunIt3ogPPc6DD5O
1rgjK11KsN3N95eKuT28C4cF0BRaSoCTtRIntxUle+GOpgJtooh4Z0W+vhS7oRUzjpcolzrap983
LpI1dYUs512J2+35R+U+xbQ80kvuB4mmff6s8AorkvVabbQDxR0/xO5vasqa2HA+K8mMkDpyRo4T
rG/SV7QbtKUTa/cuwL2F2dnKd8JoVeAql25DV3c0Zal81uVIIeoK4rBqDlTNMj/qzlgdRI+/Hol6
mUihTeJvpXez4MNgGZzIu7J+gRUvoe0Tx4Sz/ykpTEdu2QhGecJpiVuNsvZTa/zVZhlTPvAWdyse
9v51yO/acCvp4zdjz0+G38pF/wQqyX3p1xBg0y5GuhQIunm8a7AvFa8norsRN9uB9mTVDCFuCAew
ubuwUU1ZUjDOZOyBKuzFCD6+kNF9swsTccybRsWFZgh63YeLTv4OR6WVW87SxQJJ8iUfK55PAl2P
kqwaxmEqZCTlEDaTJ8levsED/41WmhWgxTPn5fDXJWW9j6W2ATPeX0gpGYaST692tPjQBXf+b05x
ofsvOkJ06JiqRxtud2wX+Uf9OiNR8mfTumtIijpOIYW6zLF6utkH7LyjNfqJpa7eALapoPzAWtzN
cIBXvjQoyC7uUfnHNGIZDAy+ZnLJfgDwMLq0E7L6rqDHVNzW8pg/uCzXGmhEMf8IB2k6TIzynbwb
O1D6LMN9pqCQIibqPYIqtwffD9/1ZqZSsLRLhMTl6fEXnQFbsyJLfIUBvTuoaXLxCjXg+hzhLAcQ
G3lT9jag5zrWZPGwlo4HsOPtEdXLUJM/nOncQ2n2ICJVKF38rzNqpIYvG/NYHTcDNJPardUQGrdL
sIxxFAffrg6kHCnnJpbAxFqkdnFeIY1ezQYKjALiXkEKOcZfPtsSnnW0lC9PQQgMY3iXRja6mmWC
k52NdMaCznGaluVt5dtn/FZ49XjBM2q5epgh9lSVaDcbtEdcgPPU/eu5BfzyJ0iAMzqoQbf7ftu1
j2udCnJE20415wrZjt+iNK7iOlx9aIUR8c5dTVccZbBlIC15ZgNSkaaMbgn4AvE7olc0OGMX9oDJ
xj3gskIHJLure487/fcZ3doW415hxDh3HSFvzHuYT8vh4R+Qj2Ld9mJEJbn6xXgETLWKxGvryx/9
8pmHDJore5aY4SPCQOk7MMSZ3PeolVAkmTvE/J8Ii9yZQ3lCSyxdSjPhBHoy9+5qAij6IuVqePDT
82e8KCwFKPh4ZT43qicy+qP/W07ELZfWj5LJ1iI/ANFAReTzU2yaqQHtJUI2N6bUTlh4D5nuLEEj
VirtNNRB+p6EUlWjMcr9ZFfzxguRmh8NyYXY+tAKvyRoSYnxT6zIEVU/M+fQqsIQFJ7osQETUexU
ziftDsC4SAIzbYoEuRwFD0hnTDyT8loajigrkBXItefpi1UBsZJ3tybRfpgjmZTLEygOhuGd9xbI
GRuQXQv7qszUMOkD19sjuIWfTbnMtnxZ0mZ5FRYUfoAEv5hNdsPjupOAPtXRFlVhZ5iNi0Cobh93
Xn1Mn5IgOJE+Cy8euU+5dC/z7AT+fOYCVEWnY1Ra5ZQvI7Fwm8m8zCSHqw3JyUD3B+r7WsaJJf13
iGrIXrQqe0w/dtkq+VIjsN/UDYSxhB90SCOG0ww9nvDubhbwjviLeI1yzKAzb8JwO6A9vivblIKX
jqXYuxCJ8m0jBeYeYJSt11v+dAwCTrikPIbySIsl9xIROTQqFnf4XmKqXemU4Pg+jNW1NaahVkEc
1b9ZYBOLDmmZDSdm0oHYrCeeQ6iBFRH7mHUWC2XUm2tBvlPc3q66gmOjEACpPpKrdAXSA7e6GDw1
EsrSvDQnNOdEYy2vRqc7rqN+oeNbzZnRML/osFBu9QoRrT6hf2oEiVKjpkCew/sSLzNX0OMndihn
Ey3dc3CziZEdDNirO//NVzxGLQXfbca8CEHEe5e+KK2ZPuftevdBi1uUlNuwOzyFYWj3KX7ARxVR
2PtOgztTaQqXFNTyEMJrPp6ozPlqAUYvJYBFmcv1vfyu0YYgaRXlNX37SsftO0Qyz+Q+FQ/pdE/g
e2jt2J9AEOqxyoKdSUoT5xhnf4T+WLBD03ZDSliS/Mmc6+scxojBhwZuVbJnNvc1hz6iyUN1UB2J
nEhIOAFK75FkfB2c6+jXcpRehA3ZK83qM+9dqcfUF9gpuT9zwOsQBG6dvf/JYNNDIthcerKCzc+w
tk17mzTdyN3ZFpFwY21EioOgxNGDtyyI+aNTuY3yq2C0Xx8MBa5U1euykCPL/br1rPRenDe8tLqZ
yA+suKOK7Al/3OKepOgsMprXsl7HPOp+2O9ixfQAiT6gSkNu3qOBB4ghGvjGL70L4Vw7QtvK9i9u
rdYIohvptx7JD6OMvJFHo1XCZCtuWqQd6SOckWyJjouWT+30GyFdYG8E2T6ojnuZu456x+bRux4D
bsrdQVPEGHwQJnAY2wlyXfiyDPJI6q2v7jzsLX4nDamSDN6/rcQGIyQbz8jus9Wc5V6qzewKi9Fs
33vjLhxJCtn2um8YUcjkjKTId8nc+2O7XSucZY0B4XlHhvCn2iETqZJNvi3Jbi/1S93cRbqf1NML
ElXsQqq021+9YRYGVNZtym/k+J22bfjEYtwx9E4583E7txTlGlnUS3vMdgp/X3QFXaBGVQnI84dx
DhMjj7dwiaTQs7pv91FDg/J/gXP1//V3pTkGX/qUEzM1jQ0yu0R4b4sQD6qrduwXg71KHDd8UMHI
e4MgQr+H463uEhKXqabfF+s+VFVqLMG4CnssayPERaj0HCBDaqQMqerqUQkQhIEcmr0UCPCVBBR/
8zmZBk6sH8fUr9cknyUZwIzK2R2rlhN/70ZYMAdXo2UdvdS7+DqWubFgQnp55yzlBZ3ahY0QPnkT
xVsKGHt1T0LMWOOP/uemWSDjHyK9jud/enIoxW6/mR+tj6CxzX+rWMK19Y37leR0vEmylW9M/KMJ
lB5BQwXX103WtuV9IuZYQ0Z7IZeLIoiXmacrsPt8IzacZ7YPTQc2iRkdwjE6mhJkWof6atdL/m/p
WzEPJhG86WLMt0iJ7zEeY+GQovp/rO3FArQDaV/70FBd+nMmSMPxrNvuV0Wz3bdDAUEPC/CxD93o
BqBzglkAO0Q3uqrRqvxspPnOLFBha+uH9Yr9QWYjY8DZ7C4E6EpuWvqtmSqjz6KYiG0K0lZ7HkIu
IuEIvSChjIi0mj5lWeWdz0gfhiSh8kZ+iRCSgW3Y5ti+ve/VwWxfgsh2UfIYBbioWoBPY9E2sHBd
UkiFpTrKLp3J3pXyeAHIeXMyCOBpXiVaxDHGroKSn/lRYHiAE/01cvuLsbAkLTz0RFCEhKQA/tcT
cR0pAwvmlPgeVMPNhmZGWMOCSjC1dbgg/z3bufVl4/Zlpcxum11AeZ3u3XhuGfc8fdUktc76jhCQ
WliHC70VwwmGL6FsINjGoAkF6v3JYoXnwA4niSpDlpAtIqDXHrYPyETSdSPjS2NYF8/1xpS54opw
oSFtDt7PH7m7eIP8qNOZncvD9U7Iy2YzbU3ZCpA1YwQaXddpvO0b7Eqx0YOHPgk2s57WWnNh9VBF
WbbTxSqLpSB2EqvhLGFyh5G99NiNSpLFMbdGSC1Y4XV6Cdsj83PTB/lAQNl9oJJEQ5CbcSMacPn1
+Pmp4KJ0Zbv4IkhLfidVHV/WGsBR+qpBrizn80lzMV6B57vH1r1gAdLEMXjhrzwdEMDpNMce4kZ2
nBuYIRWxfZeB9t0x4H/RpJg2p7W14RVTFImSPgT98FSSPXoSAWARwvnYm/aKsTzao/08avG2t92m
47Rri7xs9/RDkz3pruI6CwUcCYArrlozSSKWzbCR/II+1wF35Ut15gVSgI9tcx2OJ7rMgz16KtzQ
7EpfkegCb907ilY3QuQ1KxG1H4vJal/fUyhgCCrvxkDt1m2wNB/hJ19vdV7sIAYIA0RC5+ScB5+H
lZSHH9qptjM+OR96ZA7WJ7gV2DYayiyfZcbaBU+mkud32/zNCYz0xA32aGDViNVWIHgpjwSIG3DC
cCPkXD1VP1o9kx8Zd+/xsHk2snFHGgsHvR9yIki3KB4c0yAXGrIRMlZysSvMCH988HVQc/7Tfav8
HP0fg9B/DzkJkQhjPzmbx9ARHmMF2EQ5bp1kYg/WzZSA1AbRS0ou64ytpF9+VQeYJYpLhKjnxVe+
jwa5Ma3SXzLv8eSK00Bhrc3sDCr1gjg54ZqwViOealI8/gTx1AL5c+H8XA+Myhymd4Hj0Qkcwbn0
zvMe5wNIdeXXO9Djo0vpKkLW71uWaBorxnsqCikBu/f3Lkcv4tEOZRk1iNHo1OMG+MF4B397gEEk
L2F2D7a0+4CGKzJfItAsZ7LnORYljYD4ME80JCq3XEgxHIjmB122ZxQC+9tF1fh/LHf1RNg1RXgQ
f0KEUr3QKsdd484qqNgkutpDCj5SK+q9xdgljGrkDjEztCo6e+Sn9FwP3qMAApNGwukoFsrTJoGe
9kQ7xBYTa7c62eSMPT9a2rn8wQ6XMr0h1wrci+qxVjzttMSsKqEWOMVADymaDsPF7NHu5yH9SK88
8a4XvyfLx8scJeRr34+eDpiPjHlq3TFYpV3RU+rr8uahH6vWcWmBKs40YDPpXZJAgDQhSK48MQnj
1wos4jcVftpfvtxoc0rg1vMQvXiVfbIuq8I4lRVgNCe2glwwngj3sQnjba5cndRL5jUBLV1OFS/k
HB1aJCltc+aaKsHteebo0Eqk9F8xlXHW7F73hskJ6VJFkUZ8B2NzyyfikhqEFNQrV2a7nw+N4CF4
h6vBe0dGeIhUgLCNHQ2UwcX6/fK/w3LbUNYBR5Zb7CLhQnNOJnCEPB2SyQpwsj1+EfvEaghjdGRc
dru6BL/Fdfweikg6V5uCr5fYC9dVKFH2cE0AOam7DdK+gCDU5mJODdvntLqGJKUtYO3NaGBlXxcK
zCPmtaBIPoOoIcn27j0h4W/4dU4n22Y9TAQfwChuZ0CnykR86stspgt5pTVKdHw6ppFZug8Hr5cy
CcYkSQ4CCBChC9Uu4sAxZoVHRVJzd+Me3tqpLwx8Xm4KNn831QccsIXECdLdNWzUhSzUcu0Ul/aE
y6wcWu5lm+RyR6j1o+P6VgxaYM7SpaqND5lfuTq6BSzBlM8UIxSviMCZ5iubXCA22hszdKSiTCZ/
i/Mi2uh+PLUBv4cJn9Qdhkc0AAQUfqBYQ49Z2U+9vQmEAR6Ca9l4tmzDGpzaH9WSie1z78+tp6gB
j54b5mYZYokTY0lKMKCPlAQi9DSVqwV0ftF3ztlrZ98pgAM7NCN5kJOF/reDsZwpPUCBB1ASArLP
1XfrtcSIGlRFh17Y2iDULr88ghqdMuoCpByDgd5u78D+9BTOSU1540+KOfpyWRA9g1V1ipPZdJAT
iO6LS43u2BB7E2o2qSmc4lpR0qlfYyvhoHEGDUyItrHpNXc6R1PlY1DFFT27SdOlZ8r5AfXZhPVS
lONag+qOiOBU9dx+TEpA+EQa+CJZOkkhMVTpgnHLuHOndsvqriauTdoculR14b4INPB+5smtrU+k
+F4Rxv+hnnStioqwP2Ld+K4A12v91jIN76NK/nxEInfJfDYuqsPb6O22fd+nT3SfL3CCPbVmHIqy
Mxz6NTTsSuWkBP/5FDQhlNCR7EzFiuFqGsvi24L733RtMALFnFaQ7Ey1UtSBw8CL2lmaXkJ+AGKb
QP09HamwWqgBqy4oTQZxmMObcSKML//kBo9prWvDEgxsiN9W7D67Y9hd0TA1TYtLORSNae28AP1d
/FDpkWoYjV2OzQoifVL0Jqh/r45EthhjbQZGPNWByO8Q53VpGJOMRZjtJcq5M/2O72No7dm4j7R9
4/RBPNYn0luK0TDFqiErGrmkq21b540wIA1OBDIRYnv4B71+sYRUquCfDiIliyoLb99lZTZYdKlx
gsF00jOC0jvBsE8mOS4TmmQgiNUSwNjk4daEh+c86ByZnEasstKUcg5veUs8uu+om69myfpV3+ym
RDGYVHUiExcohGeiAs+WSCqK1XrSzQiXWNs0Y/3++KVRgPIOPZFXoHNyw3Od8M7rdiMBGjkJETXf
VtdXGCwCgfl0M7U20m61nPgQqvTgBCDlx8zXmOLCwphzcTb8wRteDG6E5UmXcWmNrsIFzrHvz93O
1/w3D1WjN1Lm6jGggciJ6155gzW36r/VXTvHltGBKgfx3ZIrUv96Gtj5ftt4lNl5KIfE7FPhoT4K
L0cTwt6OkF6CORKerXJCzyLh0L8ouEKRUTpgZ39+k4DBrH0abibLhpD+/uxLjplkQYeDAuSjBKat
MUZsRAW51J2Ao5sIlWM1ihcc3+gbK8QoNa/xm+babsSXBg4R0FoG1KJL7OFbaaHH5XvP4UibSYvj
9E+D4U3FSdHnu5/3MvI/fFrCIcYZnKAp5srp3XU0B1H2+2dVK4q5JJ9PYrIdB+dDrjfocs66V0E5
S/tx/1bXn60mLeo/6/dWk2zlU6cTDr09/7Ci2o1f+jNzdKVmGBi98UrjEfxJL6oz/4HZMe87v7wp
IlVRiNCiavHZd2HJAD+RREmyiPlPhh7r2TJwjoZFfnxHxkK5j2H8WZs75SFn5/7m2xk1LeFXnaXh
xw8WWaHTELIF+CIDwmsfn3lgDDJWvwrbeZjPotXKI9snM4bNc5GyjlcGUgchaxSCHPXb3Y6pubjs
x/pnOSDHEuG470AkKRo2oJy8ICIr0FxHaVwMh7YRuesSdkjnneJAV5EaY6kZsL+uMquU2zKLlBW+
TaeIZZFNesMdsBErVmrMeNotYblNZL9GtADfMClDHDiaUL7Fa9TpWHFD2L+6sXsLuws6ozkZT6sf
MuztUk4OA2gL4a+s/P0Akm8w1koubmVJuJSVNgHvGdifM1inGijUx3XnqGe+cWFCJoT65IYD6DcB
nqYYI2Fs+2btYnoTK9chSSSdjQU7llTlINgbvSzFvfNKtmRVB8LSpUS01MI6PzHyNGeUCVDEDAid
xsyM3ovP6olcjOy4/c4vPEiAcC3lJdiHYaWVEWo/y7o/YaTgztYSt5Yhz0BBNrYPCL+qnVLqQGil
5UhbF8Np6pOsniSba5kikIGIWA/qUAmzqabySMQtoHyutjhFJH1wJIrdpVI2xVDRwJ1iM0xw/C1y
BThLc8pn04swrAP4YVNaGo2/H0J9GyM6obXYJqqx2n4k8R5/QIDeKIXY1GPik193XZAn2xl0MgFg
rdFJ1a05E+RnMbmz3JTrBXX5iFYgFU2JPmnKlssZIMr0xrK4sUAmVhpyYviIJA7R3Bsx35cg0NcY
MqbwkGDVgvN9TlYGqxj5TFpyKU56/GVoEopl1u1C5FX8hJ6VT1mNKfWcjVwpYERk0cpQxMo/rFvf
GhHoNo8uZoWJFydGhLh88ETHXZyJIRI3Qsmq9WUt6IngDCsgDQcQSS+pd+l7EtA0RNKhdpq2rDGO
CRS38rMxMgZaFUaMWSrh4T0Q2Bg/4cHPOtb6i+y2gQn96f0rdxOiv0a2+34Paqzkkle2K/4NpFuw
NSMRa7MsdBLHEo9HR4J4JPIxRkl7iH1zXQzWRXAg0gxtrJ2c3zliku6FL1doywIt+aW365j9h9lD
yZFCqpuCVdliMNVlNxn2AxdfpikuwWYSaN2bO1SXg13wrRI5I9R3yxU/DLcfLCIMRbLYkqY7jUwr
qefgaixtJRKuw9IOZ+GDcffl5elI44PuSqLD03MK3iDDlb2IwStxCS3EyfefAs6vZmTHv3Q5vNKZ
g1QsNnZrLfisK9xUNKHpOWSv2XgMN08fZGgqGSlfAU9YJfTjDvWXsHjKIusVo6Bur2VQzDi74LWT
o7Qu1NmAPb3l3wETFLlFlQU9OKwoglFyTRHI6biQH2BNR7qd2IeUpPDnDIsd1KesWFDnDhPHn6Hq
ftBYkWGBSTde8DqpQJVxcwnliuTdbD7IwMOx21+YXo49bvuMOXDnuIWyevgrI6JQtlGba1T74BRn
53Ibl5IqJpiFhVMgqeW0LCDUm/2geZrEds0B8ZO23rwMekujKLHx1MyAfEYj9iXvTFeRn9SOreCN
Zkjw+8qak6DdO7WmGeIcmXPVISYjuhf3wEEiS4H9TXlmIg4Xmmy2B6ayCPL+7RRaoWep/d8R4DUx
Z1fu6kauyQ+2vjFbnh5FwLRkzAyBOP696cjiXz3ph65TW3qfMVpBhCEhBmRJnuQFwkSRDjbu7oQn
kUEhUNkVwyG/YEhsLmhN4b8zeUCaGRTHbs2rQgGFEd9+VYY56lEkmkQDduvIRO3yd5/QELQ3QKzB
RdzhQpaVAfUPF0yZcnxlqsb2aVQAsB7RwjLld/j5/2774HMEFES5CByXrvWNBW4RQpoh6dCxsWVv
2K2UlTEsvL/Q+Of7kEJEICI8KGLrxh6ZHmqh/w/KJZ9jQhScK1KCjq6iVT5quQ9/3rSWGUSYvfCK
5vFW2petpxU5yIIHZIxvusWrqEkCWEtKUIAbFzASbc/Dxt5vkn/tTV9049ZVfJnAPQhuRJEe58K1
ubaPCSSeuWE93HKuYTqRnAk6HOvpM/P/A8W2cKr4+3U7m+GITR74s8hVPQejdnmpU93rpWbYSILh
ddsfWmWjtYVJVUxCSJ4RqDeJ0wrrcLrFZxEun6SV6UWeRLLpRbEB5Wad5nb/ct7APfTHU14bx6SQ
LCpJHnOcFP1Ap6M6vEbO4dG1aPkaW9mZVnLspLW5Lohg454VfhrUtjQQUbMMYCFqREqM39mDprmH
bGaXb4ki6YsWPLN5VbykgRi7rWm8RBstFwZifmtHb/4PySXM+ZnNniZW4k1KLjY7UgCkMxIpSyQN
1U/0MXBWQPeGUN397k8DQW9uWzr60iWHd7hJfobpY20nY5ryZYk3DzJ31Ob7bdx2DwDPeSFTxt38
YGmsaP5epZ+c+raplVxg53EjJVNXw0wK4WwimD7+hgQC1LXXJvfx0PYUKHjtk8jJb0XCzIvFL02p
Ek3bQMCK1+QD5cZziiGEi79JtEmy+EQiGocCZwjEP5FsHFO31VFxgHJ+flGo3274Z3elKW554KlG
pGZrN3qwo3U53t6dZ5eDS7cH6k/OP8TJUA1dr3fssBAujivkQz7D4lvggQkHMvZeNr0pfAM+6aqg
BYDpD9SeY4C/h0hu7fKZVx+UDNeflJRImwt5vUEvupFcFeiPyKGg0hbEExhksmhTdSpZLOwsgpSu
Y9pLvPpYIm3YiPynIMZLgRrL3e0UeuvmRmZLwY326+QSLbnBbeYXJAcjvE15HvAgYOpJ7S3aFrnH
9z/D5x/+PixxcEYc/yogEp559JqunMmk3i8ni8zO6n122drycxux0JZS1w+CHZuTx8JdBNqD0Z3Y
t7WCI+JQ8zzpwqIfSR7/Luso3O68ZfFjqoQUO6ZLn55aKPGpDgg0ZU7PmDcfmYcXm+4+A/uWVbg4
19S+2sep7vyL4ItXxw5oohUdAuxpkZ4+AnGFYiaSQ6DASe/sZ0cSGuXhhAvyynpWWh/QVZWPWutJ
gbgdept4LsJy5l7CTIE8bW532g2bBJlsldV0mMt+CAHmFBdwUsUObeorxWuwaTptj/RI/Y8XiM3C
Fvcb5cYjnRe/NbuPOvZwPlIbslf2r+Fxu6PVn1KCkrqYbPa4IcOj6sV62Pl/A71SMVh59zMPGYsh
PqmXfGzHn29xRQZZqABWswVgG6dJvqy90J/aTaB/w+eXd8oywwx2E6p7+5q3mZ2u/Fd4GCBKpmIu
O075Mb4fMysROdTf1B+snwyRz27sPeo8ksJalCGT2LVD8W4SUkG4J+1VtYtAHcR8wXD/85NTdHub
XcO9e8OmBaY8LeJx46cTUaTGCL471f1eWp7uRWKjvchUAJmjfU8llmEbRKRWbD8yNDL/BNHw0KA9
PTFGhAAyrgrId2fdz4Jg/KPQ7ABEdPbkIbCB4Utuxb4XFJZfTuV8xSjyXxTiUjGSlYetDV0fedG0
9K0husCB/hBkPUEtnESgcgcUWmcNq/kB3Xw6ggr8UFe3ZQOEi5kJ08xfXUyEmc+COtGUuYhhDcYH
vZ+21moQsCra48/pCRWR20btp1d8sSO7J6hO/0oz5Y4qzoAnRwqHaklyH9DNVhZ8y3x/LEbJUgel
rzF/R4VyUDPoVXNVVjGKUP44dw7qmfDDv7qNTp6dVSCCyqmbFjYlRDiEr3IqJK/FYqVGFw9fsRGb
ztmeCLtVC5itXAs/Q3l5c3S/W8kfSGruTKvHOjnbpNfivJrPZX+l0YM2pBz5gRv+g9sbQQBKBruq
8gpc+hWJii3I7SL4MaI9SI5/1eXtX6nfz0VWgcoNodanF967nk5QJws0VvXzPbRSCQoYw3nY5yyJ
G8wSgEqblAQeJbb0QcKU3Qs/sjbpnI3SeUrDUrDWYbQLSCBHP91MbzUbNpp3k7blwCYO+SBnOn/U
5k3/DDy2puXDZZjU7rVQWSqJ6IB3uZ2utZlQ7Pd+3+b9WHBb9ARy6WdEeEM8tpaNPgIuKgK2g9J1
LMZbwGEv78vZz5GQssX3KEMLWfjqPmihoyOY/V/qcok8KMa2TIdg2b/WblyqX19SSeu0DTvJtDQM
zlj2uXS6zVUtTFddX4WuYWoHzVVZkLbUOj3PNtSuXZ5cqU0y5yKJ5JWzL0/ZdqW+s8grShqdkYEe
yjATduemneo5L3Sxl35ZHfHRpM62bOv8lgfu/nIMaOY5Zb1kk/HEmHRDwmq5ly8zme6z3YQDWF0q
YgLOLAx0Hy3X/eyS1yR49uCVtW4zUuzkgqZKnbehVWb8167hucpspHgFBedUnp9zLmpLNndD6VxJ
3TeifLaza5rw6XrxkAwu4Xf4gcRwj0GA/O/oJBSrOacUYuC765bPSXAiHKy170c91MfzldxFfc0V
cw0OaKD70iwEnGqcmpgmjx4qEqeeB9wrtRSgHVwJxqxbmG/1dKInb+5Oebd4yEWg8rxgKlA6iprM
NugUuMDw9VaBvWbPJ/ahRU2LXKkUo2h++bMCgo0qdWSoOCAU+mZuTdPER+8ruO3Gp7nK/ufrZC2E
5ryHaGMjPImCUFxCWgISKoVl3qdzUKiXUiidIIX7kT+6XIuSTl2WB2eMfC5PSq0nhnqZbA/91L0V
JtwUxaEbJIWZy947bt98RQoh5WKezLteqGYdT/N86b4oyGpHCUm7YCyYS6gfI4w6iqUav6k5YUJu
ulxRqN6z+axIoL0LVI1zrCBP1OhkKVRl0m/TMy2zN1I705PRojxapZHgByue+ufU7gx2kx5AZKnR
hKVZPQGzaaxuA86+PATeJX1LyJtkLdurVZDyyS5wz2dNUADNMfxeCIyeIf7NrJTU9Uil/MopYO+X
23aoHavOs+dkbwLqXLy/gr8yC+ooqjtSe9kuuHYrp5U0YCbK4gRouPBsNyVPVXHSDoIKe8Jz4bwr
GleoKIVQ65YQtuiv5UmpBI8UacT3Z+XFYEiOvjleEipLc04y2/dnpLM9RWXawHGbs6n0wHggjULX
TC/jTWIrjUEcfCLa5DNj4HYuITaBrVCuNLn6HlRoC2A0erS7vTZAuFf6xlmUk8gz4/bljABqVudF
+0H/wnRV6j7FMjKYrSKMWv+rwB/NwwnldYoJT/Q9Xcq3+EPOUJLRLx09cdvvCZyLdXsYQNaOt7Zp
4UBPmo4SoF3vJHXXHSACWsa2E+Rvlc+ZtMblkmYzA+Pk+03tS5+TJiDWeIAZw3HDJjradw6BH56M
nJsUaPJQTquk6TPvAnm63hqFi7WYm7DHEqGdlF/HKsHvlBGhosF1m9m4WOMmvx6DTRozdIXTQpiI
JFA63SoRRczCBe28P9xKSl23mcZitDGu23Ir6vlcJDbloi1F82hcCwYB4FxcAxqOLJQTjdtd+W8M
SSbbwNxne+pFIlFdtxerOeIzzPZpS19sEp6fVRLCDvNwN5VZnW6YLnhE5amQ3cTRrTj2un4GRxJc
m3U27GPSyM2hT0uya+Ns8Lnxd8oHc7zpT6I0BaAOhNohIn+aMzglDClVwqo/Y0GGS0nFG2098qo9
w5bhcVeHGI+cue7zvsKpyKXUCNVCJ/TycYeLvQ6sb8y/elfBIzgDaiFT9v5iy36Z6o+85//Tsz+L
IvZ49fIyrHwnQhTk8NG2wOesb4um8u7y2SpP5AMjGWYWMZcm5DKJM4fF54dgFbjX5l4iAHU2iM1L
BCyKJxKFyTmsEUAMj1AB6xf8Ft2ynV3VMOG8vKl8ROKaYiR3a1RaHmR4gOavEaartAqNIrhNBi2S
UbC1E2GKAGAodiDq8kK1PTw4AnZyOwcVYV+j8NIvngm4jaB3SZSsTJJRCgWMG+u9TNd5Zq2K4QgS
1hO1fJf5Qo+9kS+TKglyCwB/4ovjN0PTNCJ0TqAoi+af3zdpbEnJnUWoE9NH6AQHMH8DWQX0/wrS
fQ4XJxIxIYd2KY7VNISlA+KZH7yMjdlb6pI6B2gYJGbWCXFkkSlmqSzg6a8UGaolo+RxCTL9FZdC
HQPjARvDfgmwC9W51CfPd5ZZWYzhtBfCr1etTFL3cxezpSCJkSgFl4QEr67tm6StGh2hCPZ6+BVi
a5TDBww9SwWJwh9cxBCW6xhh5e+AQDr8/fv7IOfDHc6jM+nzyIcedERkAPj93DcnHNDSlkCafX6W
GBApVt4A1zlFMb9Ma30aEDFpqJos54Q0tv1Upi/Zzz7nrtBymjGiJGyoyWIzJC2Swp5Eqnm/IO5g
LNW2YpUl+PMgsd8wGTbDtCoCUwxHwz1tFUsEye2J1Ma1/hjMVvJ7UCvNPSY+AxTDOzqRzyUExjes
aqYHpRGUHTXblVv+jG4+Po66pY/VXRCafku3CI0y456qxL4GPWmLU+O15cFwY2YxG5+lNt+8FcBu
DN2EaU9aKAZ+SeRIdRNnThP2FBYBSPfYftPFOdf/5v0WkR8H07wf77rlUG7G860liLlQyn+rjUZK
081gbVArUELabqho5EciU0KgIdoWH04ULUPgoeQnSVX/DnH7ShDSgiT2wVcdjYyeKPa0ATkra22Q
UDoqjp37xovFWcegN9fsHZ+StmNijz5hoX40QGyqHAlUb9Om/UPSjViv+gwQqkOgyRVMhKCkHTM5
wMk/Il48695XAhZQ6W4hUFS81sTlfWFIa+o1sU9Z/A+zha/wMNqc8skWuJeJIhWmH/ZA1Hbte94p
MvHo8RAlyDGExY/KljNq7n+a5ulj9UfZgUJd9Nbn0YP+qNPJmglpNjR0xsICymftz1YrnDen85A5
0M6WaEQjyLpYcJFaSkd9kprNtAftvGNKw+ajFHADBs7NlXL/FR3T5/9UU6u/oUClWOMEzdv7wuEd
ETX3DSrD9hN+cl17SGT0F+IUvRwLmW9RjLXV+dGagk4mqEJPPBICGXLO7qM/Ear/6OSqVORp6zYk
0M7rcutu1N6kUDbRuJvrSTYv0edkA8SZbDU19pHYSpIQnaSM120Vn2gsHauv4ankx6DPsmVcF5DR
En4i2ETXZUftXbzqisEfaGpnRV0IoVQoG7r2g9Wd1z9BDrY9zYyRh4PT0l8OH6ZPmTLgYVoeWxQJ
0lr2rku+TvtlwVAeWdRiv+tpj1vdTfVr519Xuht9XijpEYTOOYCCZx1TIeqX2n8FuUWGqlT/ZID3
yg61nsDrGMNThe4mqw+NGzndY7/wgwn8CoC+3t3UJxwJVaKQUOIMBZ2Yr6qN+EMvU5LnRGKXvNMI
j4BmZdCkluWnfNGHzlvQPU5l0CdJf2G3aAFXzE+UbA87MAwCme+W5+WPtjyWBg9+GIYSxQ3i25uI
yM7QPc7p2lm8jop91sY3Bd5WdnYIFz50/FseY/3ctMiiPBlnkaUbJdAFrVbTfn2OLTdJRUoqy4Q8
xZLrDh6jsb09tsF7JVZtxYvrG5OpzTnwYZ1TWR0gyErk19Bw8lv2mqpQl4srAUH3A+/7NYGx8Ewd
HpDIFmkv5A6fnDOyXAuYv8wRQnq/rIyIqYSm8nledyhDTgJ6HqzqiWMwfpKsuWSYqDsV/610B2fw
sSWvyK2s+QGqm9/1ZeRdfbWmJIA/23V3K/oCeod58eMItruVsI2FsglQBxmpoHmWGiXlPcTopdKa
vnc0TCuHA8m09qw0DX+gaCVEGczRQ4/cHvGJn0g44sdFtvYVJB+q1CttN/h6ni10PQ1s2flqNoWe
OR8h+McrL/L0lG7oHjCFbkwKdFw7XVVTIyqKBN76Qa2GkkAcAl3fAk9cX3jrhQwzakE6jTT/z1jy
l4KHsrenaDqQLcd+D6pFarEgjsQrWDdpZCNla4CdtHdEoITON3kjEO9x+4TDgI7jQIHps2rDh0jY
p2Q/h7HqamlIWBqR/pXDlgNua3A24N4mH38O1URuKrAIe2qSiKKYWY0dDKaCPUayQvMpTIBCos1+
WEp5KScNs7ynhopsexdEFqcCKaLhwRBWPQdqWDCgHxgOWRMysHbtmkYt1V/3riY8cz/PEzq3bk3E
Vp1SXvWrkSMT33GyfIvEFGyivdho9kmbzmMiHeDBRqosnhkv2QxA59e+8M7XvPloCYrNX4tpJmxu
oK72Y9r+SRJNgLrtLruUaM2+/n2qVLyp17FmFFob6l/6pkesVTeE2o+b42H7JC+STPRHS354kyeR
z46VHmYUv5ONTeAoxjUV5NhjoaXdGaxBU5ekPut8JbLmBZARCnSDIqhLDf3XRDVwgo5Melk9DQYc
tYcPmNGLTmbTmLZ6MkUBiCq50LY7v82MjfuQO6/uTgXQPJqncWTH71az/mXZB3bDjLhMyBCq6jc7
i6CHazFLxEw6sDU0DUb0qTRl7ANV+f5rOob8X+sgmaqmjIGN+jny8QMAqsoDx2qL/QqA1b/wSnJr
W9O4ENFLu8T4HL3rXNGULMY3J2ZHVz9AQswSq8+Vg92JIHD8JRJ4/z6n60OTCHkT07DCT3OQQUct
dEfdSXPPp6e875uyJjfGH040UjDlH5F6SX24cfBAKoHCqohRDpvsaGn2uq1FYGUYT2lA63PDaPNd
VAMapYckij+809d+jUjkpuqLsCHKL7bTCF9aSF/M6eFbri+73k4odES3i0HlV11UxthD4LKk9rKj
VOzAI9ULUNuqhpd/RVbRr91G6y0yMcNasbgTsNVDUzd7G3LJeIA8NUdaFZ4g3K89HO8fPuqumCCo
hscp+6DFfL73ZQB6jK8cXFXfdelMLnvo70caFclmPOUuqBM3OLhesdMYnIQpkhDFEkKvH6BceBdA
P2FVw2oBrBcsIibR2vkg8X8LGdTasrOYKUN7RhO8LR3rahpV0A7DLWUMqaGfazUep1djD7GKrFp4
EH9solL60eITpLqesFQP4sBe2kFKZ8svUctMtESC0oskKpxgJyTqy/vTVhzqH0R3Qp66Ym4uqjBJ
xJy5UpRRvY96BnPRrtF6OCEBGqW5T6AcmUqYtOOEiVxBs3LDjW10nuiOkBUmDJhhY9RBtLbmAbxZ
GDwm7BUO2ef0WuBUq8U+dCJrYKrMzofCpFEqX7eIyaFIUAjQ2W8CA7DhuevsnC9P8Ml3rvX8SmIP
Vf0EFV3fn8fzs3nG466/2tEJY2g2VSYPLrmCQtMBIRh2rScVIM74XBQAfc/36W3vBU3jhDK4Muve
3NfOU6ObHsQrWusv23OrPNNyGdjlJeJNjAw8K+Z47t9Hvb9p8xaUHGZazbzbxZQ4sRksgtl1qyqJ
uunW8oMJYq3RMbOW/dHY5zPrQNIXdRUtbACjsroD3ABQGmEScmSOGDitl4ChtcTYNkorerB3xt51
nTX9qqkuXAv84pX0NkiPlbDnY6Sh/ouK5z0QwWV38x6satmDLmEEFIhV3BaEMJj/7o/ImdFbWmcx
MeL6Zd4OjWiluqFRbm5OyBtnEI6sYt1qWTFUJz0MiNYjECp5xXh9pdiitmh1W9CaA4v6BWZZRWTY
OZPPyI/AdrncSyf9Y140FuU9GF8pS7Foajsei/jVV7+WDan/pF9JSunxTowPWO+p4RSbC36g14Ps
uEHwpCwsJDi2hRh9IKyXRXvgUgbFTyN/w//ZsU3tO1fB+kCta8CySIeUGcb2gMfkpxv8XjjwP+Hf
Ydb4i12WxQfCZYmO14JtlVTeeOBsPm0u9u1RcK4N6MWj4LYtJuMcoyp1Ml3uj4vfdRq+x9lS32vM
6scDjKHiV8/K7jzoEXeL25cjwKyqH0lONj4A/n/clOWfitc3w0PRjI/hAulwDnMub/hC/zDyLAoK
0ktUaDz6h8J9HLR2TNAPqywqZ49QTdQ4rb6S5eLMSTGkRJeXwcuIBQquzLZ/O92EBa0e7i0UEqys
xy4WyYbvPSh8aQjJ4ik/fS6qBsfZRTrefLI949E/WdXSPg2EFndICaPOvBpqIOMBEBfL6UlQq637
Tb2ciXWbyM2zRCgMa8e0IvNNyNfqFRApT+nhZHEpEtfSYiQ0bZ/urNfDlTXIBMuKH7FCFa/r1X82
hWpC1uORP+O2fMGAX5d9LNeCamvsUcVCwfUFA1n9oCe15nAwLQnrZJeqykSHSIufy14OAMOP9AzH
hEGY4XRL29+Xz8pCrvpVnNzQZFfbYlHyjW64INqAEhIaG47jQ02TTLxBu2Yvtws0xq1lsBsk77sa
wle0/QF7/iQhyAjLvYL6yDA+9wvZpv40P0RixmVNMpSX/+rsxJZ67C9rAmfVyI/2W54PU1agUIYH
s9XJDqDqGdR2kpIsoWAvYIpCW8P6psTaY7OLmtCCE7F4FVvOX8lgq4IcWv6LA1gNOmWeu9P5R5J7
nZP+i3snOxoOZoDlODL9Q6iZx6pTnvXVaLbdkITzYZqUFxXFaJJWr6Nx62R6XyCxvykWQi7T5in6
t84JLwsJ9YnK7fnfuCYXHOFOABi9KnCV/LdsMfj0GZP22RdE5expFsI/5Dkp6xV7hvSasAEv2tos
EwXg/nrTgjNnTaU/tUXNeWL8i2593BGXc8tfqVYonM6WFjejaQ+hyKzRqlG+N6ZGmfhD4p4UYetn
0arANtH38yHDhtgpoTzLIai3Fcjhvd7bDcKqO6NiJHFmDDF1qUbTYsF/WkcgK8TGOmrn/58vbUE4
lgfuMoLRB5FC/4kdvMpPK2ZamABs5fpQiGIHp/VgUqgP6pOjKHzccU9m9w5bPh76SRk0Bm4Lcooy
cxhimYs86dx0uoSU51ymvwdb6MVotABQOozdzkmOZKL44/zTH1Duqr/vuVqRZ3kxuOA/TPhFnj5y
bUTbIEJLKEQfsy224+Rj7moHl/flmr/GjBocGel1yaZucNpA9bTzLOZ4Bth5hzFdTcbVlnLf4JPU
W9d2msFrXB23G9aP5LNJ6qAytdA/hlXN3CYHx2uqpp01bckOJXOMWIrALdd7SSFEW1r6vFoom5go
7Lyyq4oIHDDErBbmSi2qtj+1jOJloTzIJULrBZ3IcdybGbw/k3BmWDPXeVnskhV7nmtgQvfrvtE+
EO/ioHCxlvq2Wkd+n3P1stWij5pMvqQ7gFMthUlTlC58esmFIuDR1vyzkQutF2Cvpf3GKRZiNv8G
mcMx1Xz5FW6btpRzPGhxvzNPVw1+G3G69QiFHno0z9xwo9wonV4xiQtnCq9RTFt/EX0rZT+oyj0I
+zIJAPDjCYJy62VaBEvgRI9GHuCWhPiXDzgZOJMSN3MdPTBSoYSiZp3XXEn1nfwYVR0R7tws4uCy
762RDPJrnnLFDKWHPkBImsGjsApOopRUrdGI5v60OygljcMLn+NTkfI3PJoqECCPSxxV5m6wAQgW
YfqBFHUxiPwosZyiuU2qUqxdLq7VnYgQ1uef9go+JboiL0rXlZLPOmJQt5NXRz5x8mQ0XjORhjfE
c9gMnkOZDyNBinyVOhu1Rq/3E8tQ68xu513YxjiIFGtIwDd5JeTA3ZPcZJiSHBrJzARdr/ek02Tw
55LBU3SY9X695UDBom31sXFySvNu/Bl+MzRcU7r1zjZRSqNwruqp5V9XurvtP6oNuEm78FMJi3Ma
YpnQ+GQkyw/PbHgTv11yEUMasA74H/5186meUsxK+vZ3phHl33cIaFMHi4iiEl98VIA97RSu/l7J
FZxZhJYkqRPCyBcL9ngcBNlnhG68xLzKkAe3GsTBA3ZgBMHboGeHGfnjN7H27NRyOIQFYqAZcV7L
lG18P/C+lfIYZaxVBP/g5oUg/lzVXNh007LoIqhNMy/7gbthCB2AL+REJ9Ntb4ATaYCQhsKTKpYn
LdVJeNuL/GEqYpAsFcOjDBAsGry+9VIqag0wh6ix3ZqGa3fJiJ+P7SeFOJsaNK0Ej632tgU5sXYu
+1M/5Pu4dL1v3VQygfkv74n81bcKC3pyo5C3NdAMbqb+EaBeY4r9TbiY/+ynJLIqgixdzIRQQCtl
E7q7GBrOxVPFWba5Q0bGf2k2iFF5Atc+sbn5YHa4y9nxclp4b96lH/eZo6q+5Z6XoArXidw9hCIy
wboZkZTtUeqaOkwLvm1uWTkZ0+tMMxxYY/1tAk437A7MDTYhvvN2PMjZ0hxAM4+UyVz6eHLKQ28C
rCzEeb3kKXip46Q9YzYEhpcjxxw1SG87fdyFC2X2FNypUMZ0RYjq+rvbRMGeprmQu0YZqjamoHhK
7Uxgou30elcwc3QoUcWsv8ueVpy9IUMXt87M5y9ZggrosskAjknBvzIhNviBQBNld1CxTBSb3EAC
GBtlGG0WJA5ljIP4fjLcUmmqf+39zC3mYLYzMIpBeluyeGig2yUlDTgbiu2nykwrLOQ6yzIK6XRD
563Y1rW/65xbLtjF7I07G5cqYUCFmbyQswResf4qOnDLoSl+bjwoMMVvqEFWfVEBUldFmG2LYKpL
/PYg6jW780p5WoXVBsf4sdt7agLm8Mb+b1f2QjX/mbZbSHQz8whItezafpbFngck4Nex9+np2NNP
9QP4UdR8TEgsjUfjJ3d8AMmy0ALaGNMjrVnewj5rq2cIECbCoiN2wFqiTrCI9R7ixlZ6zoGKGYSN
QlT1dZgAp43d0T4IskaepBWW2FtrjHd09ROp0wBRuhz7eTFewQalDonk1syBXQsyf7Q/+OiDUXY+
A1SMKDfpjq5+2Ret1v4o0VxZtsJZR1e6vD8v5YWglkHjCrzAGLfF6pe4VCtW/ALdmsnsuj57bQMn
iHclEweQiBBA6Uz0VcAbH+6z5/0aY6t8MFxnPgx8d8KAoJK/vEV1zC/FWLSBuLT0/qrl9/g0KY/Z
0kVShqLFR0U4DyBqSYfgQYC/4WXtJoBZFryjJCydAnX4KkpFLl2rjZ3DLKwDiCMsvex2xD/NaLv0
SBKIHicVyiJfxEprPKkKfbLdtl8KRZbJ6NklGxp6kaR04ke4QIMiw2+uz1Ox3ttw6AjHoZv6DVNG
peqIOrRUee8RHa+lehkNlkoPaF/EdwRBt102nP0nhv7X9EHCLxJweEfRB/4j+KMsiqXWzSWLzyq2
WFbJ929Fc673+V4+vP2eH1GGuD6lA9MLCpIy2LaYmbxOFNVw0ldHg9Cag8vr52bV5ZdBZ/12G5tc
hk+ioOFbt1nH6voTcS+TUr/8/rMg5Kn6DbqUxgjKyjq5vBaBq+7J+QTRG9nZWwvOTo2ewAcOoV99
mchQFxWm1d42dGozvDTWStERJzhynnFLYGBw8QnRKhxth9naEj9SWXykQR9ees+nverc4hZ5eRuj
bGWFq9VdhVCy/PShmS3M8Fp/48WNPFOtUIaYnptBgtD+N7kj6oI323WCLYUNUCEtje6P633OVln6
gQzKI411NP8y5ZOx4rX37Os6yey2BTb59GZsCSSGuHKY5k++QRdgG7XXQlR0QEbzho9/GSTJ/JTV
BHsMti1YsSmahxJzcjMnYUMSri2Q0Oi8L/xzOqTwCLuTj9yuN1i/EWOSwRDGsY1XdyObz2eFxlmE
kJ/b2DMiG1iijBhUuz8BM3snn6u2jQaLe3418VgsBJHS7c88dWSGSNUw6ya7BLUS4+t/OexyECTO
bn5zyIeOFUoZtAlm0yy0g3OM2XwRjxMZGoR0w83ayzfwtG+sT7wwrtM+E0JCtFevx5MBRxnGLKa3
J0HiXtp7w/rxj6wkFZSSxmiqIark0VAoDBaoklcwoLQSjDjm1FN7n/Kx8yHbGrNXVx/l1tAdosUi
jriG3pOS/mwS2ng9yoEDLheEMlbZyFstcrNesOJxpTOAb/MqjvnYIR0SqMUP5MPx5TInyR5foK+t
F1Dd3jTpRrxsm6+rMN8s52MtydUAdYqVl5RCDY80PSxtBUfVfYGuFbnzsTXqOOVISYSm9cl+ANLy
IEM2cO8S/atam4R/Nk3PCRK9JJR3WAVlyWJGBQQ03fvcRKqsXQw+BtCZP2cxxkKc0KDJD84h32LC
7FSLg0xC8Jr0FAumr676Y4VAfl5S/3vGDJaIPQGDSKnIvF1yrDvbKIibhuBYZcxrWGa1030taz6j
HulbIwKQtOFYWIMKg9V0YhYc4d6vBLx9+0k0a006qDjcDdRmUAh7Y0078ubmml2mKAiB2AALswyH
x6b8lsu7Y+1N/h88xfIhIX2f0KjxuOv2L2I/j5xMcuJaAVzAK8WIUIuFNuqD0woWVZWjUVMgwa8a
qF2694Uw0g7tsCR6Ykg3mx3qrDMJyTqBpDEdwiCTmOnQ3Gfjb0/k8Ng8WBhYpY+I7jPS6RRsXzJd
z0PMnZJWp3pAnDPPPSxZe/bK8Q7J/yUVCr3ZR3qtVF7/ki3JioABhfrwRn1odBEi1wcIpfvKZOeB
2GGIXvpLgvJkxxA/Esh0oT/rNYw5OYRS519YURG1U8qZ1ipC/hEwMnP8Udz/pa31tVopoDEgx6kk
hARwPGTRdGzd2++zX8YSWkRgI8pjBF5tfMgLjej6OYKCmDFKV/qBb5ejBP2vbue+2YnZJP3ev81p
nO5iocWMU05bBLiG7UryTNI8MNhAQIFpJzeeuOluSce60CpJbJaesN1guWEaEXtDsexrd5BBXgLa
/0hZ1Q1LLAJrJaPU1x/sb4u7ZpDTxIAdUBf/7AWqWqSrZ0lLIJpJhsHW0bCcDzfRBHoF6ULDYXmI
0nv80gSJLgc53zBpYd23s7IJFOYkj7xK9mXrpzQlJvLHnkle9Zpi0olgnBQOPoicBVJkXS3dh1sH
AP5LlA2MoVMN3BrO9Ccl0foL8EfhDy2I3m6F+8hKINUkZU20O6Df2RJdpOx3JXSfNxsac9YGHc0T
JJulVRfCr9FV7M/sI3Ak2zA7HSxbp7NT46seh7h0NnnvHrnkXg+08dSuEmmiJpf7uBD8/WCS4cZV
PPbvYSqimRvMLEha8lqtzniVOTWq+yUFVZpP7cfqu1P/Ypk5oNn92GTL6CKQHGuI8nMXwAFihHWS
yQF1anvBD4IqmG16VwKH6GmS+WG5FmCtg6L4wQ2x9pOmqwqvUyhTwTLw3jIoLGKEycOTQguF8Woe
eRSqC0rSOwlQjNfWb5uGmJLez639/sfIoTMZ23SgTKUm8weWAnQmyIJ5MXHIJ9gjoe6ROv7IUVA5
QB+QwLBowjMFPjsoiFh50jhlwBg4fyJz4s4hshiwHYRBE0hEovol7o2PaxhfoAqFrxqnN5n17k9l
9GEtoQPtsKtXZxpfY19HvQjhK1dhGJGPYFZrA6UGdiHkQ0HXIFrnnVLzkyCrS/kb8lS5qKCH0HL/
iyIx13Crp6QkxkCyTZJw+8tBw9c8P5LOhjSJ49+PJ0Vu2d/DAiawhfovluw0euGCxRXMzgOZcfsp
J0PWQoK7im+p9JXXTvRXhhzlkN4Clvng0xVqKvLnNFrqoRVOrJFwBNj7+eHwOScXFgea9hUqbxlO
SJztUyCn38qORkAnMkCdVwgmSVUhXCI2x/CauESFNhKLLPOztjM0S259siStq4ADuUcEEeGIfLQo
qeLfw1toSZk0z80IICaqTAF1AQQspifkJNDRi30H1RQN50LvT3TWEvnr7lJsp6pFzqVVtIbWb1RJ
p+U0VicRiv2sEgEc+FF8dNQgnu4iq3jmPSn6mJHm3HGkZLsqDCust7oqLt7jnFocnB9IoKKKFGOx
fxaWpABQGvarOxl3R+1TWuKl5Kr01o83USaUa/l8An9/fd1oSZhGQb4EguV8/OOAhpcJZb6pstkR
Licrbu5ujMeAf6MG9aJeChzIC6qaAnYtddsvYIjgsR5ijNvaigrTwlsPjnt/HmlEE8Wtctqwwla+
31o0kHLtHBDkcXfdXW4+1SMMbg76pCmcJrxiCwCfvtQ6Ds/hMSa3wpW/qkdK8mPVwUduf8gtP4la
C08rzZsk+vH+jy9xgx7qnMlP/K+ZGPAD/NhhnVRmTGq4I9GYY8OxRGs0pUWpEO0j031UCCP0j1kr
pO35envS4xj60OasGaqpygSmwhmUnds7yjmaJWwMzklu65edN70dkxJQ32tDy9dUEhoLTZDpM/MN
3TOqMRvBIHcckzJHXfStaZqOOdq4mkoysxiMZg3t2uz4v7Jey+T5TKwn1SoJyit+hKQCZxcqeKxP
3nml3sRxqzx6Ur2sK8QZa291g92srhVWcP8zL5l2vz5ecCaOvwKt3XCXl3+yAy2Z0LTKDQyrwu0O
24SbDKJk3aP37Oa1zW95Dvhi6RV/lCRMQCri9N9W8oHlj7Hrvawgje2A0ngcA80RRpo1ZdF3KwhI
KoH+f7PtwRvXxmF6DIsf0AN5IXBdI19Av87gNDMLDDu7BgTrYZ/OnjPrN7IvubL+oD4+cS6g11mE
2vLOrZo81cM7it+x0RPgk54Nq9xLZSob75J8vTw2ODBkkst34rSruYdnGgkilMyUgRlZ+2apTuXN
ecRCzOYDm3oBs/vVTBgtbTCnjKN1sjFpa6GnNst+/3zYu7Er7dr/7Ldhak3+CZsvU+356hlB0OXq
/gTH1HcCT7f7eAFMlqufpDEiycJMRzOsTNTx585tL+K99TFmk1Fyak1VtPhHSkeE3rdPP9Eh50Xn
PCi8iDz6gzRZdqRi/E/6uIzS6wcDU29ElZxV9yic1XUggll2zKjATkKPVccYWbSSCDXOO3hC746I
dLR6GHA9j66wRTN1VQusxGn5Tyd85TiBBp0P6xAjEIAm/USf4hgSIrAV2moq/s7qNzAYdEV7nsQt
qdlwA9GEUR2EpO/2+eh9EDZhfbv5T5FkNCGgOLX7S2+J9E6kVb8jw7yT/qtQzLDzuG78t6kc/4/b
e2q5p5n/J8K4mWEl/7u2MN+DuXEJuWgpSoKTnc8VwMDo8MtPUSgjYjpY5px/aZd+Bl32FCV7SecL
w9w1nE1Bu0vJcDdKdY9z5EnVvrqE98+bVrkvGQHuhHObMEl2iWwPhXGh2HSSYe2xPOduT04koX0N
aDghiK/NPUJYUVAQTLwt0+vxH4gDFoc8XAMF9xK5YrV4C84DCRB3ofKw3A7o1AQHkZCpGB2h07O2
isVtAcrJoZeXEGavrwe/aQGv2ZH6fkEWAYpNy1WgJbo+LGQUjECxDYSyEc2hsNDEOcvjdhBuYB3Y
7uEm/xPPPQAoZxlhr4GLm7TejLO7dkpWOB6bs6Pc+8Eyna9isaRV5EcZqIla2OqDA/9utVOPDhsH
Tdvjq9FIkKnCVSAAJULCR7+fjN4NpIwR+NdN+hZFU6Jk2kKxVCto4hhdl3y68lXSgoS5K9B5dIWK
qwJd3sRZit7fuEhRBXrwTe4+P8Vu09wYUjztItoIiEcFRgjvnTYzTYkT5ePNKGt7Ush1re6EsX2l
IgyUb+A7ZjIy27IVZgMICqh9JLYKSE3Nm0/KajrcARAdS9q3VEge5Io7CjM8CxR9rhJ1dEUJVwBI
iO6SPjHrwRzbgg6swIV9K4lyR77oaNXLzU1uVD4E6mShj3o1hyF1KNslnhOaTVtF9PD4RY8lxryI
JOotxB1TT+9w0Pi17hFoe//cojbuRG7fNU4ZrEOy4nJjrm8oapEd/4tUiQSvRiRcs7t5C/UvG7Zj
1Suz/FEv9nPkdml5Z76ntw5duDs3LS/la59DKjYDf+lQXTsappMBlaTk1ukW3znx8OsGnTjI2aPq
MwoZ5N5CBWfzzYUypVdfYtjm0J+oSb4u/E/oyuv6B0RwFgn6KDGrFMTW1bKU/Zpwuf+UtMH++UR6
bhEQaMTz4rAZb31eGYiVh3zCDRX0M07vfxJpz9EOz1SlFc2YyVJBBXVQjC+Ge6Sf5FMN2Wqvg9ms
Ju0MfxG+8j8dljwHULLMj/9TZoLJkZnnb6E59wHkJ0P23J4etZJx6eGU3EQr87piI53aHyypI9ys
YfYc4rwr/X1ndsBse4OCW8oyxwxx2AkxjknrvX8Q3rDigsvfVbX7GpYtCw8vrw/CBDkWvT3vuQq2
1iCSLNjB4SUOWUb4p3eFn4fzCoydGAoOdRFLcPYKvqFMk2p7iXvhy457b+I7RPrND+U9kY7gvIeP
x4g4tV5BFOHeksILV7TkAkQIu5qr8PNjVoSQ5igTXv9Ewr7J/lUvS1cBTTSiGqKICkLSnGYEGM9t
0fezi1l77Ur0IjwE37997NZim5Ufa8WIxIS1/4t/9qmCtdPOhh3sQjIGVRNfYVDAAWf2ns07GftX
mQgsm72E+KEcT/b6dNoE03kRf8cSVMOF6zxnOAHJvtBmQp2CUjbJurkkgmthFfwJybaJVld7f/zM
xTfYQ0RtH6WiPaIIdg06waCB7VBQ9uYnQYDD3dNkIMYSXg5zLXdCN3KKKBX+m7kQajkNGNDM/OCb
jLhLRjcpLX96ltMwKA+FWXTZQ60r+MtvarQDdr/9lxJenNzmGspFNUFXAQK0GU17ufAxsR8Ot+Uc
3rTHT9yLxPPyctbewnGYvNZDA2AAHPHZMNAjcJ+yozSWIWZGzYZ3JN7cI4AATj+MO1hnN6fSqEy7
9288ROpPaKdlBwAuEPd0NO3IEmOf7v8ssnPGORQZpPmN2WRiAFEIZdUo0zt2it4ePLCJkF5lUDk+
sqYqwsy7qqaVXfoiW1VJys6c2eKSVRBe8HRwF4gudI4el/VJFn05i2OGRSCmmnyX3RP23/IBVLE9
EpwTXDkrMydLgqyjdNPnSveF874TRX1+YEmJt4E9VcnAhOdBUR8P2hJXRE3iHOpYojc3lVWd5YfT
XNVClET2C7mho5Kq3t7Npl3eyKhQAr0LYm8Bc86Ff44xGzOLurf1m94C0A52yK4KnjWIYZ4kYsKE
jIa8fH8y+yZC8ZMnkeB3agnifWtiKXWSOBYOp+mkG6EzyCKsLqVnIVxIM/Snm2l8pW7t4XW3LDsf
PsJLst7KK8kjkTHEeUZP41XVW2zADAIGxHFQZ5MxoXaa3RUCJfxspywuPL66fOerO09IQa864sXV
soSTm8QbR7t3FS/FtT9QqOWmy6NB7tw9gW9xldRSgrgzJRfs1LagpSpgNszpXZfmN/7rqj41rNgS
8y39deqLE7mkExyxyKwFszApcnpqTMijz6HZ9woNu6+n7MPVS/l0W32P9nRukf4OSxADEgoNi/wH
/cRtGKG/Qze5Cs6mXmW2XWLfdKVNNgmaTjbYGWqhEuIBKnX60Alnf9rpI/E+cWURaS0rXgQgEd+D
tgar+Wfj5VJ2z3UEimYOvZyanFJ/kT17ZIlnOElUQJvTc+WUcbjttPWfYVAoJpGdtZxoFYaQGiFr
1eVhBduf5zXzUQlmrDfVNLQGPjgdD5CkTAUs4ju1pQMKphUpMNI2UqFbawJVLPeg/PCufaBgNzP8
Zo/TPI6IRUkAFZE17Tj990qNYKKWsqL6MMQRFBgEpC+NLvHRv5DfC/aY2avDNOVKR9GMmTyKNDos
k1qsOThrS+Gckh8kHVcj8jry6XAS79nRiSks2TdGEjF64OPg2P5U4sjPM2WhAqpI6bFfYNyWW+/i
iGjHVCMdZeCEi6CHj/QYNQ/EFEFdxXO6KcK9f63u3TPvBPhD0R3kkS8LLIaQ1cz0NFFqcG6nyle9
XePN8NLofLKxTjqmUVxn0F06Q5updCUTpoyRy0qtHAj5r1y99maDEOz7mvCSHlvl7cBEK7q4qCrT
MpssJBKlRFvNu17jrkoKSWufoxjiIqFI66LiXvIhfFT15UutDd3tAQFeZHTu4Yc7zpUDxaoKDhbl
VOcXwjUIIUYT5L8gi9Mx5JW13ZJzf5TGeW3l5rZpfjqnEyJ/Py1N6ALSeK1O4wyrpG7sLCOVUDsu
GqBdvGtpSQNVcXVvRb6mmhVaYhwtS5irsmrGsWJ+KRV2Kz3lEOoDm09dCytMQM7NRyYUGEXEXeH7
iZDgZA6vKKLs8B279dTarBCLrhdzTUd2aNRoWWkpAVthV3GW7kzZhWS8aQediqloYiJvOvyaLuHi
ygvaRAN5GwZ4/lOK8NnXgCrnDgU5OAa1RE5c/VSCRR3d7KzurYrLfVUe3+TDP6MOcPFs8My9Jezy
D2mpHJ2E+31HUI3gMSswfIBRv/Rzgvy54zPXRlY/vOe5N8HUOzc0f6BPI0K+WSQFhjPdWnk4/RGG
dLzwnuOFEbai0ohOnjjMBK0NM2FpiSdfR8K4OaAUPLDJU7DwOyP5l2tsSj/czsrZKlNLrNpY8+Mm
83BZsOGxBiKNVoP+isGRyoG823/iXbWC84hHfCHdre23m6PKcIT48hR7xug75tYrA+SxBYCTyZVI
l+wgOWXPDztaDKQUiCYU61CHLiz+wAg//2d5VPUmGuVzftj1MZIR38SHDZqD3yDM+J6GZyfmqTYR
2XhdMCsCsHBZSUKjpPx/J2jcWLDLRtDO8xIpDGLUt5dlMWfyvb4cF4Oyhi9jc7q54Dxc9hmvLcEG
P9C+MN2cBSHhwzFfkXvTc95EZs48il7Ea0uJLjJ/8FwXTr2M+bw0rS7mjBiTuHPcaPYWE0e3T32D
OB0jzJs/5Cq/vN/Oq94GH2n8T94euOMoYxqTI0QzCJDp9HRJ14G2FhC0f42FTD9fNKjNKEr4C4RO
l378BjWs6wSd2lnk0Dpxzxzet50h5zn+lRRe++nXyBZW1Xeo2gll2n81w1YsVkv7JvFE07zrBK++
5TVc23EXKlmk69hBQgpANSa6yhROSKJpdNtBrsD98y9E0smUwg2GfBvqUh+lmQ8cTXRfHgeg69RW
zEPPMrQiwWrCP9lAt+yvla7WaHfPs7FeO9QCdQ6pwQUDT3QC0Zmye63CGarwHDH3SL/b3Yn+ecPZ
SfZhlG08fx25oU/1GeL75sHGNj8rTdDai1Ac3vMRNg3iRCWG+a3Usu3M4pxwQalEwG6QXsxsRSCN
M9XMIBDpWetTLex0wl0QRHhdQfBIMBrtaCuIbag27DbN8+Ii+o2A8WmyrRleugiv7hX6zGHp+dLX
tH5EMjgni1ANUwU3JtDGzmP22keD+G6OfSux87y6bq6WZ7vYmI38hAePnCF01o2bT06wPnpTjPOJ
GGjDAlitTjm1d8onbo62BdFaLir3XEZXSJ5JcoQfs9A7sGcyIqH4ywwk1a1Wvua9NVTXN+NEpDlZ
zxdbXpxsD87aJ9mWXbSf6pCbR0SFWRoir7TXVu8cparS2yW+KQEJ5WCgefLaPADt/TmWHvDaWXt1
9CmnuafqSsmc2Jh7vaYRK/grAMNP8+OOrJVQI4VIgDMn42MT4jR2FrmS1KWWz3kTkXyuHpHvjDTO
Owf512mI3VuLLUAOfc7/YBorn5c7tTfLUCKR71nmWR88yreOPQiok16FsxWEXRR4Cw4KmQLWsk7o
gPmgGu+eXZFBXGzFllQ0ry9NAsgPhN1GNco2zYEhKursVPogpIUG9VVgk3aHqdkHBgLEnXcLvzVy
38Sef9zoQmZk761rUpsjXTBeMSjOPWflYyqWyxMxF6AZdl0EI+9/+K8gaR/LQuKNV1S9O9Ge2xlT
1S6zGnHYydic+IwW1w4JJrCoUb5ms7PKNCaAx3WMz++1sjzb6ADtnZjSUpMlLIANPrgd93KtJpbc
fBuDW1NaGDbBrvG2awQmRApmVkRGltdgAq6FjbZZ+hAw+2yhiABFRMDJLz+c09qJSj/RoZW9bWa8
2ZCut333ldxqX9ZQnYrWrZgh1gOIgoDEh3cklrVJEUTx2pjWTkDqkm1fxcPbCmnM2SA0SZGFiPIR
8otaM/17J7Kb7j/IzsmU2AZtGaaQzPz7ot2Fq0NKX1a9HDKLMpoN/IgFPy9NMkW/3EiejH9uZd6k
ZuopfhLnKSEp+0GvW+hp59Ddxn/Jm34hTFB+P5IQEekSSYVggV0nuKjer54W5GrKVHETwlBMYbcQ
6V5gBCv4+8axxT4/XTk473NpwshbMi/H/3KQFuj+VuSm5TmP8rOieNmXZvA2aWfgGiDGAHQBbRDq
rtPx+7BAWYIyczT0GXA/rDK7I0YlC5KjfRYsMr4+qHm4jcbWoLHSAEu3X9k8cX1jmvdcOw9Oqi/M
s0wnqY+Amc5okmfucnblacQaQr28yccwj2izkk551feW9Rlov1AVYM/Zl+rN734mVCKBEGwmWRIV
zCcPmwrvmyT6PM5GZZLB7COW7eE8y0pK4p8nJTegvtCR+aXHKpH1U+GOYC4MRbE1iadhveyLJ4Bg
FxVEk5aGhtpVkzlGqTVKw17ujVYXSMvRfWjfz+HTnT5kVDlYpzi5AcTcd4RmF9SDzFB8WWBFggmJ
bZBNCtr4q3s1/cAcJ+LjWVwSH6AJzkUZNX851FBJtizXIxT/Jru5qk51lQDc+RZ4rfliYzVdQQb7
EVTWQt0GOLVrZ/Rq7bm+05Cym0HgGhh3wgEkB3kYnJhyNm2FhT7iMVXU6B76gHNY0kuMxwdL4bE7
Ke9S38ysNxOHfVyVtVT1VeMA857mFT4/3tfPiijAWc5d04JiqP0Ed//+ez1XjhXJnUQU6n+EL88W
CH0mac7mgH2jbmDav8BNPa9jvvrxwUvi90Po4MoDfKUoXmCalTWmBBBM9sXS50v6CAGf5k+mWMoa
oYbxgHvj7hRoWwPmhTdL+dP5pJhS8M9Inql2p6lfdjApiQyB2m1EwPXl70EVvoR8lxwEL09KYFrc
gfnnjCsrgTMLLLMNIdRVx2sgQ4j4T2mrws/La+D22xLbM+8jUH7nfmFEbRavSyNombjXVN6skb2X
/28HkmpIlBv6sK09ji9m3X3NkUIn6cgKP9yjW9UtIsSGhMif/Rr0t2QrG8jhuTMvmTp/o4/8uvMM
c1ZhXMa1vvc09XaqTxLWryxzmiJdZPpXmTFoAJryySTAgH2Lgx77aCqC53RYGZkxAj+7SXpyL2Ex
3ceBR5sU1ZAF71yt+FKt4CZDeMH6etubepVX+KzmEeO4zbGDoKpxBPEKYR3Pjq+B5DOl7UHWcmil
X25DuHcEe6/xF7mg0H+byyQZCB5hxY/Ivg/h4fgCVXu7t7DgksojHihVFxV2EZ3fuV2sFh14sguj
gg8MgxoNHugb3Vp85uYtAWzfNBIreKM21JJYF9hLkkMAGBBKZI9RXb5ATf32KcYLSA7ywRYGY9jw
zMm0BfU8zBVhJ4JWvV7Vfkd/PePhSEPf8Xp/UFerNmn/6g0MPB2QV4RKxU7+8MVgt8MrK6Lu9X98
FqkE7IZnK4vThm9YySS4vQB3qdfq6eLNgQSKuOvMwMzV7f2HwF58/EZUA8NzfPLLRM3RzP4HCxw0
LN1kAomeK+u+pRg71LpDQD1obc1Rrn49FD8tOKouT6o/3U/YkaZqL4cV7fgdY/AoTJtQEqWhYBLI
J+/CoCVGUdQEW5C8kWy+HmbA224rXGBErgxj89RQoGZORiY83OpOHGSJMUBarF212RfzWt6546lR
EcLG8tebMAZeutJp69hOzk/XINaoncOo6LPZzKqStTonO/S7dyoBfXaVJ5PhksvA25xAHRpsLBfZ
eoNttegVqZLB+kxm+NDDf0/N/ykIx9yzn15H29MCALDV24yLVTChMUZK3r2FHsbrn5QN9LywnzkU
eCOWyoMeB7Jnt25HMaMxlyreX4wspmXCMFphHbDjj2C16JGdM0w99SfeG7PFEkavD9AFvC/S/gsK
XB8jR9CNemAgRXRwM9D4bqFHbrryVlZLHuBXJGIBVVvf4IT07KFNyRIHgjsW5ufb20PPHQXhBW54
92ol1vZcZuTNCj5dgg6NkwuKyMMmV6aknUR2/oT4kBTonxqmMh1aERRRXYtegXFYmjowHQi37YPz
iNAvqQt+hyIcQX45oiYaOc9L6Z9Cqbw6PZa2frHhCI24anPPsFhBQRN9FfpHAnI7ODmWisqc1Ltb
QEs2KUJMgnQEr9TvD99pvevmgSyQwrDeJe6MxzaCjQCafasxXn2RBmXzgpKCUud9uTYR1uyUCYUH
t8plgyGhQX3O7+DsXJtXAA402ppUt/FbhcZ6gyb9gjuWVTAkFLICBLW6KtTVECmf86IQxxqxZgp6
dSz7pqSpH0FK94NZ1sEeOYvwFkge+38BT23ko/r3tT7yswv5nBrUfo/2wpi6g+znnh3cj/mchGai
O6QzwrUNzkiD9+m7NwmOM2JFr99l3XAmQZ7ibJa5IVoS9oNUZzb2cTfIcQ5y1EAP0McOMjmb3tQ4
t9qSXlEcN+/7MXbGqq/Gv3ZS9UFSaNPaal75mpYYgQ9PPmVpc3iQWIYdbBEp02BDDzs7dfXo/J9I
w50s3QBO0lzQq9m4SszDWCE0lGI8oHGboNJic+b3uHHImXtj/AW+KZm/89lcL1RG2f9jmu3S54sh
Ht5M0vxW/WaNA/Pa7Ijel40eVjmVKUML+ySexm7+//pVoP+iNYECrKbJ+CtDSUh5GP1AeQJ3Ykv5
cU/eJP9zVo7QjgIOxv8Qsbo+1RfL7fyVUa4NNnxuR/dCrI2NlpVP+1VWXmP7iucPgv7HL7/driUS
fdprZ5ZE0PkVaLPBt8gjxLkGy2GnOo9S2ksjtIwz6ERWHCmQDBc3lmE1OdSOH+E0d/vgI3FByB0j
VOS1UAgNl/4cYEWROtRccQNpXEwzZotBIQgYA5LKpmmVRwUaATiP/i5MhmAlP80U607LMlNuAi9m
MDv1YyCK6yNJib2OpDX9jpfgMgmMvCfWxfoAZ57pjzgowIMLMomMbElF1CN1O3WQsMOAAfeb2PZu
FMxYsCFdKPH9uCQtorlE9UzzEMiztFBNsHag7SykaMZx39UFr9qKH5d9qmSqEfb2306OPQxWex8b
U9V2hSQxIFdVayNozJmMHFGa7SXHoV2xiCwGlMGRf6k67RTzWEZ7Ujc2GVthmwjDiS/V6SMy2jZa
Y4OLi1tm4h30Vgp81B/UhsNVQ9MJyG6a/D9ZVH4JfMbH14q7C3o9rqGGhFnl4/mDv6LNoax8OPc7
Ltjn/jeg9olP5oTQEp7ifT36UK9nzDgBpIDudib+i7orI88ELeeP5yi2OXBjgxduWeq26w8TC0O5
4cBB7twaqAPbBWLEVa8OxyeSpsN2fYxOIciveKMNSCLOi0d5TV7AQKNQbjan1D0Itar9OMISjrOV
buo9v+irgA+reSszaPkvBpdGqt5ypX3dkCITULOABDbl8V+7brkMwsHt/bKpWZHsqv3WSZRMYpzb
abE67yzmzAmIfCgVubiNXG43mHqYi7AIx6medFB+gk3rvSXhDDAlls7gmGXvIQD+CcGkmM1aexqH
/W4YHWTP1eaNBDnlETKI0ZyfFmx+fi+RUZQI/VNW//0wPlGMbqi3rHGpYsn0KyLO/a5NCiPZaZcA
Ai2c0jKrj+YSzG3ZgvgTuVu/ToaaxbrGsPJv27nhUKGz0swfp+AZvIdVYPoU9PW07IZke0uPsdm7
/G6EnJ7au+AfynStO9lo1NDe+5vzJGtuW73gPEO6Jz/CAJoIJfhgmAmfo6Q6h7kRGu0Ds2b1oXuO
paa1I4fppUaUYr3QrlsbNp/ubTY5r67q7y3n/5ZHzFp4t9upocfMRcohghTeoXGBhyiPx3pK2e1Q
aRPrT5viPSVl++8O9bcYoocpEyzCq3Abb4YAY4tsEzeXspe8lk16HUba+W3dPWey4Y7ggySUCNLk
wXaUozfE+/lyRwJJERuBWMz6N0EDryB67fXMnpe1IKEntWNKAzdkpMEEnfl1748roIqx8w5HufKw
0Y+3nPv0xt8WaFNg0eS69pbEFLABz3qoF0alZLA6kT3ZNnrT670pzbMX+sLzDnU77Ru2aHzSopSJ
/E7FhZngXrH1dqE+Vhy1eVNPJUcRa725Qe4q6Qgt39m7f1z6sLaG3KRYM34tw0PC7GkZFRePjJ8i
3yGM3fBkACHblYS7ExB7pirH158NqZ3T2WmPvk6flQlfxM+TRW30pgPqDV1KhADqKTP0JtC+CbOL
QHedBV76IUy2M4iiJ+3gk3QKp4puDxnM3hO6U5teQvxFBEg3H5HfYCSfrY6IF4UCKKfI9Ovn4+rc
zejgx81/hhmrG7INW0qOpTG+qChqsptUJ0qTQv6Nw2RNfmPLvold2PZk1x3AtlTFrSh5BzR0+dT5
vH7Cp7gL/vZYfV3ThwK2AEmHix3nR4ErDiM/k/uD8Fq8BJ3LM3gh4N+tCYefMhwsCrefwGzLGGUP
f51OuRH5cWZXexarJs1ohvcp3iAYocnh1GzHE2cyTtMX872MHbT+Io4mwlAfJBfcX7USjoCPspTO
71N9tM0k5amwS5939p/urbAq/56li12S/Sw0l8YA3DsmpO/F6xQeRZd7cK5e0yNVc4IpZiB0Iyay
6hrvxelwcLcRZ776n5R30Ckl1rlCc1tpz9nFM/XcmIeiXD5r03ixpNSmpunCI0Hk6a4E2fIvFdNk
4jk/cninoY5BomUo5n+al57o5YEKP+9iGLm4+NFD/rLsYEiUa/8Cp/4ocDS1MD7MoV0M+tLhDEUq
OKUKR3jDl5OG2wLzmtbLJIORk16NFBpuWhECBcYCFL7DjmpyrxXZ+0CUaChDuNbWidd9Etn6IZDV
USyOQpsPfkY7Mu7YVh5vKz0aIhLHy0TOS1fI8PjJwH06dPbWyGgHbipy5FdU7eAbgfUYzhS1zycN
Q9HDNk4RCZScoUue7wZpRaWzrOrTuhFq6ohMEsA3c82+S7I2Wl7E+41XES0b9WNtW9kfHrppMFMb
AaDo+GtZsjzEPeREyZbwZMLsjNybr8w/OTy5h2hKKL79+SLMtgA/rh993e5AOz3it7JysdWRKeuz
wj9Oj451gqtmlbjL89km2QcbTgl1LCefi+eHcmNfYnOsG+MAT2WfKDfxSx/NZTgRJ6rjqZhZMZE7
wOvEz0J5eMKi2bA4sBnaa054OVOzeiG0OSIrcf9FtI6GRnlACN2T6ExSbznhaynsaDQkDtVzaAsA
Ny0VyjxZqu1O4ehrpZ7yIbsQP7RMoiCEEj8O75g2WoSQ/E6FavybToQnu3PfVjpCHvr9kx0UgFuZ
PjXQOehywV5Mn3QS5NLrQ9rSWiuLewLQrUYmE6oXWv3zMBJkr3evsy7vOzT8gg+ey7hMqIxGdHg2
GOKafRse8bCd1a5sIxC12gFaK3+I26wmjITee4mRSag3iFDRVd/cDDZaRjXdAMfkBCSgToGjdFgo
LsfHCQypmiWDtiCy7PcCaqJP5Zy7I52krGJ80UOhicwiUwt4WjbV1/VM2BzXEDifEntgq04wN1Ar
WXeXWWHrQgZPO18J8D0QZjwZ065jmOsXMB0WBL+M/8CzuRaDzbSojRKXAU7STIRi7FzK/H61I5pg
+xqQqxUd6jnWg0LsinONS7v5pluq3Cky7qiZt4u5ZZ7NSQL2mKk5dIbq/XcOt4aAmXcxZgxgOxjg
2mhFZfJQw6tF5ruw/Op84caGD1XoiFTzV/MjMbJgym0CmJrdCGjA1lEBhTQLY08uGzjGigzATC/Q
KzJzfIVIdGNXTcnHDPS3PPNLI1X7vO9v5E6xJsYBycHPfF+40edhmqxgDxVQEOD3TGTA8bT4huPE
KaliT+g/0KYMqUhSLnkXkGkg/n7O7p1/rGAggEHq7OYggX6lgEutpxgyPgDyJG1s8MF0lPAm67Ca
ZkfjSQtK6dECxbbTyFG3xeYbJqY0v0p5egLDNURZPvUnbdzu2YcqdaWNmDv5/xvsntO6gGDgprmd
M7Flw3ZGAs42EFEnZnTXyNRHD4rloQaRxiZ8LkrA4AG44pKOMNLu6V7L/IrMiHarEDRVCfuU1uBv
jo2jsF809DvAWwjEOz24YOmCz6gNxxBhvIkYO4FkPSUyI4cTykuor914YDNXLXL87ExqhY0jWe2E
VPUDBQ4Yv37EcoctXz9na6GjiAuBgGql5ZpertXKRqEj0PkaSyVQRQP1TU6T7kW2uHhdp/r5hRCI
QGQefqB+qIP6b6n+HIIeK1o9F1LIZx021xxtei5R6l8wHLny8UOTHvdEylBDdtUsGmV9qE1RQb4M
gR4Aqqy9tpAS5yKThVKYgRUXRAgKlA3yJV9cQkpEm9B+zeKM/W0JMbq+6hPWgI3W1bxE+Bw00abm
qdQxOi34qvKjs9ormHbxJMWBCm3V8MNn2aGFLvvL83sIK1/1RaRF8iJKXw4WI6YoC3VeY2+DCmiZ
qE4OjfBQ9qQNMWnyleHf16tY/P+UuER5VPvbP7V4AH42sy5AiufeDLZGNP7GTzlcg7B/eZPKYAbL
4VaFwG7oQa1NpEmph+N+5SzT7AAtJgVBnuC6pJ4ZoSQ+z93lD5engOiyKDIGJJYeYjQCh2BdQ3Cw
A1yqwm2kSpZLf7cn9dLezQyZCGXfZt4Cqry+sB3RaKsA1ldBee22NMy8mDtJAHcdvNcDta+IqvA6
JTbUzqsQKowGC2NuTZQ1kIS9Fz09yYeeLPuCE3mROGglRLCTK6e1rJZ0NyYRF2HG2cYX+sE3ikE8
k17t+0KuiukqtqAKN5SEqSL1SPY2tTfESyAuK2iFTbw6L3UWAJzidXNkjf5N3hJiHBUrPa8YaZMX
Jixo8KNyS0fyAwDXuzQzlUKXOx/K4PDXK8PKDlyBDe9pXXeOUd6x070JkRXqSiVqOnFkIxwtV/aE
oowqFd4rrzg4dBrNqVgk72s6S6S6pIV5VJYb/ElNHYkkPcps+lzysAWmxMjZH7Z49RgvsMaGo31a
eLIy1krXJ6xTjwLZyGfmFmBmoGVKN/y7hgxMqPp66Fe/VCWDo8d+GPEJ/W9dbFfcALcHgNOsvSIk
LvSgPSpOdf05rpIzBbDkj4SNgU3ZME9p/MlyrhDuELu/6RnyD8XVliOBCfsI1ErGXHPcgWO5O2YK
RUcS8oU+CmJQjsD1toF0Fpnf5FNb7SdiTkoCWpqoCCuIEw7KRJx4JFpHa9aLrFrFCPy2WS3xZNbc
H6887UGFVe2WeCHlMBqAO/QiU6e6X9Lk1GUeuL9YWJ4Stit+jhivlLPIhO7aTiVb2WrLaVji6k14
7CjpcZ8zVjNyLDxSOF/x6S0fAmgn6SVyiu4IZ7YlicgILur0V4uc6McLrFUApSWq1HK3bGQVkhAH
c/J7fC/PpJByLsPhjY+sLxwAUcpuwETfScyCM/U+cPG6Lb5gCa6eYHMhGsbxkxORM6rLw8zLXW7q
+5whOENAHTNUctGzJvjgW8A9y0d45F83IY53LTGr9rqQJwl/HXEnFvJuavXsQy94w7ibHQjaFt2b
1f6mBm1k+Gfv5mdSutCkvZbUddtGI8KaBkARHkrtjfXSupR0DxV4eqRJbhxKbmUnU++MaYi9xLRb
VHGMa3hxZONP2ggC7E+ZiOhpJ0PHukYbdHtfqKAHuKn4Aa0BMRd/4pSK2K+8mOdFW7XpuffOiBFX
QimZtWKBXL+B9nY4lHwZnI8W9cTFXPcaSreqzU3wiNi0tUa3QSRq7kfly+rlZIP8H/0A3Vkl/WrC
jzZVGMQZAn04SwqUNe3n1dclOMIrccawylcx+YRgLHM3n6c+ozQgpwDsYWYHW6YOFloQ4mKAOGyj
BywwlNzuz81YgzhJv+M5FWrgzU6f6KHL5k0h05pEkb1bV+myqXASiH/KxO3FbF3f/W0WzEy8d8Gf
alf6Nrw67AlVDnSFZQ5rujnj3PZiyJxIPo8xoWNO3wqqeb0NfCMqX1XGLcpiUY/XSGY5NCxP0E9d
0I/JOIV0P6lR1d8IVDR5FrFqjUbIL4OE2gJauAmlKenFJj8wfvEgSw/4W5asSRtL/2yHLImSqFdm
CZsU0dusgccUazTvpBEU9VeQw67bLF/nK7Rpm7elpJLr/QbCmUAnGkkVQBa7EfXDYXEcfrrPPrhZ
ePmYU6aUkhDWEkwCSazk1YUTok6BWmCGVR9gbDNcbE3YksHWsqcNKdDuvyXsDLbz/KuBZOjvMSfg
zzJ0VC6iMXzKeRk8gbjA3n5HfyAEJKEol252OnGtrN6Z6xdhXTAsORGmCRu+7b0AVKioHesr6znv
lo2fxPqkrFXedIy9EL/1/+bXxuzt1oYvJlPxIuTNSdT0BtW+gthJMhVnpLCAFaMNFBFS4TCZ2JIS
iGUEh/9RLriOyNvS+fYRoYWmjM99x3zRvQSDkePd3aQtz80LG63Gc90JdsJgtdrZCyZN+ak0kFRV
JDCs0LAwuHOLNTOHXVGtc3DEhMqcfc3PUca05GJX989nu21A7ckcH5/TMAmhupmsQJUlMACxypIW
LRAGIsrRmyfHsiYRJWV99LoXHtFHNVmS06HyNOKeEfx4qxtFJWeoz6MruCfLfauLsbnglCnkI33F
74Q/ez0TMaXv3njKo+wbIJW6HD2VwxqkM4f62497dtsbZUpYFt9cbtiKwfjlaqQFA2RzdPRM6ECC
zTUOppWl1q7PQbNx/osw+MqALT8wRMWSeEqJe9A8EZq/uZ9zL3D16HIL8F4NKeNsLyBqy2ErQ/gW
rHzSQM9D5Uh0LGAUL4K+7WdBJq3G71DmH+z4AxMXmvUFyWyz1pBkhnYulL0yY6OZ0Y661R61tHuw
+DKtXL3I2ebEns2qSu4x41/uNVU4r4edsia2OZbM1WqCOlfeR7IZmvhws3uHYCIYki2oFq8JSRQl
EaOjgw758uF5jV9N2laWEfbx9/slbz6z/MDWUXV0bIne6sVXOQy+v3fg83GTVIRMpQx1J3XCtO8F
qHEOahAE50dshTNdmXtWZ6/1HVCiPeVxpEY4Iggk7xDcTzHxkxZOyJN4B2B7VMtUJA8NwqmNqD/u
kXV0f5QMMa+rg7HWBfwg4lUi+rs08pblmJlRchZIw6mtUO6vuYz6BNyltEQ0gu/t6ihi6UwKHdfC
mua0EOO+5msVAgn2bfv4b52eagcBtwtJ0+gSLm0cE7V+7p0MAeLc9liO6GIsjERYR+PaqXzUds/x
6/U8iAwYl+/q4GksFf4Uw4ombXQUTCwLpUaOSCEfdbX0cbyvkhzuvZLG2FxNXV1Ur4sZASpJdKD0
Isl7Oug3Hz8aSvZSq8X+ku7IHL0pxXu/QmDPsekG8u9u8pYJezmbWiwwb9Ppc4ZM1B6H2eVAVpBr
RsoDHR9g2jF6kmYtXayQnGfi7mH2Jv1QjQTKOJ4TvrzYti5A3xQdCh1vgKJzLDvXsmh96hia/DI/
szt8Qd4YXPRocNjEOZe8OMSR22tSbLNzmZbbuuZfGU/0BiKQep2sEh3bxfi/m1r9KiejcUKp3VmE
zcjp69YjINd9BPfxMlNLhxR9MWVne2WiCqOX16tlgR1Q//IHHXcKe4g/quEhVjN0YLsppaI4nkDY
oZFR+jd7qQZx91ez+S4CVdd+bf8/qKqjC5OXvFdoPgUPuISJuUdjZGkIspYTyFY96F2gOpFM8tZY
dFT2r3a8Z5sPUWxLQr1YcZFyQup4miAKr3VRWMopWuLYjw3IQE4k0FOuakmNVxETApG1pDnj7284
tddFlVLk/cvbN0SOS0vP7SutU9LjKjRoKnor+x85OAAVyLq0P0msfCm+nXjK3y+kmPjCjM+xfoOF
0AyULXYLDeoqeWXjMKu7jYyv99bmfDpSr4kIH8WqyKeNe+Pa/X9csvX4NO2Nkxbnzpp/f+v/rrgu
FhzuLTdlo+EmehQKBtLpYlPdury1qr8zKrVTa0AlkF2iGXFt/Zw94mXX2BLX2LxPMxqhb/qatkKR
q6Fu11vuaBYI2HK4D889bge+Mt4Rfcj0VzZbuVkeFnk2A8H139rvOXVTx7S4tXVxIJtrXUXB42jl
j4TJfAF1zTA4H0SuyVzU973pE5Fr97UPpWKRZiIrND2wPtAo8obQuYwvI0k8HhPN/TnFu85qC253
zBbxLsMCOIxXIGgT8sWk89qhKJ01y0sILIAqUYhl7xyP+0sGcr8AFSoi1m2RUxjwHfTv9queWSSB
pLcwGSQMgz0VaBlnYH/AWVyrYl709deT4/TwSfNzG0EcGVqeKFaeeatk86CneP26FJ0WMAgKV0pA
neLUBMS8mfbs0CAOUvJ10x2zYbYAa0n7PVzkqX7KRgeEvo55ykdgZVafY8Tez15FODvCKcIrM/W+
98J1nUE7oB35r0UEOCqECb4MI6QBH0L32ikTiudhPyr8wvuW/vQ0UI+1jRTKAyh1qp0/5erMSNdO
2p1Ha4qVQqZ/aepp3yJmr0Lv/uo5f3FJekGK8aXaT8WfWVMGffviLk95YjM3MRNOSSyBItOxEs52
+JHHlwbcbNDA+9ftt4njw7w8qAjfG0UFpziKfyiih0PZ+6IAK72uzEm2Ns69lirBivittuxLekWK
LTZUFzY1i8UWk1Fnj2moNXv2luCosdVP406GzvS7+K8ZvIb/bbxoKbxpbTdWKf6E10ZnRvrcr5a0
hFzkg4fMDmPvmEXxSI0LsVxdxw5rl3+RjbPv7F9NAN0O3fbYZ6CtbfZKKHeA2KGfhDidfSleIC3Q
DIJgY5z18PSyiM3q8DuOKgt5UPtTgNJGw4IxhhzrCB0sh1F76zYlKc8/iZkK1tpHec/rvHjURGig
E09TSosT5YmJDcgRw+D+RGpggeMpA/k55Ede0sEQWA6NfmR/U5DERPNFX1N5jizdGQbDSezA7icV
JMUpuGxXVhDSBTGMmgRJqtl0hiVlHVl5IsjwbTQtbdIvRIDtMgPwBcUws/7eb83J91S7Y3sUFUNm
YLyue/AklLQLSxCjg8mywHJQx7IQ/v6uwH2IU0Gis8R1heZaG8Fcsih68Pme1tauFhbVgnqsll4S
AUipB3TDOqrm1CKNO6rJlniHlrNmOGEk8OrBPVA2fjAtnwySfmt4Pr/qmcnlC5co3lnBTR1rN5Td
f9A2ETJJzTDwa4NYBmh5njxP1vcYWYPoQbqqLscYdVb+bK8zRap7BG9yVXon/FRSEwYur3idlRon
7sIq2rQA2zjKKjApWp6YMnQtds2Ezbqip8LzPepoGZTfz4mY6Of63mAdaOzhExIDiKwWqrFNLoQk
jad0FqV+fWWtD05X9NJx1cFd4GIrECICdwoztE2NX3YM07iJEPiSFYq6TCPt6igFl38NyrQjcJAw
gCOxvRanS9OH0J1X/wVevu6oHfRncdV2KtnP9vYUlda6e6YbmRG25ro73Mdjs6wTFxCqB3QJVgac
jFhae0TWfvY2b1KhNjWBi1q5cyJm8eVOUXRT8zgDkF11Dn10l/Dd3/CCks804YrcFTuLW05e89Ma
V0gEnDWR770hmlBGbjCSNEwHj+kO3hEAd9U0zTEaKbTPx660vd7QkW1/Zux6+wmxJQ3FQlkzXjGN
qnbqif0EELs7K7kzzWHa/8giNCWBTwGMsnz0hFTlvpjuzyxPBrY2PeUt9WIaou8C2OVv/TM+d1fY
CMEGxrjaJAQ9lOCldWCQHsOsqLvkmhBj4xkAEAaGPP9axYrkUEM1P/8VO7odQk5bXwimuyHvflwg
7e5wES22RH1ySWyJzefmAEOwPn1p9ANw643vo1vwbyWgbNSASIZ4oMqU7cdSnc6Dok6DN27t0H00
ytIqd+3IAbvxoBorH+4+RgbfYxoR8rd717nybOlnBiFpRMoZsDQ/grEq7eS3d0mJJmdtHmJ0K56q
SIzgSk/pgJmXlT3Kz9oRqVlaGYUqsBFq5ljsm5KePlZ5gP6zO7QpoCIFGIiFG+GakD8R6PZykcii
Dm26YaYyRcsDDOI50wOgfIM7V+5I4qGVpGTpLDFdtHq5BrkKWCKa3s3cOUN4YqhwjgXEoUhri48d
T1RykLcY17KKfPZzEQ6Um5Y5f8aCREOGqbOAGpJbavTPsQVufcqagYbDg5nhc9Z74jzXuAAtsxaG
wDxX94Eg7VO5NXz1CQFcEGIA2V9L+gzba2Tn/5KMAKM91u1NWvrakLucEhkCFogjTDtZ9HpGlI4Y
ST2NXb5luE+F0ep8bhR2aayN0y1mUI8B+9dtO35dzH61KwE8se5o7FtVQ7R4JVZ2J5gbbh+ko3gy
cWTdMGJqqcVE/HnJPRfAgEmvVNSi8BGDwDyzTo83aF44nXj4mmjMjr19bWXuA81NQOp1wDCwiZ+B
6eaYkHtdF65vIZxyqZdXF6klXs/ApmjBsnn+EnPoAUKkW1SD/GhnEczWIOTqRE6Q0u/rBdSNltVt
5BGUqsPLG15cuJHSYYlgHMiByciZcMSqxk0GcykBAlASrzdWDE04oV2n9lLoDoUFrFkty35jg1xR
DLnPooW9jpawGfI1ev4sXZ+jb3cI0PsMm1Smk9PgrrcuLnnpAqhD5K4oTI0Oa+VwDSaWhNypv/F1
EG9CEa//b8bgNwaEu50vZoI15X07ugWYzBZiXup+Eh8IiddJ6X8WNvG3tzemqdBNe0sLixgMnB4Z
bLj2q+lZIpdSP3ToOcOS9P1FaiDGIg1dMiBrXa9iBnExAw2uMpG8M22CbEAo3pWjVNUNa4mM5tm0
dG0EZ5gN/dhncbZnurixsyged0p/4HvLu+1gZg5EDgP5JyKpn/msAIUNptdvcapqqOKHCaCjSaqX
GNor6zxsU0vAVvO+Fe4t6h9KsJkz1BAZlMKpwHBw2SoruBfCmPE+oOjm5sk4wMt7ZKhr2RIROXPZ
mIHVNqFG19GMLPJTIHiOJuBROejbwH9ML72R9EM6V3Wi2/knX4rSRwjF9xIliYU4/qH8NfOYDWu2
3XGAGf3i/zdIfLaXOL4LRUG0dsGlI6SX+mj0TcGbeCEQQejE0CoMoST2wR0ggK2W1zDtQgc/7lMw
Kc4UlwkmxqfFQ8QPyrRLkrhldB1602JbDAPUwuxxom0qzjyWTGcWlnSSaitxYte0bxDM7CoXiLPL
N11Tb5juuHegYGwGR7DvnoAxk2SGrEFoYDSw0eiNgkLl4F92wzA0IVLQ9Y9Qh/s638pgHMSTnRlO
pBRFsUgdhpugM6BusNVLHAggJqciSA8ofeOAaPc+HGExBhHTWta2BofNhgl3R15mrF55C3HcC0YA
9xTNKQ+px+qOTLZmpVeA67y8y9G3lZ5YAnxSsnv5j4HWzt4000asSIljQ4logNfn29kjCCwvopTm
mPDF82Nhq0sVkGY/U9dDAzbTeRWfRbTY2QIan8dCSbBbmEzQeUuqE8IRRyjqWDmydvZgDChxK00i
lPwA6uUI/VXB3fpsQlLWdXVa3bmBvQO1Opay9V2btHcemCtct6cywkAxBA1R5pDp7DtokrnlK7fM
hA4BuNt4Tpe9XxPkWnrEdEkj1XUASXRlJRplaXr/NX6uXzo0BvnDUWLwGcEOoSQpyNwchUlpgvmx
cPaBQjzlcjieky0Jgnt6ovIDr7ARgSi9Q+QOFPi36kfeg+Yai3bd/uZl5gDTokKPqoWZI+eJMfFE
4xu+cBFBv+pfyvnwAgsGRzDKP5fz8g3iD4rA/LVSF5SbW85N0r0kk9JjPfX9AKCt0YQXSylsuHCK
0/SBcv03LUGqE8YqRvzXe93I7kXKOtxqfg3lopEROba38NlfXZ0qpCrAQDoQWwTqXdQHLICT4MBW
8XCjDzpz1+4y2FteU2pyVOfCIlqFe52YA6p6rlfPNRhRGflEb1SWC/kYz+VudQLbRYgSJBJtGdeP
ORaqtz2lytwPqTVfZdNmNYZYlzkg0k2aoyVMepeUms6UuODMjFuLorBsmf3qY2Y2KSovS81SEo2o
ZHJZzs0cxbD7eDgAm9R+D//+0RXc6U15iTqcNkWTPfnghHayyPaaj6tM1VYXFGdtHW1vkERfY3fL
jNuBiwnfjNYE2/p9LHRe3Gi8cksF2RFSYAPF/NTkl20qFD3VZZrb1iNg57nhhYABMX3mrEg7JhOJ
N2Z55wQj29LVNZ+hc73Zi+V28H+sGw/AbUIVMMTtrGvqMaZzpz+V9MxrRh6HJp1G1fLcTOB1sEqI
tw3ZrxrFN1TxZuaP1zPh5VDuzFnZCDGiChV9dufgLpQydpH/7t85PZOG03AqZiwT7KAoBxjqX1hE
V3Qr6bDV9V4IfE+2XBOXcjjE/PFn5eric5dFTVeJUsRjeHQOpvMJmyVvOhzHV0yVqzAWXwoFZd/5
M5vuXA1auhLgGj0ydCrACc6PRt9wV9bTHnYYq2yDLC01bz4hCrmrV3BAcDPuaTu4mQgNHxF9DDby
uAksvMZ+Aaj8YxIAQmQyL5mD49aZQCLCGRYJ/0jmsfLCDTbvvR62tSSdbESniC8IW/OEtcmN3bpv
lhmWXyZtuAPRnwSAHBxuo/J6dUAyYS4XEN6sX+AB2r7yevWFODLP800GglN5/CcqOhxURGsyYk1y
RCZaf1A/YOYzsHTBhK7SuPq5IpDJFDk/G2UBI6G2Qe9cTiu38hPZwdTQrGMINpAXQEZMJdWhFQ9p
MYt8hKXDA95K+5BT2t+QA8i0CM3O50qvyn5OqEl3WSJiWBoJe/bN8dn3mFFIijVwyqmIdfIj4T43
RFz6MdkFySgAxbBAQU4sNvlimisxPH6R7HaUQ3QASElB4xU/8olE6y3rnz1WL6ZOdHTMbUbJskMQ
Ts2+hI+zkvHo0NmObs5v1g6XQr3aTTuBTAoUIeZL9xVh76RbjrrMjWyI7o78+psgshAVpkV17CeZ
QLA567/PW36sBIGniFiHz82jeykjLYhc9AYjVmconjRIxV17U0ywonu1D7QzoEsWVvgqpxODqrXd
z9cjgSGIIknXnOUJ3viCvXpI+gp6/WHctIEhcDxZAbJwRcSKGbMHRds6DHbwzxjqGM/OLVXYGBMp
0o3t/HpVI+Hb1qr44mxou+EpaLbYqgAD2PyHTdyz5MQ+ysXZ6EjDTUgW+ImXBWGsj6PBTVvrSQVN
0cFljsEvkmQbLLN7H/hUg4HHVmMhRxcs/lUAo5lAhlYTOJRxSE9VPxNd1AT0zOsyj8pAF0iIj9pc
kjMxgEvw+5OiBpSsvJXGKKnk9vOXSk7IoxHpnG6TEHz4AZFQxuCCX+tdS5ejWtYMmTR/tC2PKN7b
hZbbzR0XtxbmQYk4RKF5NJkTaYu3a/mBQhmebDN/wr0mW9xojv+LoxRUguG0GVeQ9s8WtqrVObec
dkHR7PngFAxqJSjz5/i54nzezwmtW5hphSmO12ruhH+XUvsD6S9oEMc28/HKdQSSt5+xoNaMPSDC
wGo0BYm9/zM9Fk1s0Tm+kXqP+r2AWfZgcKssrZ48EO4ogfZ9KUNvscdVs5Ugt3EE0EpVEUHsIAut
NRnxqWXIGucZCTYbbDXBVCqGEoVCEy14KgnnQV5J5+tROevy8IlG78iL9xZ/QPGdPuDiiO7qd4tG
oTdps9VckbCnDVzlSrhCtO5PXxaoPZN/omWm0wo22VVKtKhWj8qgQrz1tRJW/iNW/Y3lwKqxPAVV
2kStjILtu1TEYGQMhJYhuO88c02beTohmg87lw8QY5Ql2acerH7XYz74DMg8d9t5koQVVtVCdmpb
3XEwRMwa1Anb27DYa5qd/o3XgvuBggJ+crU5yVx5rf33yG1DEvLxj3BRJVcn61JiwyNroBc9MsgI
s5WKHYeTYvup61u0MhiBKJxorHv+f6dUeRz98nN2HtclMYWMkoYthKyobT42+Jz0RAdfqWmspzeT
Dvj8c939D1L0ovGgzGRSQfTHlxut6R54GjZRX1htcpG71r3WtJfkqwbUB2b6vIMXqwrFgWaWQQ1t
xvBYFOHH5hGx0mv1vrXr0fazoC/Mnzi2avY5iEbULtMAhtFCxY/7G+owy7QvFtKZVrqXNG6T0t86
VjSc36/6KPC4TZMmkP3cl+dtB0GZODd8+g2FGzBltLDydTrrGsS2aiDhzzAsq+4sSHFZ2lE7RkNW
pCVD/Gos7RavpW9FmyesySak8AjWpkY+eGDK4GFJ3cdE7CFZ+qTQu0AVoi0ltfX57cLtmCM/HbM7
0iCDw8qGDLugbSTDnCQ8AFMtm1mmu9Uet54QXILV70U+30D2+1rf/Fo4wd4VlJj6dMlUhfA/jrCo
ci0XiwePATIWO+89FNrgvvy+22vzp8mDtUoQeCwXLoucyaFi/sXBQX4v44/hoIKMV6IPE2KuArqR
QsU2EKCZwsPTHiBW1/Duaow0Hi4X9ZsyzVej7PYavoEnDugLorWqllrPKNmpCurce8SW0ETAzX/6
vyb659Xtnc74uHj3WS3suP3XNJBFaYTZ27g8froM/EHHGbF8lUxuY9WGF4whPcOuyM4h/rkdX+G/
mUEMduOx117PY7Xbe4Y5+CXL+8XPdhw2aVcc5DxskhdikdAFMVB0nqqKT7q44AIR2hCQxw5su9rx
MuENiGHMsaCnnRnKOqj3POGr6y0zDPgG7rVWTR7jBthDd9mnKj7YhQcz8Vt7LTFzrovG3tGVPWaG
fISkLhhTr15uLMEYwSp+H6D+LSr6NDjsWz7GOjh49C8nr8FmnFd1Uuq3G/vMR1zUEL1BUCaMJ7qA
pf5eKBVl8aClVcvEniysKvgBSNnijbH5PXddRaKHVNxDlWI6kq8UFtgS7WS2lz3jvNRXu3MkDDXT
kL0lal4Yn4/J3Tt/Phy5zxznQKFj1Cu+TcxnA9Aq1b10L8NMEGOxtsvumKorHEMvbGC9nX/jUkqt
elVV6vF0lTZ+oIZjQ5ptqxyuv1P1mnpIiVT7zHtVVM5DMqc/WJWnDd5ZNeX7Vf3bO3IQCQcM1YFQ
uuWatOkAyj3cUNaiT4Mdhm5dbfHINgLj+m5OTiiHVIhtekAnCD0BnD+TdoUnyaa9/Wm1GwJrV44r
/ArdgKBMOKFk+jjy1vZ2e6yKTcAeEvz2utuuJO15NhO4sAex/TFrrSMfmWuAFDxr0TXGFnXiroj/
s+GI1UpQUve1ts7iZU8GCs5EMQL4NONv7mS5lgyZiBjhpew24O3JsfXTDOdoEuX6onaZIAt4oOAQ
4f9jn0lxvQm2S8PAQ1uilTDHRuctBIFlXorFIr3Alp3N06FI39zvNf+oIxhYRg0ImPvG09gHQgy/
TGXv6TDTBC1EmfKMUBOgdG/C4C8HwoxNGsDK41GwexTXYdiLkq0ROEzcPqQCzzcSldfc9n4bjnJn
y/5gZV2Fvdw8urfLcrx/Gs59cv9JC7syHIigf92w/h8eR1trQBhGIPDu9qs5pw6A6mYzlhd0gVGE
mRt+KBChFRB6ycx7D9IRTrTAsq98S6OPApUXNjJqNvmeg7huNbi2Ue2t0fx2+yTbuKF+PxdwoB1D
OXiSRkS9GrOA8hvY0BxcfontXqvGFHyA0A20lLI+jnaIbt5Tb+LbQT16fo1TGtmRuCB6wPHw1SYb
cR+DPxSyENMZZAAxiHoYcBDKk/3ar5epcALQzBNxeH2N9A8lQhgIG52SzbyxkjjJlF1hT1t/JIZ3
oZzyYlYRj2epYp4yA58OfhOQcGiawVKRz6prSbjAXwhZP7vi0BaR6q/jRRe7yI7qNbZJ6VeyBl7w
vbM8AF4AY60Kk4ptHNKXlgyiKG0gL7yDVX6WOfN5/d76RgaStWiuB4eNPxr3cnu/KTW2LhYKXSVT
KF1DhN3zGIvNqIuKWF2LyZ0M57CnqMPrBYvbWOFtsMhCvIcn5nT1XfxxOSGWqhykwJTrKsKp9C0E
ElMX0XbQu2upqziZNI+jPH4aXHbQ++3Cvigw47L7N9Sjn7/LmkdIL80aFyIskeeVVThKSiGCNFar
C2dJH/x795khnJ3dTJyv8dprSstAkGWKMbqA3031iTanSp1v6bVQpH3FOACgqs+MfS0rsMC31bxd
9Pz2aPH1I8ICPu8wwyv52KkSQtIF5y0f7lGJDuieI6t8WF/8aQ/36nSM8mcATwnkYlpKnWBOCGZ5
NWXeH6+0YLcCzc4dD7+eqbVIJs6kmL0nH41rhYqYfVZnuk9CjLbVsTKPjI3BLCdekVfvM1JyVI0Q
d6gGBI1XTib61uzQhAtPpIqwNYblCnKxYudNuVtQkKIw71G395tbPr2XoJ+XTrRq6TzhVVA4GGnT
GUYsGt8+yG9AB95Pr0bu0cpnNZ/xDmBZvkegqseUdBxL6IjiVKPrhTBYfXowj4y25PGBU06lI3TA
tgNpKi7ZkVHwT+E8DAXfi0OdmRg7n/wna1HB7dU/RSu5kdCISNJRKHb4EsG9zJpZZm5VeTPfC+p1
CvBe1oK3y/dpNRatTSo/3UnqZbtMfK5GB0+lJnIV5AyNWuMqxLR25nUq97KUhvy+5MsEYetzI3DE
a7uRQT6sa0SgFVohpwrFMEsldXxOCzbZOw3nbLkxS1P+hUfiYSKKNvUzx+93SeJtYu0r7wWb2Usx
7rDKwYLAES70YuqHpJIWU1grRzX9SnE54soGqBi4PmCflGexIzlBPLFLLjsK16/FRK6h+GWIFTS3
Qv1M42liZ6CNmygrCG6oShijvTylXe4QX4MzOGVIT4/by4ebLhnCnVDv2SoSv8Dosm+8Eov3GxMb
P1FshdWBOSydQeW2MXW8i2faeWM+rFyY1DtAs8IYMHP5Mp9ESaxckm+JMBiNK8++32k4qOeTRwSw
JU5pUAgRAiE8tCmSnKXVfRdk83Wd2v+axc6lbHbS5MjhZ2euAR3ZjgondwNFgz8hnGrBI0i2VL9B
rEMtoNzHJ4fRi87PGvEAZeJJxzHV4SWE5WgzHJlDfUsJ/jX0DJl8eAtifBB7UB/WqG6R2wpbg5qC
7dtqq0R7jpZYsKgNDHxMs85J3Ag4imR0y8VweH/XvMQt1PuYvuE9igZvUMVwIrRlhiKuGhubRXSD
b8JG38wF9sxcDI1SQPDRrkGN5kqXx3dM1K2evbCyTb6pX3e1ecYWIeBBHepzCuLXhACI2rPToXGf
JpuY5kwewe3dV7sGzAKZ2w795vDtmCXsHuVCsHq4yExbV9DxF/C+B+TsOw09JMEdfsrTR6JL8xBg
1nXpz0n7q7rSdrLu3kyYYQHQh4I838r/bXBVooTs/Shz+HSMv+d2q7ARB2jQ3CwXmihzvj5xu4xT
M2Km235VKY8I0H8gzxVdvwGXot49otdqYEiVG6nEqhFWVJ73U1WomKvOg+K2exHpqAQrPgMI/nHW
vf0x/EcyecWTt0AUs8Rf3KoHlyZ/a5fJwBYoFrpViZEjK/F326KjSfi4dqGP48wsFHDbFbOg47WO
ibo3Iuo/V4QEGPen/Pr7o9FDCZ186r9M/+Cfp6ItQtW0WtlChYU14QV/e0o4Mo/ce7+izjlMhiYL
XY69AmYS6wgmpv+y4PNwDZX+Nv/vxO2xvJhd2U49Q+T+Yxk0NPg5TMS5eYHjK/D6i6B6AIO1QTg9
Et65hdPfkJaAwwDI07EVT5ikZqb7agwvDbwUsUYfH53QSCk5M6WDxf8WyibZjGeIyKjhHiufpcZp
lU+1+G+s2gm4wZqZ1+9QUbtDhfZAxLdUOSNxDe3bKRL3Oh0qk1W16srOiDiuDJ3h2Drm/wxqdhpI
3Fx3J7F4qrpHG+/ZNYTfsgJBXxtSD10kbMur9tgmz0uC4RQm5oDfWuSCLDNmRkQsgwiXliWj+PTl
lzzF4RCOJc3NALjN0unbF23SB2DN70N6fztmPLJGdUinal5Qja5CM8q4OWEyyyiSKXZt4YbeUM4k
WPF0zxoUMKYwq/TfAW1HBGOk5rSnTQOxndZtC6XpjR/8Mpz2+QpVeA1fpNkxK+Apuno50f0mIiED
FRFSxeDiCDYe4DfE96pjU4dPkELIQy+H7CSd4sPrNFACW3KinV5XNV7L+zGuVY1yxwTg4smRPpRO
KTgWlW2Ha57bQStdl1YdEdl+2DhpCbrubh+BqaC/04QV8EarBDSvGzWp9QR32tapvGPw4hIFXGU4
MN/foDOvl7CB3zjvdYukkmQmndrpJ+/dj2LP3nj6PT2ginwCTSTctiWcY0+3rdMWsPwXgTw0rwkW
/QqCHzKNANPvk0Pjsbo7UlfYOHwQAQbE0sDpoe2G3fZNn+PFu1s23ruxsN9VwjjcSMh5e9d+ADoW
mNu/dB/zFPX/RSO7i6im6v3CL7IsX2taaLUk42UJnStVi9SFCKi6iSUFnXGChIilont2GV1YIfYG
QEqC7RapFLmwlvbS2Oyt/viGWlyo/gUUbsyBi7gsJDODQ20cTfwfxs5smzWfE2PxDYeYmkE61Iil
wmrWZy6HVr6sQKdbNA3H1CJ8PmEp4n1RRS+HCzuwqfe8TPMxGAHaoyLyHxyylV+MMStK+/QJla8J
FpEiZEMSD083ODIIEiAvtyVM8WL60sORW8Lo5WQlVpyog+i1iZh01EzgE0dMwoobCqsY6p4sdt7V
LjyrCrjNd69beBCDNUIuTvetTts2/i6nrRNEKr0/+6Tw1Pdz27QjLY7S8tH3VjJwdx4U1iQOac1Z
Dd3eCHlRz/aQQ440XCW/dxrpQSx1FQqY7K//p+TqN//RxbYCrePEiIbtX3QPGVyY+JHM17f/QzrS
y27vUb5VNbzpjdcLFkhxbxFLDd4WmHwjvcBVcaksjvm5Mf4BYdn85iqnWCWKSMpljQSn3t3cjQqc
P8OTZ6jmx4QD5zzDamq04tBclGxHJ3a2WfAM3DRa1lKEistkoJ8ibIG2E7CanL4M68nVOEK0wuCM
GbRcf9Es2cKVJPR5G25wWBCrJDaSkrvG8cogpYvpgB0lQb/7/7M3NFzg/DgF5yXLynYNuevepowW
8w0woCVxhWGzjCUPvScsxnWm4Z6HzKdvZ0zGUAzYOPaYzEDq7NotVH4sdkof5dmk+Ns6Yn3Hh4As
t80elDw26s7jRhvjcQdtELkoACe352Dy9x5TYBHwlYDzt+HI7FjLnRcILfmMM3wYhq2NhvOCOdiy
QvpJOIJwzS3dNcNwWo7gQHgYqHz79quSReR5fmwj4F0mrVV42wkXm7/YyCm9UJ4GtMmyXlof4jEI
PhpvM9MyLl/NAewl/9I4h7gUaYnfVyc2os7cdOPO4016PAyjhgLAyrOleRp5syHk0Fg2qEzPNOwD
X4LBCO7MKVdCjsJG2OQ87YwWH6hl2Imk55eSiiinJ5R1bKqsyiELYikjK4EW9oezV0F8m8LJQc4R
1us4batcOqL6cZwGRxFmfcLRhllfg54+hBiAOS6kBrS/yn/eEj1QHfurYKaJvwQ7vzur0FP1NgRr
ja1zoKP4YFvfSY2l5EpR60jwWymQniEhe/OadiTvs80Br8qG/J5ZZvR6prQ6SjWOT2p7nZhSqGgz
nYQzpoLaV7r+s5PhU4aN+OXxw1MB7674VV9p3vjNzgFzHaR8DU7OTceZ0Y066i4WNQahpvMVYz0e
rC/cXZ/Z1HDycrF+bWBZiPXxTjuAwmM0l7pQtKUKRD2JZWCXve6TlLtdUATVEcj4xqQSknQYobXw
sO9YSHPbG33TlOrkJWglAy4PdQ2RLfRPuUheHNNyYEFe/60W2rfIQqSXHibbcKSnEanISJlNuxII
RDbdjHLdUl6JHZyQ4ZYdxsB9r9i8tF5UwZTTakN/ul+Hw9a6j+4tGA9hHqWqFJ8DIlN4f+LvYph0
lnuE09QSNMu6XBHI6ueUnS37bCUxbQHN5+KA7jVI83coADGhcC6LzKVx1g9tKlmnvMGytmWZN6Hg
5hjDrJP8SsG3nnS9x1OfVwgp1r35AMgtqJUvh2HMMzCzFPY7giIVhk3cwZ3D/8U4V1//WfDq+30Q
SjassHe2ZIT9j02gVlH1GUbkQ3I68w0/2Bk+NUNYeY3Ln4ETB8eNui1Vr/9EJV9ubAI1vwK/i+iC
CHREtQqMQbuUkxcAP8pMFcI4J/LYLEVF8HYlslZBQt0RUGl5lqH1tto3cCjUs75hLVn1mEe0VzwD
hnluPPpUQugSbfKP0IL4kmmMeKCGXs8PPOGdzufVQ461GvVGQLIPFMxn45najMXdIIwVxPXx27eJ
AuOlNoc/UibwOMBF6e4q/c1kRLofJENMqWQiPLdVOS4aWlE1xWSDYb4GjGr3tfdqFALMzhFSt6wx
KrKU+2bEZpiZtUrFuiHkFphJFOVDe/XV5UB4W4JwXnswrpL5uvICa6sBCUisiGLs4lCvyH6p5R4A
4MTqsf2gs1dVki6AfBl63JKfDpdf63qcpswwnDyak5JPgqSuDBRFVNkVzf61pBZ/R46Mp0Bgi/gI
yFQAdBDAAaLffr89JBkG41YsE2F8TxmoLUuCOHHbacZ5CFrsh0F4KB6L8IPyRmbFp1Du9B/A/4TI
KN4V+CnE96FczCqIFgvQ8jBuoFS+9GCzuKD67/1tvwgwklpdaRLNEdjVV0N6ZYY7dteSzxwq/mxV
M4sAI05pz2Wl+jGR5q7BVp1VPjpv9/QnuYQkwMT1bMaJbGzAV54TfhE6kTa3x1LhUmfcLawcWYIj
lJHU+AqkWdJHrVjD2az+s56vgDRWLCBz381/UdShonqMV5pTiW63e62tSwZi4Y5w+JzHcsahSI+n
eNU1y9FEJIQLf0o4lp5cZLfOVQweTtpwWkWxbIc+IFocKiEmRoKnXymsw23Nnbt6TO3fNVZ+61xN
YkVHrTu7OCRtYM+FsdDFZB2+8MVMxDiMnEvzZLVx8iu2gc+VzU/n5zHgHDDJdqxmH6MI3dcpBSd/
gBm4gN0EXBBpBBDYfQOY4TMSm+yIMkEDpxVjeTLwC8SQdk7pbgeqI464LN/e0fS5tmYx+P/lngxn
swom/BUiG2yhkDdk4w3pDxMAWrQ+KjAwfx5V7G+o5cTOTrBSASiqDiTX2zEtU7886QHwJfbLqx4w
ifQebji5Ak35oQUdag9hHvNFMdIbzr/+PaEgXXXPgAlK6ocU2osrunnOAS996O+1Paw2BCUsiSYu
IQZEVWw0wd2kM3GX3qiZayh2M3v6rIMpbws2a1nqskfvXWjauAZawYjBqoaZsKQbpTG8a9eRwPvk
NB2VEkqADdzv4m0tjW+3pmdm+4fa2rPpQmU360StxhqIQwOmQoYs0ecjpllyXYXHtIvqNcY5nUEW
xpuJALlUonWT3grbsgnSUZpoPEpqmVHUo/BzOlWMv7UKErIGEGren5UHPpVvgJ9psmL67P3Gtnb5
yGy+4IosGxDEMVhOZ0t/rzPnSTo015/GmnCbQLDcyX1mv/GHwBV7v7m62WAZuFzAy7k7FJOomp6C
r2edPJ0ILt0w3J5MWIgfnPBkE/C36sbla+dfUwFZ5Po9j50qbEtGyb1Zitxx5qej7bzKksStn0FE
rqUrsopvJGTFxUHJKO+9JIUc0o2Zd0gojnmV/XHmMcPq5TDJPg870tkGrGBL1M7a7+hiGm5Gv4WK
zXZ2Sa+D+FHeDluB9PFndLuC212Kk6uHvnHxGQkZxrldvk+pq5z3n5NPw+GPPF2MwgCTYr+QNsjx
lHTMrFDs5d19rurooizGnHrhD9Ze0uFLUJ8U3TPucdOasAezF1GEWJwx7+Zzpki/gHBO0doRvdk6
2NTqhzLusm1URVr9mcAPMENM5Guur+a8wUTlLgoEYhGC23lECUzKkkfnBMssqd479keUVLSA4GDM
m6krfj5YmF+JeIY+4QbFvYdy8mj/Azwig/1S1WtaEkr6JoK7p79V3G5orra20LKf3Pfx7AzqtbfI
XXabFwXDNCBshf4Dr4HyUL9Ds0M4fdJRs22rkOJp/Lfi+Y1QRnLCK5eWUjHzdSD9O+hG3zbWJ+dC
cxOVfq8HkIQ+GApAzDm+ejP8quGCUC5SWepzOuQhnJMCr5eLEZTVv9OWseOXR7L/7Ae/UF8PiqvX
8/7k71iyUijuEcPEQmo/2/+ZyBKhSFjQLOoppEk1jlsHmBZU3rPJT5InZUoFFBn6lEcJqRUU5lcf
3Fl30aKDRDVz9Eb9/kAJMM4/s2lbjofCO6455Jj3ZCTNWQfgoI4E4QPspJyZPYP5hsAsi/wiYcYs
YnAiuQjbnJPMt8argoOV/mzjLqN35KB4QDof9XZFVX+ZhMpfQb5kSU28AlLuhbJ/k4SJFDN9HLIa
CcVCcV5BbY3HqJKJmPBHm11KUQj+eH8Ydjblv/BlugRXe7oVpbB95WhX273Yz4h6th6ymc0q3gHI
KEzRquoNTtR/+ygcG4Z+1cF2oIBQkh8IOQKaGSyuVYdSNQWD6yTt/wYDi/yVf5PB9A3MzJFA1Fdc
lHfsF2eZJQQ6Vm442JatHEPs/4Hvk7e7qqFuvIO39yixwEpESZJ5VHAoGzObV2ckAqcpIhnYGqAo
kTlILLj9GDmbvvQMvm1Q4XArkXiRER5driu25Gn3/u+8WV7kgvlWkd8K5aF0z5rvtKLsj5qOR3uC
MYygJr96m+Rau5q82um1OwdtBuxoNVTZofj0gMNw7IX57IKFFB7eWBgUuQXMvLVEYMgZe+pL8BVh
wb13hZlrBaaYcJ802EsoQo9iRPEUicC+c/3FjYRrH9zAAxHeo1sDDXwM+27YHsKAJwugYqcKViWj
Zob4OZCKgIBcC78EIy/mhJ7hB9BEPAs6yfwZoRyLSPsBTk8fU9fZ2wMhn98zBNyBeY6RhOEdNNN+
QKiT+NMSuOKkAyALmzrJL5yOuloC64RYy1II+/DU4McfLq+PZ9WC8UehRvUmlJQ4OtlUDrby33W1
7XADBmpBzAPKPpkdeKkS3xEiFOBGBYpe9zQNQBS8yUOKIJGGi/RMvrHb6xGFHffVcUQtBfjUiNU9
4C1aL+ykJa9oAH8BP6jNa/aoVg1CS01JZfQfJAPHXXemZgt7AA9G8tEQ3CYNzlmJRk8uvBzfeGpO
elUle9/7zgzcXIB9pUOoCZe9kL/+xCS3GJees2N3AzESU8YjGDMisVcsXLsZYkJMb3uAVLu1DpTO
vIXVeIimclYY8g55HHBcziAH6Xy7gcOlQvKLuTr6GVeoX82rR+3CRk6GNBM6/OrZyuQX8keuLvtP
54DH6xl6adwQAxxYsLqa1PBOCUdh4XbtXEP00c2+QrbnBj510ye4mr+I/NDwXgVm/weqXw7L0l1R
NeH4hOt9r1iD533YGIT/L0aD73OV7iisfG/awYPpQ30Bw5QU1ecsy8nQbZQhuTCQgBs5ftdCkOhR
8lFBjsBSQwvFiNjW6WnKe2mfUz0AW9BGIrMiCahkdrGLhqvin5FMDXaRmonFED/cVA5fV0OrUs7y
2IJm2AVHG0B+s5v3Qf30i59vVXBgMoO4u+rngfKgZmKjN6QVZ8gpZQhTxOCPtdR20q9CZMGzjweA
Lyp8Plz7ncVFAST3dVMNlnuj35tupmTOISsi6G4SDTRGkEsu6bWPHb91XqV4e1gsu+Zj24eRGWlE
wuVoJnUGgem88tzCY/M1WkG1oYnW5E6ClkPhUDlEsk3QG91y7n4Ef+axhcvDUVFihK7ozx1JZ2sK
DcIAJNA4aCv6gZlJ36XwunBOIo9oj+govEG6v7scImR1+ip1Zx80qKzX7qYvvzPv+Tqzc0hksFiR
4v0Juu/eFgsPVE4JemvEuPc4Anq++lSrATzG5+maM4s1D822YxD1gqLHO7SMpwde7Cye/JEDRJOS
2hjPHhJT5+9URH7dBsRJkzFv+7Ip7C+FS1ZrxYoEi85Yj9SWiWVGjMbLCfwVaaVcPMbicKpoLk4O
AkX9yS38niu/DuRHgo3CMQVovl4/3ySxAxuecebFGpGiGd4cxZjldD+KSs0IpaxjrXD11s+N6umZ
htWp+U9Ufqd7HQ/K8JTmBpbp9x5eYTl2AdTleiyHnSkTgqOwktmhb1a7+2WSNs98RcCSElwccUvv
0LkSB5XC7bUR60dpaa48lENBgCWoYzW00Ct/KCJxQTggMWjYjbI0BR4M8MQb3O/kRqrgj5FF3jGp
IG283gKbYUwaSuep5EhjfkE4iWT2nsVsx1ohXqFJPts0ohMYyS2ZlusJP3nb3X0cRxSHJDedSeMS
2Lfi5X/p9QZ+lIEpEOwnV4MedBQVrAFrRi7IP4B1a2RvQHm0GEAte5d/7ff8YoI8PsiBWkhReXxt
t9EKtPZk2reMmLjNEmcsyyb/n1HlXqdftVMDzdCNrg00v/Auo0tBnCIjKFEknVqQBfeTPx0S+O8I
J62iik+61//WAZKWguoZm+cM9U6x9MuKOnA+WQADCK36FSwc798r4W5IkQTfgSWxgPWos5XaYSPz
Xf70tWvcbaqSQdweKjwmyvWSU5aZ5LAL8YfK4arGhUCcqmy3UwkJhxltPKwXF+fr06nhH7XC+hF5
lIS7L/+0oeUF88mPSJAJGutDFjJI7OswJR4f+IpjMtY1lzvnf4O4anc60n+0Nv2dFVw9ljRX2Ki9
5vzgoFXiB25KYzQyQlG/+UePl4+t0CKrOK7Lrwo6zTXKIcYT5VoJhLkpsCVLdDynMkN2L8Nr+94A
ZegzhmkrmQNr1697DRCl5lT3WCVEOAD9C/mMJmVHEPRWAbo33j9s1IkOuXm7x6o/64uvQMo4v2J3
KDr9qdq9tFmRNQZtp4aEikRhXqVl1ieiz9xFlU7vihOMsZu50YVakGx5d7kYa5ORrt2KiIQ3DAhB
1bbiVhl+MBS57pvCq8DRSAiKlYvJMeDslPH0oJc7RHd4yKZr2fgQRY1Xto9CnIVOY0jC736jzgqf
j0aYPzvZEYH5p5GpD6gx7OT9ik4StqF3TLf/pXqSsPup9NQ17hjlXTvkFls/u1gv/pwq+RmRVxcx
XBOJvsZIOWlDiCb6uQZSJE5kCCLQsCNTkkf/qfnWB48wkTAyDbnuj5Ey3jKfuqy+rHbYw+7y1ERY
eXadzZTk1DCNhR6ASnGPY8kjP7k9k4ZMPOwu7fxdrxclgWUC3C77qzvmALFi8HuG9VAXTZIxjTSe
m4u5FXhIxynXY/7rWQLS6OKd14HnMjtSSJMXq6oCdxlMSBbMCG/Uv5zDqD82XfVdtGPoU/AjxQC4
TiAGqshQbJZ5Obk2sX9/y9Jv0LZWTzjIC9q4dDFT/55t9o/4uy5y/W5zS1Cb2UxiKf8CsQb1cX2u
aFzx9HTkV9G4C3QU3K9WNaZMg6S5yk5pjhyzX8L0qAt9TL2TAotP3hO5BaLFH3V5yys1gwoYVa74
ykUCVPt8B4OAQqrBPzGHz5QthgOuCS5BynazIgdIdenYA+V6jV9jbo3cnFfFi6+wjPYIqaueDQK6
y5ZYumfH3hZY/2fZvx0Pp4p8M9Ya/ud2dG1e0Nch6c2Jqc3TC4yQk7LTPsudsgCXlZoGiUCHTF+E
X2Qq/r4+t+M7ihLPEvdKwB/DCOQYArFSntwRsUk2NFl9FHYoSCdnw64EaVU3kpyJYdk8wXc2jn/e
Cx7MTxh17LG5R9p+H2uAu5Dy2phwc78f3ekwdJh5xWqE06uv+w3AUPUhFyC238OgJsQTyGWj6ZzH
7xqbR+hVzFioyw1KFCRtzJAdQ7KmVkZEUQ93TFjy0OiHQlFcmRZ5oYS+9c2ZA3+wzHYpqS7b/hrg
XiEM1nfxNNtKpACIwmUNM8WvSIXOAKkRaeKh1Y+YzYljTkM7b4hZZPXzLyx3GxCKU9ieTJqcMylk
OIGUKy2AZejm4yfCjJntHirZVVN4atPdoFwF1FB7vUM/AXn+zBOVGnE7/6Y+3Bk8CGroqRgyypvz
BXyfUBYJlBKWCTlxo2Mx9GoRUIO6uk7QBUu9u3wej2GMvisvSeVl3n6+nhTbjyYbn9YccF2S1iSD
XkCPQxQckuM7wshCvyanmCXWD7C3aCtimCrwawvYOr1r9CisluxXJenubNL/QGbyoK+3Tqz3o/q1
tXyrv24nN9BFgkzgnOBaNhYxgZQ2ZxLTDWL+hyoLFBn9Uc3f5pTMzX6iJ7TwToqfZKZjH50+IfIZ
/iKxLYMXHW1dAV6nbXdPhV2l9XaC+zwCKihWfoZbJD+2uaJcjAQrItBiI2UQGOVS2UEobEY4ekzX
MbnmKNjrjhjDiVQ7nbGqTJvBUU74Abcl1DJDjCn1+Oop77l46EfKB5NRTMPQKwubC/+q97bDa3Oa
G0cVuORy35BKzQi5tmILsNv1PdjtzWTNSDHKpDVbQzpo2t5GVFlkvJ574waBLIifpBST1uHH19OQ
LG0wwTq5bqNxy6wnCwz3qO11pStryJs6oo1TWAFkfMKFSO3NTgutyI04ZsZDjL6gVXcdGzr0VhOe
c4lBtjyECWGNx1H3p9SOv+kSn7+hpwETFvOO4OUe3ub3wbFgywbP9pV9AWRZ65DOa0/FyHXMdsZO
7kVhTO6xkK1ZLFO8xID+KdX9Z5ZtlipBNe5K6HzUEsGgmILz3IXfgyrH43XtkXSmo5yfBaNkNo/u
XcQzsBJdhGtmMhbiG/frDdG8KDHUP0r/NLzxwW7oSu9+4rvshHzBxjfn+E2N3/5sZAc/Jn0dldPJ
df7Q9h8npCF/utbnUM0ohRAd3ELXw4pPKdInABplDzirwnn/d54bG9THaVHm0nuklO+H6FtZYJWf
Wg7ymHxmV4QFBTSoKt1MLGIgrLU5GSMHtNcpF3O4sFEaDoCAOFflXCnUBnlj2fSVRyissbecQ9BX
kRdDnOx18Pse7y9Dca3Qr30/1UyKpeew1og3EtDi3NvjglGEGqYkpDPZhpSu95NkShA1N1pE2elq
Ayo3mBfTH9AEQTcVYI+3SDwvSjvLWbLdaKw7m3Rpm1gecutsNkcyVKgOIZTXbp5G5a3hDDJjeIS7
QdELKZhmieXWtVLOYWY7PfQZTjLCBS5haXIZxbPlI5cXT1Shew9ulrIF0wwolhhm4A0SrZB9/El9
NC+836x1kwVITvueGSgioefTj9Kap/q+8iYUiXG9tme9aposcebQE44UiFfEedYPN4uEnIlO+8H9
uXLRNvHBa/H/KJxgWNNIGEYELNWaGeP8PDTWVZlVCQlaXCL2HtQWFDvAZeIN3+ANzQqfPWeoV4rz
UfY9oLogqkCyu44JjOoAAMv+FYkGFyzppSpTfncEWlzvwalrw/ri+gKljtqCSd4IWRdx2QQux5Ja
sacf+s97p+6eQwXPpviEoNNC/5bU6VJCCOpF7vfJxpASdixNKFeE1Nfnl1heQGPf+3MjpZyq8jcN
AGlkc8npjbqfX9ewbDZJGhR4NWPxJQLP6wuM7gQhBYhsCs10qI2vDZF+ks+xuQgKylWFVuDE4TfJ
ck+t3j2hx3PXxNWZqU2j1tzC2zFv3zKn9OWSzTg09IfhmC1kbaMFIN4TZX2cYozL9UyWJ5ug+L4X
u+jw8gOLSBteacN7V8zIkVUAF94a5WabnoFfAOTioqbIRGdu/bscYZe6sa6o5hl51tKnPbFZgx8V
zFjd+eDHZO6M6XFS8SK/vy3+YnQc8y2fOFxdbWUMNc9/l3zUEfLtYBrAs0IHiYUgxLS6oYiBCbbM
2Ro5B+64MQHFJcMnA7bH40dYpZKt1EfE0aaJpeDOrkp3fJibxyH0xfDdJQhSVrFECcp9W27Ty++k
26kobaENxT/lcE2g4MocJZVsisO97u5Ha/dVsbY9UtZF4lRJjlmGZRRNJZjUO2ZvmhdZe90pMZoD
fPkeYFLqAr9qXpS+8CgwVdrVIDLSPx4dgpYKOns8N1cayZz+BE1UvF5PH9Gsfddae2iFoug1EigF
ZjLLn/LSRtOUU6xUCskEvqNLCr7lZ8FeoOutGHDBoquQDYD3EStlOWx98yrJibh/UWx67ihNKI9L
wrd8eeWgotg/jUzWwYW/ytajNT7TuAvrDTaV78F9cX9syA1uOEE/CYN5JrDnLq8wNkCJsLiL65d8
LIyvDoB1QDNOdt/n3jcuv4tG0wMa3DzwIYQWeX4xYEbl/nUYpTyoIalYEZXaV/ptEIlhQAt+gHYT
LZlQkL7YsxkBlEnsyHMR5qGPolyoWe/guYVFLsKgNxP8hdiTCm/5g5RN4n+0ghzOa6DWns2CbKUs
ceH6NxicK6EUMAXLiqFyEMixQTKO6vxKE4h5xFmq/qAmsP7KF7aY16ytjOBkVyx9ulFUw5SF0LmD
7eceo4im6h4myxjrLXI9Fd4ZJQdpwlK90dSRtod1B9SYbbY+5VuNdavRDpKZCFuX7bwjdGq00MM+
Y1eK9PqHlyTKykYk48rIw2wVD+zG5aMQJGMrpDiWQNVfjRMVlE6resB8ITbCK04y9mBoPKdqfCzT
GhlLSDjdT5arJ30950TUNv5ljwNR2MRQbWlBYFaShy7jD/+8XtrtYG07TiWM1VMqGkYoEsigLBmQ
Ok39C8gWQF3+adYHz1zL8U8/i5luL9bsiszHOez8zwjcWWJqnbiPKHGof/JLcetCbqXV78E4+qQr
BL52AAN4zfItwu5xx4fDLWuVzaU1nXId2cM4MHaJbEbpZO1eFCLXxX3p4T2JFOr0A1xuP6EL3XXd
XNPDM9EG3NZFfthpI8baImMJa/7rjmxtQYLmTqXsZYghZuuiESJLSZwipAeIhEy4TjEDAOu3Zip5
jaYLBq0OLQgspsur3ltU0Xncr/NKmDmfJHDVa8rrkklnP6RW3hTWqUlI+IUtgkHw2bJbTN+CY5HO
kn4NjwZEJX44ETrrfkveVmBxWJvpQjM4UqCqyB06pfPcukr5gKoRgZcWMjXeu+fPO1rvGHheICwG
9bjC/v6iv+pTgu2Cnhp2SNGRhjeDC9l5ruDDhfLagdScrJfm0jU9fejaylzoeBrIEg6Uulj27OFA
44f/npPEF2npKbuHjrNwGCHEfynnG4muLovgx4d2tjTnXwg8kDfKubioyavI2NfFiU501fgD0BXO
FvV3IZeMBF++s6LB7bErkBhhY2bHFb4UxJM1B11fVV+sTpjzWmP/UO5XK4m4xU32PoNsULQi1+Hm
rypJCjhmsVYSBzZlwjMkmP6VElX+QxElvshI2+wys8rczTYagIvBjWGcyvND/Hm6GruJHAze/Bf6
sD4JtPcWvhJvnER1Z+ZK2+Z5BcT8JM8VWdHRwSNevRpGq4hH+UEmPobP2GTSZWUUl8Cu30hArbcT
qcwa6Z1uyq8AjCQ3CjH5u3HNqxXOAU+XVYCTgF0Swig9sHJyw/s5J3dnQUedipWrFhBAA6ngL+G9
VueuOJZlJfNm1hWosOXznxJDf8DVhO26Yy/XagW+/TtcsaPWtl0PAenDcPk6UN/PMwphjY6mV1sg
mVkWpGYHgo89Ugw9xcTQF1UvL5h0cCVBnHVMFYm016yg7sn0DY4Q8H9cteZa21VHXWtKlq6i0YNt
iBa+3PxRwKvrZV46QJ1GVXyffJHFZMvJ6UBnzPm25USC4kQzCnyB6l/JkJdcpt/zPa2hIq9U1wnF
kjFCGqvB5NcC8qiLUKWCSgUUd4T9MdO7tlaVKjOvL9o1lKo/yGM6RzdQLCzWB14WYLu7W3p354eS
oFE7Ud/mKFa8jZrvg+ZQVY+LB+dnZUAItRcJgix+dx6cpnN5ra0FUCoxHmObPZGtuE/mj40G/wkA
oabzphHwsl14qAFyIhwgoGhjjAR0iVUPA86iFjBaPj1wjbMwGbV27DvZGeZgv1LVR3rB94jrPIXH
iWxh4Gh54Idk1ab6ZDQWcprl7HTAmAtlm3iyZQAbR8YhlmxN+7dxywjM2qBnnOvJ2j1l3jHKIviZ
ILWDmOfKQbswe0dCK+s+2ZCBPQTy1lYg0aKWYt9UsXYGyKjdaob/zRxS/e7VCG1+sZ3kSh9gROcR
m2LMVGlovubzOkVB/VzqhFOICr8WJtHvNa12BhnU2lqWIHobF5U4nHt52h4FLPH0uY0g+0H/sCms
rsHG1BSeyGedd07ct7TLKXrwgcaavZ+/9mElUWKKHqoRpt3+14iJ8WywXCHyoYk91kBfLRmQdZ89
3rc62jjOJUMaqCmcEjCi7/sgxcxJzFENB0tBPWtBUDSojXi+KrPNxbdg9IOEkQUlgD6dy8luFciZ
ifdqQ590V2N2yqoFbVSkZY+OXFBvWbCYr5r468zSrzxILe9/ewl+QfPA8LV6M9FIB0VpXi6M1u7n
AKw+JLK6MZh9ckzDyVkuBVhtFxLfCuD82Zfc6+PN2LEey9UMnes1HAptcKCD7obS3lR0RyyYConI
6ii2B5ouqx5BkABrFQLhvW3v4F0POlewcAOAYX5fgReJQOft/gFf9l1R/3Jro+sFG1DGZh01HnMb
GGc9oYObQ+JJT+PohZcDEe8HN1wOfjf7YWe4sVA4B5mAv86dnUSZ9rBOcztux7EobcWdPiTqjJa8
Byt7SR/HaEPprvk6ks5WyMtg4EPXPhx3RzOoBOE1vnYMpiC2q6PUaIWM6Icoo09EDTZui12HnKgk
kUA0xIYNQjFIwaamUwd622O0dJmhSHd6phOWsf0FTJOvA9hOpK+/wJFBnAklCOmchHibdd6GbS+K
DzBXDF9OlmTq9rlvMCZ5UtqL3/pmgh8/cnSWyNdrMG4mxPLsZ2XtuZWlqtCWrnuA3VBcHv/7MXkV
o1mUN13ANNRNLd1hA3neJ7qp+VhZzBbjx8tK6cq5MUEE9WLfRZ5x4QbJD+nxqCNf4Q1xi15w2cg4
SWtXk8T/I4lASxObXqesJ3bsoprYR8pxSWM0uYnvUgTNSUcmPh1P4Yd1d+SzzPok1hUE0geEoayl
BVEehv8YE8I6GAsLZqacuFEFXhJNvyUZK/7WCl7ELO7UMPRCXskmr7Keio0yIjpGUGWJKc+KEW9Y
A2Wj7wJsOrn8wZqHsMQMWEmh/3B1TvkoS5mfysboNkMWpaaxY4hNZoLi4wrb+CRyNhmQBSXEQ7k/
UH4gojIKXOAxTXG4wrRLYQm+k84QZ8YGUILYnNHhyqc1ijmcf341oOL78Do9V+3GRu4xVZx02C15
WvwWTam912sXjPdpJcubEZfub0QD5x4dVos+2OLVJ9K7VH6S055lJu3sIB+OFLhIVJcdGKldv09z
kZ2Q6Jt51TDcZNAz1FaR7C+8j605Vdc0xwYIsFq6v9HJeWa6OI8JO8cYFYJRKWjo+4p8cMylVZxe
JjLV8aHodvDHLn962lsfATqOr+SOof1wQlO3WW10RHMqA1DICyJLfhhwyjupbX4YTFVcqRGtFiXD
LTVKAsLTBmgrtV8qRGUvfgMhBo1R+nokD7qmKSCMTegnD35nqlrGQ7isT1G9xjBGhZgbj817K03O
ul/9GYIwLEvwL4NTMLleMaZByLTq1wcROx10htbQW7J2XzMz33+WZTfWNR7Z1UdysfqLJgCUlHr7
ve78VjDwrmFvtvvVvPXUKPg/DlEISjsoiZ5Et2wwuYLBYx86x3DHMDVusOyqYjk1fhQoMHLW/QM8
XtR0P+PKaC3uHLQE6gC2QWGI4eFsEHssdfE1OvgJdxamQGlqLXF8Shr3fT1yrMMOYcgelpj5nZyM
8r8tetFoDXnnTKziIz03QxRznYFjjwoKxJs49q0CVyNgBiMhQ4EmAdNA7iOxty958IybJHPMS91G
xpKs0dryUGkPJpyK2mzKDAYY9zilomRpImfVZ7zOR7/YrNNIN50IvUKqwjvsJX/fb3hgQsDkcGtW
B7SRlJ3kbBsICP8YUruGRbzYnq7GHqoqDR90tlEyuv9UkTVe8v2ZzWe2Wp7Pigd8g0D6bYXlJYF0
OfldDCdWmfcbfK7rNLtTSsm6LzAmSe5o9ws8SCuJJTQR3daMkqxl0JTFAQKaNp0PrYx1AdKMEqC+
5qj0j1NPlu3YyhhzLFISnEM5MYjkWiHA5hFxmzVP2t6LwFPbbsQzqXXUFKJemZc+rn93eH8CsK0z
ptfScqhPct8MVo0DQhqqAgDdjgcWJnXj7Rrywffgtl+K3CFI5aNlWzR/M9SWNkmljZm37ly/VsrO
26QiA9VAUF1SP64FfXupGhq6tqTXfqebT4P4gfS1rze1dHrQTgxTXst6oaks3M5wuTY6IGyWpdMI
ZfuSTjQLJ7jtXnPaLB2CsF2QlQvYMG916KBpswzGtlEiaFQJJnmcow/Ae0wp3UiL9INehj+U8Lf/
oqA20yuIS1EpVvkgFOmkyuNzB/meWlMqEKUEE06K0mFx8FrQgbwkjYR1diOGn8NGm6GxfVJAIFep
OL4sc6mxahh0A0rk1ISE1XsDAhLqZhJof2YXjWQB9vsolQE7WTQ5mogTfQrGJpbacUcozO4j+qSE
UapQmGgqwz3XtOxPhENxHjV3amF5p8dIbfDH7enGnsLWJ/K4ptS3tpqoafUTcqQXiseju0tcOCju
xl0OLagmCdt2u0KbSI1gT3uvwdRxDLvv4beIkB0BO6xFnwybctlXXZqtkkDmSeVwFN8JTctP9nBc
tzNFw20O/AvTMzoFGNAL73ItKJ8w5ywEUS5HsgzugzF6UVzs1Dk5/NwwFzehPD3gRgQsR7YOZMtv
lAp3vSShTd93eB2rLmViG4JDMv3HXj29JjhsrvpPmEkItBBzgeI9g+E1qetmIlM6FIp53yb6I1kB
CwnQZGLot779N2jg/H6IG6xCtQ17sB27yo1OeG72yUFrxh6qqu4kogd3Ir0tmPsSQueGLmhhSwWe
zjkdUarEE44gg0hNlcYz31kcqIKBpDgTRys6VdMpMbWlqkZr/93CLnSLsujclYmidNr9/KB5ettQ
qyTL29J52TNfr2QOTy3zcMK7xKVfdYm3InrCJb/KD6ZpBprKwKYjnLedCXXd1WMTEZlEY4Wv3/RS
/NTpWQM0BNW5F0TH8+JRQs8sD/BvSWwJvhKJwGGTOcwE1nle7Ni/RZTYvVhvp9VZNbV1AiNcJQIG
4MqdQXLq6PqCRc50/SgeH4u/GWT8LeAPTB2IdcP++/YgZ6z9TVa5Iuh3wRT/PhAk/tDiXGRVcL/m
xuV46j6uXKGvxDaFCR1UPDZgKQOG5rkjkZ7ZjBxtYe/mthdM7CIi2TbWhNy7jBEg23yK1OGry/kh
NNV4SLBU7ndQb/V7BBdg5tH70ppUP84LQnAJe1boBvj3DeUOemY3iSNXOqezhAEIAeHY5AkA+O5A
L8UmAfebuU12WnF2IiKNTH9RrimFB1x1A55jAC2Eb4uSgWopT3Qj+3N7U4M4UxtRD0tunft0Zwee
N9Do35gKExmV5DwJ/OsEZzqC/O/sg6OwagOnQ9jDUJXlc+n6g/4cOZo/mUsK86XmUlT7CQUAH49Y
7gRAJg1091AEz8v0j1U9zOKEWhva/UnOgu6wNzzZlRv4Vf/rPtu3ASg5+u7WQRTJ2UVbNMPQC+MZ
pcPSnmj7+ihMN/EjgoK2Q77kycfMso9c3J2V95cT39OaZHeWc9xcap3gt10STuYAbwBsN8Tf07cD
djfmfKPs41fYidfm9OoAOdazU1yjfDRitR0Nj81QuSlvu5jic/9kaZBgDNpfsMIUB14A+FyYZirf
lRivA+Sd4yTLfpa2m0USIsgl8u/fKvq7/curwjsEOR/jgbZbNMfJ2wStYQ3mK9idBKhTAfSIoxk5
obZmNcRjcm2LZOZrnU8Z4MNDFgBUerugCfP3EynJ1iI0AdJcWuk/zD58oDtavA5XIFSIRf6TtzpK
wMafvT7go/I8q+C/ZFgUG9ME3uk9nh3V8JAIiyghVi0aURnTLnARR3BZsGoDMzSrVEdptY5m6Ml5
o9eLsE4JWZ8aFFoKKJUSdag3B9gviHmec42X9OBpMCAZQQYl0hq2BSq+3mYKfRK5nV3sa4SOBDL0
Xe9zw/SKaTzbHsHsKomiw4bAxKCwMcNJeMgeJBrK7E1898wS1IVamx9gusW4K9Nbt56YwThD8rlM
I0yNRcdzqZ1tKzTSBCAx3tHfOdqYNLQCOGQ6OKIuVBm1FUK2CMLULVkp78ZI92DXZ1o9iSGHZpJ7
b9G3pnnHkgVeURC5or9e/PXjwSa6X2r1GpvYOtxSy1HLs2VbXyuilPBQ+AahZniFgxy8LsuMJ9E4
QkTibVzRFZm17UBDd2FjyfMQ11nEFkrEdES/dbqSs906ONQSZNtMnuYcqjWY8XRpufXvbpDGnmOJ
7zIlDNUdhkF6hWFSxyTXWG36j9Hvm2bBhLUXxjCBvRa3zoIyjHiNerXHmvwfya8tu58qZcEYFeK5
XUmVx4bm/5rI+yANMuer+nyIcryISbkQH7Gwmqc6EdGbbAe+FKp6Wy7Y8/+3rdNDeT+CtdPeqxvN
vPWwPhQ7trTg1ZVjRHruO9+3/ERGvwKJxla4xcX3P1x28/lhRJtdUGVYpdwkHUn4KZHBoswLfzft
exQYwduhJ+IMaH2+i8eUbSanLobaHKNjno9G9hMmZ05cCalQ4hCspXMvRUbJqJ79Ajucb3Ov6h1d
3dfe8X7HVryb907WM+4+PqvaFxZ/PyqXnwuYwQ7CAsePiSAf/+2V+wrW6owVomYwJBQZvdlEk+Mg
dN2k3GGuaMounSTryVABKShnXPziqGAByfgffZkMJLLBGIFnf5bOA3XT7XH4nQLVwosreG1CY1qU
Hs1oxF9VsNPA8rKbzD5Kh2WpXZA3zZZW/CXpFwwxhIrNLJKLSuwtAG7j644v2R0xbRaEchVHzBDc
OgWi3wEfMnIxwMAGIGiAZmsAK0HTdJw5wCdAPpVc0QpNPD2EvVEEdCrVa3jvcYm/zfTxb/Ao20sc
zxxVDznFa9sCQb4HyULSEf/SYGDeLwpHMX802GVTjpx0vcgV1MQmLPPy8kcaRPIKNLjrbOexi9U2
RoT+FMp4pBaNG6br+Gzx42MkRlNNh51WOLsB3KFEoproHophezOeNhiitC6PO0SvPg+oCrYqngml
lq48kybI5jVSZ8w78iIhD/MelXVcDGCZM2SXi4847Dkkx6+GCual4RGhWW9qE7yrwsI0LaEwU8AT
IABQ97Zyf/d4KSxo/wwctvJCLJTPibiyzk0AAazMQlbgzu0Oa8gsByfE0QDl2gzb8sQ6Jr4n2dBV
2gA23R2vDGzAo4PhnbH5axQvCYV34sNNSP4zmLkysF5p7Ph1X37Z4dsH0F98SKm1IsmQ6a7u+QpW
5Pj0OJJWbYEylPUJVPGNfKCo7U3egl0by5FLApw93Mh5w0c7h8X5F7ZWO8LODNQN41FfU0A6pOrB
yOMUOwzR5gzSYySrL06yA2Ia5bGe6RYQiV/FCh1uRMDyD2Cqj9Dp9OFO1yZA4+l2qDCbnZ478K9x
TW5g7W4y63RTt2zkAjW7UDojEoYgbwBQizBdWn10sw5cqvyQJI+DDNegivIatjMBcH1hm9jO806s
RVArId/XJyJHpPqpUGv9GTIrPZwR81kxD5mEHaPFUEPEja61KUcqpW0oiJLDzhxLF9yTKiJgeL19
9jkh5lhLj+WjqutIZazBafUlIxaN0yDAoWj+QAQCMI1ojiTHzyCksjMr3n8TEbcz5sLCBR63+bpR
6aj6Y0pNHNZJuzZfSNJxHQ58XtK/5DVgY70FaLdffT48NXyAQ1X6HP6Mf9fpmLfhJBBfZwJmuQPp
jzpBgDizs+LAhtX4Dt+TXToZeWe40lvYPDPDR0ogfYHxvRTOejVnIKM9r7Xj/t9xuAEQvVjt+tcy
90KKjg3t9z2kjgF1oYjxfBgkYkHOtKpHOB8T83Sc+yFuVSglxYBU9Du1vttzzuVamd0C8zBSZXtZ
wK2hdrIaRUu/Qi9hoOR4UwIzLc3yaam81X3GbaT4gBiXMrdkvoIaOz40VeltuZUNOu4o9qMWBsW7
/iYiZerBsFPlJAGT+dzNK9vt9xdMeUkZiluma1RQ3Nr/l26qTiXxWZEq29RJzGK2DlNoscEEVf4K
BRuMUMvqSIFoV4tNb3fxOrSWaSoV1F8EFammbbqdvR1/IoD29++dnvPII/vFHbzMoJKc1V4Y8Py7
6wUSlQ+lhuaqo0Yj8vW6t8aHatOhcg0dwjbn4FoWFVexFjPTSpJK/NisLtE332g3D0R6RbVHT6pJ
D0NUA/HbmJuwGHq6AU+KkT4NvdQiyAoibg1iCcmHRXYEJ7kHRJy+nkPw+OPshBda3pcGm1rLQHcI
DE/X3wh73brYJbLc5eP2lTbdPvfSGQunozgv3TBG+kpBAAoQLyDiB9y731k2Bj43F5zbOYtBxaGD
k8N8qTQUW5V0jx9MXCb7k+Bcg0utAWRjFpqbnWuxjJh0576QXHD/k/3KBzuBsMrLsHMshmXZYBi4
IjnBAqZeACDXZlcYFGnqCHvxVkXgaxudBZKJ3H3Vf0u0qQ4mAM5ZYE5s+Iv/4OT0taysu3zjRw0e
5kI9kCSYnutg1YSa+qTX2YX6E3jgVjKb+9X3aTpRwzImpOfkSYdvbjfRuWlEdGPyWVjA+9GV2nkl
bfq17+yCoeBFIWubKmaXtRf2mN86AQveFEbcXqyUAanzhd9HKXoI0WcfQyfSI9pcvdddsRxrdeak
Dvr7fbegCEVAIJWsfKmYxrTkbkBJJJtdQ1/KDCvuPSoaZDKvuK0Th61apnjw22bt9iM23wvlARH/
Kx+gwLdPMgKgsHOQkXVG9WquPR54FQejwtalp16Z3pyqQ7+ILaSozYjRrAreeCvfOt7HTp/1jP1h
cst0BwTGJzoUkD0wr6HcTza/dzT8ZMB/PSvbEqVmT2Gg6jrsKWN40vXeLQHwn8dXp07zhRVh4zsy
2fSsTzrxp42bKoOhmlGzOjUmvxCsdSgOI/6cRDRcMdbpoeIA/VFtNSBYc6qEgS78u/Gm5Sa+X5ff
wnWp7cO/BWUp87KBw8c75bFw/XPHBTkBMoi/NemVYKSxgjldV2zJrQMNgZLawbMApWZi6pcQcmpj
imA0/rOaFlfmmTYizg3mi3IEdPJYbajzFAI93bQq+ayXEFjvWGRvH2rbcLjgBuJcPCPqDrsXJc86
D3xeOQ4RlMuaNwyBKj/uFT7t2mX3sjZAyAl5naZ0ZFt4JZ5EZpF6ZlKUDqwf3Yga0iVVIHOo3nWA
DSXbLu5u+9yyDRUaAzK8hquosP2sbkRf6voWjiSl0Q4hA6M9iWhR4iylj2vXqRX9fxcQipBRPVbK
bpVut8D/xHnHWD7niGYxL0mE4c19Ucrs5SVDLlw9ADM6E7mFR4V8IGvvl4WQ78aqFTYsmIEi53vf
vK385wZ62R7xUXvwNnnixvaDFR0zCRKjHr+J0C7SdPDmFIDF1Zin24GN4rl8Ek29Z5TiObByhLII
+dhc3aFcMdESudP59Wa9wn4vVL38rRFshLmz1rt1rRyV1RrZJAoFKf48OP6e6yDMPXILVeVHZRyr
lyxVdHEfOiXBSXk++bEAPPLVF3XVYQ10Gof+pop/iGSSzxqNjGMgywsdjdnWb4nkOfwfDg244wWl
HU4KhT89n91ylnLmPuRM0n1aYjkVveMl7dB5F/Pc3OSQ5DS3nKnkRkTX8eyBJxyecBik1OGo/S37
7DuYIi3uRzxt2sMfzTVvn3D2dAwYqVe549sfhK5GmjC9YCRrt3DSyf3fMf/qrodClcoedwfApHkM
pJ1A3eFcCf4GZNRtokC4w+9/Lr5dIp4h9IJ0Is9Ck/+xJUVMchgsMBgkC8RP0cpAZQqt3wJdeG7j
IpGR8WSF7+kGncYzVP/DeAz4dYhqWjHsMOwnXaRqaUuU1Pe0yWkRlNvOBcX1AUokB5dcmNDInK7l
TDUu8Au0jjSzt4l22ygy+F7PWEGaabqB+QUR9OiF2rF+2SlO/u+oNlVNZtKAZz7aHLLZFamlVMTR
0nrvpPpFcq+JMXFAOK44XubNFj5FX/D0BYkzlCHrbzEvxB3XlABXoiwwhyYp5da77RccvxcABUnz
MduqIKsx1xhYMqfxfqL9rQA8mOfZVTCQr39mXh0Jjb1QV9k6DX3DT0DJNGfw1R2pSiLvqNgl3mkR
YCcnqhHYYbyvZ9Vc3v+HsKIT2UGPM7EfiE8bZcek2k9O2qv2uahX/h/8ItK7fssm/z21328Im7Tg
4/I8cZg/ZVZq0wQ9f4HW8DJPdLC5Q+tJ1O13E+wsXtArJppF1HfPKuT9Y6F5nHAUhtqSg55KENG+
iHBqhOpSBVzt7gCb3D6MBTx6fcKEsYXwF6buoKYuyxvU8dSmgdG80cKO7xK1MSM6zjkTNKMzAQBZ
eeQYijyMM1eRkxq+R3EwLcObvLYW28u1oeD/2EIhPVjrAVtCJwEv2dNfYNfwaqromMd1oLBdm3oj
bxf6DS5VawoFxfZ+JNPLFsoNOY/x1yBSDuDlhRvXkY0gi+fm0cKRQRfhMaDteQXD3Y9QWnkj6rSV
nU4zcufnPUKzq85e21EGfZZq/u/mHbExlLZW7PWpSo/qBCKxIRKDryf05gqU6WEOAMdnVhGQYMHG
RGrercpriqNtGUzeyDRn/LBcV7ZBp6jwe7uAXMBg1/w1q6YS9v3a+1pWtp7fOhs0yoyavTIVfo6C
URKQP0OsrCUp77bKy1gyxZj2S4MP2Qc2H1CLBy7z3qHeFgi5c9X3+8K52JbALdOaaDG1N+lEBzQP
3OsOdOqJdxebsefmMCcHK/bKDmuKcl4igr84yre8bgrO7WP6wTDfnQRShAnjlmnup55yywPnIG0C
cRfRzVGgEy+nDHFGNf+l23EmDgQ08MR2N0BKQrIqXNKoiM88xAwKorQDNYPPkeiA8tym2PhTNHmh
UboTZNZnyXlzMyeovnsF7Uw+2kkya7WUZDqzOlbxVlmJ1JGSEo+A4QFdTA2WYIJQcTQwsd0olohp
hau085BHa7rJzVA+IHSXHd3DapCrvQ8dcqkAYhQ+Sx6SD4kT/wGyHdXVOc60v3orMffmqT1iaRt+
wesRjeIeZPVd+LiorQ828CRX2r9EI5U7hMSpt5160nrDcbopzQ4+87MLbmdUfLncrfFVjotsR3T6
eHG0jeKfRHhoJ+WdNvm/9HqlUNIo/RSKG6wqTg4rBiqOo+c3MmSV1rqxXrICole5R4CxhTkxeuVD
DlslIB96RFaYNrunsXUogKrR/HJSGxWyRyTCkbUtmf4YxI3SYNMZ44bvpZjaibte4NDI54DQMgbm
oM9nFQJ/zWF+0SNnlZtyDR8W/x+NH9FssLF4fRCSuTZWUrjjuZFHOmJ1dQLMevUmTJbOhw7JEssz
Pr9t6gEmtixQJN2C0Kx1+Lrm8dvoxyd9vhWA4mkLLM4Q5/2gUPITABgmc9Dn0NDP4zX67TNieRrV
XY3BlC9W0NUAFSAQ8t5RvQRPpJBOxW7phOz4FzqNOArmrE4f/Ni4dm95bwHB1KXdN0hZepOoOWmX
di+WYyK0Q00fdF3kiH3g/HRhDIg66MJbqrnl0CYR7+16ecXmKy1S4ufXJkLveVMIkRW59IToamXk
OcP7hYklgoy+2Ee6C1mKnjG5V40Vgfsg730nsIPj9/Ya4/3ViBHhOIp61CPu/rVUAdwGOuEq7lZX
ZBLNDESlhiIeE6d7SZy86xgMVn6hxmw8tNDO9X4qxJTT9hN7S75DubFkZ+w5nXQTjOmQ3dsdodtl
LvgCWmlpbuieszee7C+ISk6OMMsGIAdkTu/sxQJitEKLyGONQX23kDlQWEiQ2KNEJhNHD3824tQp
7Mk5RHl95rWReoPfiQuoTW+R1vEsrfiTtEJo/b10BLQD9VNNZtqH5iQGuICgJbIMvMs6cbWYamln
Oqf2NnO3TgxjCOAJTCDj+HcflqeMYYoyR79NyG67o8NsOzTO39UPzPoB8vBvrApGW6dvK2kQCdvo
KmqHWhAHGMaR5vZbk5EplPwQyedOYAvlcOjIQ7sbqbQGyZZ+MvSdP7kCzjJn/LH6uoMTF4f4LIwP
JuPDEGBzGBrHdstWv/U5rDoaXpheRUDskbmFGXY245zICg9BnV28Mlsy1Jl4dHiHpbJkrYAv/ntr
c9ew8inAqmKsqvlfTzV1ChEQawHR95VqZVThpEPtjh4iJP3coae/a8cDrPJn6Dg2uxKc2dgBZRMn
bxbrAHkSBBKiswPsg5NclQKw7i14hnzGztTwfcvybrid0TMYjPXUZQrqbdQDe+Mw4QFQRouIXipn
1z3cy21dAdSj0P7EgIxP7YwFNTPlyQXcotOzjBe7z1DkZPLNK9+3fW/pkaYV6+GQtUOiU5y1GLuw
fF2B12LuIQo3f8nbBHNb8LbUud+/gz+WEqOwqGJXkE6kdQnd2+bcXVrBlf13z5m58NQaNwz4eqO4
xVCwcQTF6npbfqTNAyjuysM4wCHtcMBT4crsukvU1xDQKUaqfZtfjxhMhF90Pz6kSVU7+5xbA+Ie
wkX1g2sbUK9/id4151Uc/sMmEkk8M8Zieg6VQ/C4NCHxZ6YiqxJLlhwlkJe8VvxiLLLAPEmF7Hmw
3ibcpi9ya0V151XrlL6FShxLl8zIkVTfMM8w1dQOLEGAQxCSqITXqWVpcNFaQHvPcRJBeDLtrqaw
Wo4miL28Ga0F6y8kjuaDhQT6K1hRVJOBy/DcKsiWjVhL+wdVnfOQLbMQSJC+meiN026K5k9/BZNy
9yo5S26ictiRuYfYTHJbR2Bpn/El6iwGJsGd2+DyQo0cjDi8v1q5r7A7CMIlonqas1xA5J0uTWoa
ijlBFQs2VC8eD5qz0cMRB4Ce2rqAzcFnvbeorp/uX41HUHnPRsrqb8/F7wbfVlFNJhDOV9AkAGMQ
3a5F6CoJly0lafSMOndZlf/QiQUjipL9aOhQiKuqGrUcK0hrt9CsTTJYKahgY+7QLsOfhLiIurOw
FaIJz4FhPAOZxEhR/UpXcIld9vyTojNMVw04Tafi4kK8BZ58gspYphGvpQn3RZoJ1IqzkZEfOhxj
8qzXhk0nrWiEXlgosUU5c1l3CDN2nMi02ZCFCfLDXxfDVuABtsXVR2+7/0BZn4u9t/kn06SX3eni
31YLdGs5hYMNLZhRbN/scPXntUrVT4E1gLV57JAJob8hbr8SteAldIXG1FaIjb4LkPK0UlSo9S+G
yo3sx2axqdtAh1IscSycQSNXDEjAflBRQgxcsVOJ0yzkwoH4GlGJ9oCkpwmeWCB1Jmd3V34GdRtm
/ESH3360/ecEJ3CwUnatjf9dczUSMrXprFBfhz9ggRmvFyn/THgXJTilUZm8quix0141+PezzDXg
+VKipxgS/nT8i5dR+Uz5kagt0rlpyv5Y55p5kU5VHtGAq9hXKaSorav8FWi5h6z/mqsKcLRcNLdx
hOqt9ViNQ7n8rkrvEL4lZLhXDUnq8v9jiEMu3dXhNkOWyWTRkdUe2UOf4TWZuBJ3xxfsDDHtJPPl
dedl7IhMskl+ELXE1OWDBt7iaCf6R/oPQe8dX5YxK8fYO43Z9WNLQCa2GhgqpTXdkQlL4BnoMFni
FXxlzDc9Xa8/6VBmAt6aCzk2VBTfA3BlsKDPffiPZp3MmaDtppg8w0t4XbLGZKGP8VaDwNgCnGbW
FcDiuUdSfIbxCCDM2an/KXLxSWifH61s4RC1hYyvP6o2VnbDC2RSLDNe1dpPwmslN5AgknFp8Ctf
4cZU+0cLZ7RZMWuHpGoPXWZHbIIB9HrmyB6vD5wsGeKCfxMp0rjJXXNpsdxS8OpjRKvn2Otq5KwL
4MLGHcc0NWBINtl1VDBe9pZuURyVMXPu/m25L4zYtD/fK5YKTQ+yue9TcTUZjSxKxcRcOfAGlB53
2pZU9mqfYi9YUD/zxEw7KctiOClL0MXJ5Ohk8CDQxBgU88m1Id5fRWQDrb3hQRD5//q4b5nLmKSu
vXLNqE4KSIE5QEg1s6r5DQcILhltZp9s97/3rrAHgph4VFSBKcxbEp0t3yRvyLVPZ/uibYe08WU2
yq+GeaPyZgIEnZnNwU+xBIKWOILakMu+d3/YF5cEaUgPD8c8RKZdZ1KNNxhKXsbsY+N43u/tz+Mc
FXSEg3mxJi63rQyKyuis8uKlqaQjVeJpSQrg9sykD0noaBi748HV9QGq//48IIKW0tmT1+q4Wr75
ZlPJOTWP0dCMD8IjXaBWJ+53PgZMCoTSSk98NrejAc3XAfnnTS9nMpZ8wJelQvoHbnmuXglaB25x
HdTmuH9v+hDf9jzvs5Obetx9MyES6SSmBEUhcSJkBtUY5QnXjpafh1bpRC472KSPezK3w8JEIwT8
x/sAekxrSjJhLDxgswC0ChuuBAcKgbRZYagATP9Lg+Z1tj9cIKk1JO8JvyuoO2iUc+VWm6ZF++en
5y4au5IPKQQ3Rbn2pplVeMvWXu4SzQLdWIAgxj2MYr2zYQ0KY6/tFewDxpCGKGoRhEfEXFzxWrzp
6VjEUfKWl8CGTBrXx/Ez4dDUDN5Rqo2DStk0SPMNuWAnUxLKfe3X+sR3bNwHo4cMQlZ87oIYW/8t
g6ifqW5+QpTgRL9osRbr5tXQ6igwmh5a9u8vHZ6qZ+qcdcYLZxzDMRsegJP711SQnRlc4KfCR+xW
jE82l7Bw5XPA+l23/Pwht2G9Mepyz6fM8Qs4MAf3RMR+WA4M4QGNXZZ2+a/CUNueJPe/n4NuK6q3
ImzKz5Bybq460XJuqUl6ILcbm9BCgY9tOZW2KKxwWFbXTv8AIAVzGbs/hZxPNr1per+Fgw9LqMGD
2Jymil2Og8mzC9wItDwwLZDLlfOpykaSHAoh2FcC6DptTuU2LMQdV4rW7r0OwJFOlMiM/ep3vo3s
mtBymezlsBI8RW3vl61QGjXOXW6/CIJEtt0ziPWL8+HQ3BWweMTnmR4ATK8RKRXCpQdQ1ggH32ty
nTlOyAsB+4zzYAWZndsdsQSB/sdRVwG8T5o9uIEyWbMuzODww9NcUWibYqtcRQH6KzmCioNbUJAK
wWTqbav0XeC4B9K8LdRS1uvWHCo3yQSellbdrK/mMjxiCG/reORDDLxB+NWWEf7HXU0C27hR01zM
Zkoj0zP/rp/ZmbiQNReTEGaYWKSOmWY1co9JQ5lMDaIY/CXZ6fLPPNh0odRjxtdnLZViEfrpMy3T
eDQ6mFAYtxB5OJfqq57jjIWAqxbMyON3HNRQrgBx40rrcD/+v1YZmZuaCQkhWHiu406q0dwbOKDs
GnnponOHhCmSCkEI7GYoN/9pZv5KA4DNq5hYOOxmbTu8RanJcbozNlfu/zPZetL/bb6YUn4BQFTN
Y0tK+zCp5FGXuO0QztQBOx5UAwftpqusnbuYP5r+a068jF+mZ9MHXQ9JKfTQYZ/grXw/qwHACazJ
gFfXdeyxKQ+SkNbf1nPNxQ0Yv+46U/JPnQVYWPWaC7lgye2dhuW/pWDD77ZOL9HWBicc7fhuXf4C
9qYInzb5/aiuBJOgMLELoBk1NzxQro+F0E3zOqCxrVsF5lVi7wY+jnDICtQ9hxhGo1x2Ixyjxgx6
PR0kzlGNxf7fhEPuhETyMAHVMcc8nJCzF3mLmT0geWIdW7SQjfKiXYSMxpzN+aTb17avyVT4h3lr
oYjQ+uhe2MLjLeEIB/YG16ztTH2sxFBt9SA6Y2RQNxnOEgkcxIWvnotbOTpbPQKW/50FoHfeAb67
afIlnQowK/1vvORoY7SlCP/rWYVPYPrpOxn+NWT56RWeO/VBDe32lPrPMikwvK6Mxo7sCt2Anwu/
XGzxvI0d9I63F2CFpgF7h4C69jMY81AJoJZKJiJqhUttFgviVOsGQs0lXbN5qYU8+X/qxNUXW++8
ew/CilxGWyG+vxh4pqHT9mW90VkcowRvBSicqRajkkGSTdou/Zhs5tpTT9Uxn9FmUOylJbL7ueB7
gdUKwsbWoYdRTCh7P3UvECU9/3m4PXLPxLO+uT2XiEMYX4dd3UBXYUres4LiDXZsktaXQngyAtVk
Jx7Oo2+Md10NfVJBvQ3g1T8Kfpn1oeF+gGVsRDRER2NI5HXlDkx2dQuIt++ssHzZnZL+dI8fLwiy
5wZPDGS+gCQ5c9MT/YxorW+E8Tb1pb3Bi9Wedz3eS/FO0Nc8KxTiOFqJYvk555fPjrUhO70cuqNg
ACVV+3ZgmiSgDu8XV+Sv18+NgZLMRhnPrtK4IliGM5W5AoCUU+9s00MG7heGIAMzSJWDAdPtpT43
qL2LKElwD7mkdOqm7AoVsW4EP5QkmaUargAuW7paPNUAH2ph7kdfqUCUUIdlvTt6ardb1HOT0Q15
kmeqUMJF8nBDhYKPqS62GZKv0BLeaejbfrKY5yiKNSX6Joxk3r1tGlgDOAEB2i6PEiMTPj4vVOwW
jVkcqxmN+wjj20EnZLZvDsBwZK9keZ7EWbfjGw4859rEXnoVdTZJLuECjHjY9FV+an37pCu4My0S
OSGNw8s7Ty2sbvthPGxoO1epRdYys1w9BDiOVQha7Ow1YsgeVKPSBohyWYWPuqJPyFn0HMzv9YiF
0lfPTOJDINxsjCwkc+ny3A1q41zyFxvI9a+M5LRM7wHpDraeTb/olH0Rq57tHTrPxpCtngQLkhs3
Tu1mpf4gq+AvjH8opIarLGVZX8jK2BvUgxAgoDBKhNHAnASGl3Yg2jVkTlelBm5DB7H12d2C4gAZ
TOX8K8kgX7EbHQ0HjHSPbZWRqjiBRTcbTAdZJHpULygAPovRdRWE+gF6Yh26dQPexA+G6LbcgylL
mNYZQpqi2JPH9/qkqC5bsz6AUB6g78PtVJFrnJcQ0E8MqpfZbJWvyh5l+pjSrR+ffPrq2G3WGBBw
Y4/BEPJZwt/3TcJ/XwcMOZCX6+YFxqtfK/MdAICeHt7pC5GwU3IgflZn3U7Zt6aPOmnQWMkwhJ+p
Cz7A1eD/UgwtyZmoHRKguSs1F0uHeaTiFPhIKPSewsSlQlW4E8gH5SlpB0Q8PuvOHDz5XSeX4Cb1
kr0OhbPW0uTq+Y2YjC8kDtR82xYWBoxvPov3JSKnRePs52Zb7Hd/LQxh1nNY4XklwjSJvpRyRe5P
I9yu9OpiEALCOcSZLwxtysWbPYXQqqkqxRMk51hEZ8MMtCffWJA/ZGLkyCiO9BFRm9cwBd68CAPY
ZMA4C8RzxNNY0CMghNoHOxhBNTTKatfZKIS7X1QJrWNrqHRxeTcgrtcJGvtL3v00fDNGTsICaGH8
KVpJCUmqek9ec+OzQoZOkGDC3pWO0yqjgiG5ymhluwi8+ApZ7X23L1QQS6mnkEbSD56D5LwXUb/T
gi3A6l+WH+X7f7rpqIwhU38LvYiPJxy7QXeJCH5b42Inl5oLw+oFNtLPDboJ8LHpfCaBOevY2gHx
ufiGOB8Sgkr0QYyye95aMjjMvdxPpIYlzTkRUtnwOHDUssvUbtFpUw9EIb+MWJfLIqhXJx3nG6Cf
TYHHNVdFCM3tURtSPEsO4mi5TpImSmxb206sWXpm5XLeWvgXE72w3wxcr7hanad96/woFE9gzc1g
oIPoode7cKm5gNSflLTEmc0MS+ruLCy7Aqds2idep4YD/7u+6iz77KCzIPVA9lXZKP12aEXQj+NB
SKKryI0g0caV+vDflqrBNh3bAvRQg08JIdIYbpnJbb7RKcO0P4pHLiEGA65hqyHmCJbVf9rRUEvH
Wz0L3Ja6zSwzzmF6S4hn8A9MKVu8B1FSEsokkvTZrlNBONx0+y0gFewqHObfUvwDCgdjTods6nS2
m6k2+q0r7Yv97WiFzyzp5FNk7KrP8v48eLCvSmSnpNIdLKAVuuxHV1RxUpUVrwLkC4MMgSiJcSPm
oIojAyNHHYFU4c9pbUm68Re+worPMceYNH3LsHLKAD+m3TrXQzPHUybcttdsdgcINpcWmRUVYnXp
SlU7yhMllQhOFOHKpywjAJedqYUB8vtRwBU4HNVaqQIWiyZNgjM4ND0zhfoHVu3kQVf1DNPkCv9l
etA9wgzgtaaOxHOYEN7VqHprlAm105zY07XPvC9BRG6eGYsjvRYwNmQlTkdo1ZRuxroi31SlE/p6
PAuio4WuEAT9ZKApeOoLkxax1Id8WRr5H7ilD3KBEW6LVnVdufDWGfdUrgIiE3aHc/QqK/z10oO5
NUARSZfwZ65L8S1mJbKo9P2wi/lk4SPU4ZUhd4UQxvUppllq6gq52vK572gq6ijRv2mFeVfyN3CF
FbDZH3Q146jQKXSFdjAdgkTnR55CXYdKPLBFC83hhGYHdkuXtLvla8B3TAXIFfrVyDMABI/8PveE
SIUUAPQnbuWDk9Yu5Tl6rze3EPIrskqqm0cgin1CiPV41eflr7Ep/X/kdOav8jGOEI7/+8U/WFtw
YxnGqSf4N2tY4dl6H3WwZ2l0V+SccoGNpY5840VZD8NLOp0NgiqjvCfxuOvDXpB2hh4D0c9gRS4L
paSx93UE+nUzPozFuZqKjM2Mz9DDAle9NoujmF10t6KC6dbzUn9H8eO2F5gMiVS6DFZDzEHJ/KGO
pDrQaA0+HMAhyGfkjwxpr1M8kWk2iIxtMKh8B7u2GgGfP0SodM65todeEONRrUQzzA2a0cfrOnLu
oJKUvyI24G4YfY6LXl42Bm5i12tKqTnPkeYZJrGKcwj3F9n/yJ/UOPsfWcYmILIpLFK8h3z4BZ+K
fTtAkLZ9rEKdkjSEfyUVfeTUDNbooLevNOXK5le8si26GwOdNdNeOGbEpFa03fnZIKcqZ/+2ERCx
/vl9uzDx/INzEIeqQA1yfuqUxiIDMRLeuiytNGWzzJxurP/dSEheZyUBm3JvVH19TX6WaXWNnEey
BbwwdVY2ghsFl7PGWUiyb0JxHMTRudc9EW1UIyADvFh2JgwRAIE+zeGsKPIUctF1dW6StDZLPxjK
kGAg91xVKocAmVeSmvjSEVxs7AwE6hmXoczoIch0Z0sEPS1UoE/+TbAXSzJJBvaqlCQcWLxCUEb3
G//psmWYzJoIirJBVIKz7+DOuQXv0YCRclTI9fjeMYFaGm5xLbbD2VechfuCe3B68BouSbmMyNt5
POhdaunB3jSpFVbq6qzwDn99VaNy7bxmxTzoofdXsfzDPF2TxvUtHjlC04llQn4X/YlbFVNuo9Sh
/TigN+TNPYp4+IRx5bKv05ql5bSrUEqw5iiMvP7z8qx5NON5bEjM+zzxhcTbDHNUVKQRuWwv2uGo
PfFa0JUSKso2DnzvOCMOFd8buK1VBaSB8pIxZRbQ61zeAhsoDGzQpnPokqT8q9pmSRK+2zlZvSR+
ntGjcVtffsku35FruNdSbeHo9izTkJaIyyYgDTX7OD39V5LOu/DJ24wSxm63bElRuyi0V1JzIBYu
9JpP8zE/AZQ4Urt7HXdASPNyVuTZFRWDzPIp02eBRYgJ9iIUAxS4fyM43uitL3JrlhEFGFOlGkGK
wc+Do2Vgcb09ASYZBmbTmRrlp0kGRY+ivNELBFubUWmGwhAAocq7o7N7qen/nbhcCuimYB1kfwnq
IPkY9b/rYURVPVgGI2M0B5zrpT24Gox95ZNc+lBdHwJBbEsvwGLwDJeKvQTNaf0var8fgnWrUweT
uktASKvAiI0yOSQj3PAadXL6aa1uCGaXEY3k/u79dpnVKiiJYjbFG+r2mGYVjItfHc2eCnBiwVFh
xpIUT3Lr+LcRkNGtnRUZ4EBlVViT39ivYKgmdvH3tP3GzbVllfeSww+k7a4+e01c6DbZwkEgPDQL
qiAWCC5jDvQ0mM815tuWgjRjqJwHjNrf2Y6v1xvD/ESrefbw3+HpKzdu7SRcIRATJx2WYEFJDHyV
HRIlEe5TlplsVj+PwtfkXxv5TthZEmyPswC5Z8F5ROW6i2aC7/1ClRdw1OYVpVzSnTIvf0e3jagV
TTZUkkuKn8DdzIsoC243TZVoXfH9Gsa/kiKZh8zQas8Jljc8ZqBeIxHB6FHvEv8f2rtAr2x9ia5X
3fRWwUcEcP9JDQf/rg9uBgX8bib608U3AhQY0LMpveGZJ1Lj2/KRp3Z3zvSErZ/1KOTkgIzK337g
YmMHRfbx1cTjquHsWG7kU8Y4UcB8yDMqfuvo8+I3oihu9nc4OmjEg8Mwj+DwhvY7EFBYjFk5BOXe
3tpeyconNwmsRlDxG2D6eiyUDNz+OcW68jbd8UDDH4/BmGlxO01GJOs1PeQrIlWBSYT9m0ki2gED
mrCj1zi2RHommi0HRx5aH2/n7dR5fqKF8aKsJQ8peEsEMMikLGhcXQVzIOMPENExGj8nGrPniTR5
lqao9nJhebraRGe2QAWVFMURlhmIE+7px57eAOumKvMlI/C6iIOTd774dwn0qod6WR+wmkVaBCmP
OTWkgsXKfGw8/kfIks4WsX+DjXxj3EgME1GG2vJuqUHnmo77OZ9n49czsvCQCL54kNNWGKEJhd4S
INFqNHRN6O4ap+Cmc4ShJvKJCRxW984JEEp2A/kZ5Yq63dEP+3ILTH3lMAV9nfaDWIdXWmBa99Oa
i42c4Isio6n3cMDAr1rIQM3vlh22G2tkCadE/RsOIkWc9ctVm8TTuDoG530cZzGxQprKbd/Fch/f
dnt6i/vvMIOqmkdbR+Jb0fPArsdPKl6//qsptgAdpNmFj0Zubhc83GkzE91ifhfeyEMW3lzesc81
+FRzHQ07COrcnOGvsV1PECv9z2Qrvrv0HTTSA7YjpKJsu1ZDmOZutGoCfVpz5Tk4l1aexuk6Tl7k
VKwT3GK9n0rZ8cXg46cUZetbyGVH040JnUZYkeKKuuQPNh6ZHKuMHKfiT9QWDgWFA4mf4DOOkqRr
fmk0/w/wg8lyycSWsoULJgzWugADF/DsV7QBJgd1C8OhS9AuXJS9gdPg7jcheeG0RiiX+wpgafNW
e5F4m1wVBD2r48dC0YC4jzz25rdby7QS4qbqNiVs/g/nGqnSFaAptAwVhQztB4oUh2GISMbrPmye
qdft/l4vlVq6Od59c+knSTqKfbhhyj1XdXuI2cyeHr3SzAIHHC3b6vStkap8xen9f/y2shnAye2s
ctorSZ4x4sHVbIm9guAHlNt//ly6CidwYHoPmJ7wzKhfsqgIvoDZIoudgc8blI3QdzkpWe/DH1b3
U/ioWatULYFoNbbe/vlaVIImBd/z+zHqiAevuJOOxEcRKqNx3btQ/Vx7wcjnSqUAwq6nAiirzkDb
nW97wNC/NJxp3dR3fdu59psk6sgbjCosoR/OTxvRrvKfBOvxcHpWA3/MTOs6z4bLokDEkje2ecTn
QGeQgFpoxOJHioM2cTFwTzQ5Y76jMVvo6FTvlEGBdu/qvjjTBKlJGTMgEpHzxaWzffvufW31EmvX
nTb1R5+9xefCkVWFCUEqY0hFQrr9SggspuE4mwTZUVRsN2v8zryfhzTsr2M+25TqZaJpkWORIErQ
GpBIeQbKiE/XxI90XqXZe2/+BE2uEOdbqANNYEBpRXxFeeT1rAUOrzDzja+yk0ACN6F6pN/Jlb6Y
mQ6/85DaqScYM9HYzHogPU9XW399SQ6ORXr69NmWHTj90X51aD7CJqJYXcYs2C0qiw6TmqxRIMDn
kVzzQO4/gW0uuq3zLp9Ma9V5qvn4m85sqzvsdbySb1qu+JoVlWXBikF9pR13T4pinYXlRza5CAmg
7SY1/4fLpO1tU7OIKCLQklEp6K419Pz/nwcU5m766DlVl6/Nca/X5Qn5l0PkD41cNHvME3Ka1Nop
8u71PExk7vqQxXTn4WrnwSKt49YB3oen8OMLlCR70d5UAsWn625v2A6Z75jcXdmEJ7xSPHJECbBo
suYKYfau4KoqN7YBFyba+t9BrqKietfspYhR5YoxhOVEqEnU6fdsBlQbCKduzWaNd6AE2+borUbJ
XrJPaVNw4eC27Gd7OCDZl6KNRe1TpfTncaZlhF/lp6zlzBuyPwa3Xj1HBSFPHO399/p1sKBUaqQF
+rFiuYYw4LQXepag9fXTJEEq3HatjV7WjcVpwNRWPo5WcnHdaVd0Enmg8LHqzGX+pSZIl3I1RuNK
9W2CScX2pnk8OoAQ3COno0WTC1SaRX1qcRsHK5PmepphlQ20TUkIhu//OtBz1m23zzwymDgHBa34
AbupHYktMLkz2483g+s9bdNSE4BWVZzJsHmNnWIJ21vJDmJUsEVRRmJNKHaFHVR66KnfVo7mPKNX
lxALeN4kBna0tgOmHxt2UI2zzYumHQRSq+XFZiYse60TNLvvh330SkbUqeqSkUuVYf5BOmBtL1Lf
wX7dUobS6Ym/BE/tiLjdo+k/UN0UEE1ji7p4ziFLtgizAOW0hNI+wPxgqxTBwCO0inPPXwJLtH3L
s5NhAwSRaOtQWrLCutYuy53VnhJf8t4MS8E8HP5m0OFCUo/unQwsL0ANYOX/JZ4jbsNDih5LMJri
ElmvDIFJcsbzbvUcGgc9eJE7/FzgeRN0hG1eE1gHtdScIsA62LpuC/fncrlntVsr5j5v3MSIeWHw
UFfxmJqSsvGOkjyK4IxspbI176C/FJE2zXaJ1//yhNT1oSr7EuG8XZsEP6mOiFbZuQkr4JybHhm5
QGaTG/R0+C5n9+xVIgMkWTQlSJB09FS+YDguN26zx5z0n4GXedAZy1BBsRPqYID6Xl3rpvGdNq28
OggLYY5h32aGVIgue8sfFbebP6psVyPOwvvhiTJtDJt0Qo1shx8bWvvUgmEGjwqFjfZu00BfCfe8
kQ6nTBDAHeOYeS1cuQh2wRLlKTsBWxxY+c5zHi449esxIuWq8jSCnLSqpxQqBx6YaakWyxCS8iD/
SeowyRWah/XzWCVGAuIpK7GASWUWruUm6zD4R5j3l2S95s+mKmFUG0tjMFRfIJceeSSlNROwSV53
erzsxga1umT45R+Hgx8U1pliWpTlAQhE8FRZWjhxG+aF+VbAuKkMF8iInsu+9GHE2RSl6MiMtC4M
wzCSA6Pjrghl363wk6eEAXmXhS4bIZpT1jcJJd/+ZKqYUWZuE46BiqWaTyapG+d4jztiCjDR/t+U
cYQOD/0i6v86aUrglKso40PEIVv8W/Mxln8Iqnd3N0dcZ0T6X+vZRAvQM5mXWu65IsMNkaZs1/+8
UdcvHS1MIVrL9gEuYNCUkGPEIke4NlL4adC4ZEQA/GamBFabAfqJzTgUjgakJ+JqVT019BtBRlMS
NYydR6aoRMJjaApYQdVS16B1oHAh+Wy4Z4+qhK63JBwDTtstU9gvHyZlOq/2Du604q5z6MCwHv5m
JYZz5NbQ36fqFox9adSiIkA3/awvq6+zWc7xgm2CW9t3uAVdAwZdbAXdRlFG8eCa2i3aYDtPhahc
4Ku8VPvZdsD6nKC7nXHEpFeZfUbqrkZudWBMEzyIVzULlxnLR0AdQbD9YtD9CVn/eWN59eaiTLkR
O5NSVugiNiRO+RU16F7gRhT0IrgPWZr1T9Yt9Z4q32Sb4vZFoq7NYTo2IRJVES+bTtMqvlDHw5Av
EUyScVp+lI4vacTP4GL713T9q7FcBqPTz6yDpmKKmMHF/M2xSgY6TGrAIRq4A5q/FpWa8LyaY9bo
ZR9CmyprHUvPtjL0lPcSR2KYCOCw1OkJQUFfd5tlFAL0Y8Uhjx+GBkIzXjElVXODqCEcgjC4RuDq
Rq52czuJhETUMLJBUrD9/v+5zWd4OWMsr/h8n4gAOSAfoav8TVz2ce4yjHq2W3kvCQJn+mxddcEI
VddEoRkxA2tKEI8Y5fqlaxslqOzksujrNw1eBVgzFq9uO4iSAjOzEnq/ioO2NkVnNG44w7aP4mDh
FfGxqEoX2jyFqLSuJ8BxtqVeASRLrJmueK3mBO7K68wasKye1O+nupVxhI9hMcGHX5k+SYRMSLTU
ud1vhbPdDyz6kdAQHDmuVImY1mL8GAhY/Ds5COSppTyI89soSmwiNNFOAaDqs6WFPidl071fI6eK
bHt7LBuK6d8/OeDAtO3hBDj+9fPiTiCw3k+QsOJNXUiVAobMc+zZEhp2lUuNom7UVHjTKVBn28Qi
hUWSonQXTWZug42VD8aAJp+O8u+GOKll7M2k/MXfnB4BhHl03xyIlFla5rXsXO/deTNx3E8T03JC
2U8ZCEIIGzhTVn2tgYkbzMQjfO/maxchpIV4zUcMjLdHOZGQl0+qldZwr+WZ+MYBeC5Pq7MtySl3
s5m+UQbpwU3JNeGi9u2KVamb2CTzwzYw7W9ExdiqOO1qp0HnfL+FqASIwOcP6q9FfFMDKjEgEXZN
l1nz42sLOWZFnRN9KspkX0YJo2qUEpBt3I8S8dUfzajSf6N1c0QVJtXdAvC13ffu0mY6wrFlIrNS
HuEgr7F1WawbPKCOei/7yC94/tc0H4JN1BZwHWjjEZP8U45N+J9/4Bvs/OOxkaxAOSOIusp0SICz
P0OXvMcOHsFwI2RYxp7K5kRlz3nqeJ46rBJPB08LKsY0xKbgv7JRXamuaywSv89Z17FP0ZXUNZif
2+mGZfWlA+7YKKL2fAnK+s5kujOSJe/nOE96AZjMNDn12DWXWzxvOYrP+pIlacgsQoR+a+Djs+CW
M7UqpL2LqMQm9ONV6fKq4BPUdJWsxs8ujEMkc/j5wwt9OgvDjJNB+YXnoFQJEuxBFXa7Y4T+ZgrP
Hd1vcKLR5Z68TZ2E+YGhxzO+mXkxYnFyOonYkQT7jabZsJ/lzKUf++YRVyHhohn5D2GoAOmwe24P
8mNWBaVKGWCTgLpIDWxzGnpKxc8MNFdV5YF/V1Hzo9b/N73zysJJabBFpZkSQ2tY29l1fLFiV+vf
L1kaXaRoVDqBhiiTjb6kXgce1MAko8mCq6Y7eYtTjhQaGJVR1N9clB3el6xgfSaDYro6yTUuMlXL
lrkM0WU1Xi90SuY6AJ9WdKrvcBdYSh3yLmU7xjQp6UptbMoy6bsDUiLu3V6OW26JN+/SnBN7G5Yz
EtU6t1soMlvpkwnY8f5/Zdqm1p97GsRtcrXAVz4qiiC/2oS78350zhS0p7NWFFSPWhraXd36A8QD
BM58QkhMTh6xoC/iL86Xxi5K1Yi8UxM6VxGeKURldgLsTeUYLyWgZtJEmpeYKVlxXvsh1rMF+c1V
Rj00kDEx0ymMPD0MSkzZTUFIZQ2Co3TyQQ6hduI8wh6e92FTp+tn54n6ATgH6Nq4Oy9P2Em89Whh
3iA1pyfFW44lVrQjEdPLhh7BQ355OzN/u8pdA3NuvIY7APkFAvxpEsDZupIZborUedIb3Q/QtOwT
8+s5ljrFrh0xa7tNPG2hLcYAbcXPXw7GvYWF9kKQUyDbn/7AxYDMe8R4Jj2Hw/7ebzKs/7t6NAYk
RyyK4nJDv1k5MTOo1QZuLfPLjow32e0sYCrrdGkVC/lFcO0Ec2UBelDv8JpzYdD3tIRCmzBZuweO
QB8uVo9z3cOMvtdhVamUh+4dIjXCvU+w4y8bQCvMQOT06AOjKoFwdAC1v9M/j1XKlKv+LXVQrFC6
XnUCA1VbBPpN2kcdpDY/HXJATZTSghCmaVplE4y0OhwiWe5iZAg4kOXO+sN3TMxvy3l52o1r/G1K
JICEmMrENT1CmwXRfKaVWZmZ3P+2raaMOuQ7H6bzC4FPnM1bkujNKtTL/Su0Mag56PT2Rh2UX8Us
w8/dv1DrlPxSvkZkP0MbT5chfUfBman6HaoKovZytzUm/2GMxFj01pdo1l+IniAY+/cpODZqRCyC
N6EaZV7uAIOilAVu2HNO+UcIzLhuWRA7RyejzGt0PHO9JHXXeMjboJ5freVRcfvSdpSsrKPwc/wo
eWRMFE2yCTWi6+0kpLTrSHuu8syGP96bkQum/raQBJL97cqCyF7yvdTKtnT0rtxN7B1j5cgrmELH
EOiftGRUjCG+qrASTPsdxnl6yAyFyGfQkHpGGvDpH/9Gufi99fZhAauGSGdlwjMHQy9cczEEZljn
DxodnO69Z41TZBwjS87kxmvl5pV5ZtD/18/Vub50fYxoLtlbQcat0fWsOP7zxi005cBckDQ3SArz
QCQIbDgpqzOn2hbQ0P4AFfffDJuLFElQaa/J6Esibeip6XaAI307QVvjD0WP+JX68lltH3y3/OmT
tVCiExnXREwqPEHuzj9uidmdfGg3540BeZUSUREBwpKMk6xfe8oSbMtG1/ArjA21z6sOgxrC1Pky
Z52hp55Bdqan3RHgFFVzJwMDVOfCTXigCR493HMR23LjQnWp0l7OOG6eTgFpwqkF1psULY3wEcBn
T7+qDLCxYRLEteML+IBGfyQivgpvfpF+zSbpxblIge+imb9zKwhRrLX6XXmc8af0r5f0UwJRHJis
6YXWeq/7C7X29CsYreAhiSOnm+3IXrzbOKhHHubrTyuC1PN9kNgkw31k8Wx4R+kFaoAch0QHcqGf
Fm6CnbHFe+0rK/7+Q86UTbkIYRjPQAjFMLyE0Mk/HFGEKCYsJKZ2cORSxJexD+5IQzWlAQPEEWlG
1xemjJFSQR96M2NY8D6T4WygT/SayXDI1Y/yVgjCxYFZOawptvhnuMROk1RhBu5T1ZJOyMWCiYO4
0nnsAPelvYvRI+3FklCTorf3enL1UwVewo/ZO2j+Z0pzpv/OB5FeQ70DgFMJqoPg3fU+UlGJpwfL
A5dVjW2ZIjA1MvLOnyckiEnG0jp0Iqc8p7ZbKklmSD50TuUpLmlFc/P30Ef+nOc035+KU1gcMGw9
VerKqworGGdOtr81TFmArbPdy7xzjnvc8eyBoPrIHeAqbSpeK6IBloxfT/mNr9lQk/oBbSpraBlM
uI6s4+N2AmSrWXz+kBUIzw5+/1BYa2vu9AGRMHoJ0fGcE4mhcs7dB061js5Aq0aEIjKkeeFhTZQ5
BBgo8xZ7fYb2hJeT4IlvsWz1tbEyqQ0pEvW0KwJDe2vLnn8KEWWHA0ep/L8mrs30ynpUwhC5b3B0
yeJe2FLKoP1ArIPHhlAw5rqgDmgAXyi1oIQicDVa07nCcnbzeW1BhlI0tdPsWSKF7lTWUKXO2Y4f
h9ZJEr1fIPvNjIkdbOOCswHv4h83MiaoW/DzbfCpU3SuiOYmSARckquHuG5AgeKv/SAFDyGetoX4
OvBMS5Md4J/MxQXe7PTAWPVPnAgq4jbE0QzwCesi3yN4zaycEpFohrtEn5NTpDyOOi2dVk70sGLG
5wyZElA8sgA0xOmawkAQo28Z42gnSJKm6CcspF5DUxB2c3menCqZ1ffqezqaG6qgPu7rExiPk9Hv
UoaZgoy23bX0djao2vn5pQbc15sbHHB6rOc88Amsy37kyYEP+XxtlPAZOQKTEY6II4l98RcCQ3ZR
VwdQbDzDoZFf41GURWTXixfYP5FkCuOTxaNvOY3eMIOdr9vw7Jt4IDGvhoGpyMiIhI9aUeDsiZ+r
61sm8SJz74vWHuTiFrZK4ArycxpELVtMRy8Xd+hCe1pHPBlo9i5KUpUIxgITWdFr5K+5OU7YUbYb
XOBY8VuKRL9QZIU1g11Nt2qiSvtgCc5bZ+acQh3NFBrZMyp1fuDQ+1iAQ+zP/bDjcc2iHz04Nieg
HX5TSC1DAp5+6JBAGi9pb0GG69qf43Md0ZHOg7ujyocwN4w6r90374ycE8K4Nl6JFYUGeA0TO+Ic
saCWOCq9DHuyQCTv5/gbe2s3hm6N+16ShNMunIkLpkiF5/Tchmhl9/ygLrcWdcnZj65oRv2M2bYb
diVdCdPTTyriRoLiuzFQzvp+eFLDxYIAsO6x274/vkiEyq925xDGCbQ4dVQ6id766iaSWwzgUl0O
J/4kJeiupuGL3uhivMZ+m49DWh9YlwW6is6wqhgiMBcqUXgdUIaxRYsqBEwU+rAla+WriaKYsVIz
CSVersfdhLLJ95UzeNdLGqNN52nH56p7Y77UxCmkNLz6xMQzMrr3EX3BIzPOgPRmpW5hkKS/euFN
w7r+b1+a5w3L6fxoiPstflRUTC852qgWRFR70vE+AqiIqzPYnALfVmJETBBt2tnvdmHuIvzXcaq6
4BPe8xm6T3cha0XvgJTBeb379pspmETb9B6avhpzUt1wayQ0AhDINhMrptOuP3vGP9mD3uLIulcf
t3LpiwbWIu+egRzRye3+2N0jhQH0CXQJdWWmDNZxij2+X2VsXxjml90t1LQ4v9Ey46EUcGAauHH3
4Y7z26vZ8UidQzaumGXSEr/a1kFhHPak4XpjgeUAlkJd5Ubhcl+Jvm1qEnrw2kSeQXnS/hT6OBsg
r7jekj1tuxp2D4yUMykBa/QSmg3M4DLI4jDGJWqpR99q42cIeWnwxQLa4vIGjidLNxV3q/hF0gDa
KMQlC2qsJqYbe7tELSc8fJ0s+xEplKfyu6cH7kGPEdMHTSPGtbwXntmFvNoBvcpulANIpZV2DCzQ
zPYCdmZ//xWWKn6Dj9Iz/hJ7v8gFRADCLqU3KfY9G7Ia0x1RIo87PcFij3AFXm4KKjq6Isc2BTFZ
RInHQaQw5oRScq61KWCHS2OkbORQE9pm5JENmU2UxSfiFlxZ3X0rov21veZZaBbRjuNL+EcQ7e2K
KaqoWInND2Ul3wGnhdS2bb1yZYpSeSnM2vxnxTUMy1Dxx5JZY93z4gHa9Z2EBVEdr4P6NPNr4XNC
bcTQMvKrFtRPf105UTfNu+6XvKGLTwVeYum3x4yqS0LJd9kqeNx/zSQRrxef8IkKWu0IxxVQGaLi
J8O+xIT+pQQtmz1QrjJCjMxqepnW520cXOVUbbyZsx7Kwf1IRvBYuv2Zwr3WY6dWRCTRaJr4FtVi
uIMvpdbnAEW09oZIF1BAiFD+N+RmRuPobX+qlg0f0ZfEBBHJcDN3xk2qmPTWR2Kra+DlqqUWsa1Z
9YwNfylMs433J+w9LGEqwLXmhKD8cHAesw8bAYIY2f/9GtPdr27VzTfk6Hdy3dwcIhm1Axe4T3hy
odLXrOcojQ3IfO+qO8nvp+AADbt+xNWzjglsyOKq3mKti2eJ9fT6TsHwwX5mzKeCPiADS3NjYL/g
V6ztJKwz1ptPGJ3sJkfX2/tkOkvKrRG3QNVUZD+2O/nNmncJ3DgWxyfulX1UzM6RUQ/Vz21CDbtp
tMrxSYfA4vCSXYA4CeZtmLNqNTQ9P6MC7NeBEl6AoCyNs01tvJvjEIvI/G5iTUNPEuzmh0nai+0G
4IrmcA+/vQJc+7kUqm85nk1IMP/M1k1UXFxAY+FPj+oipKfIq/TptKkY1quv2EDQA+KCMJR1lBow
nitfO85vaStr1DXVA7h2bZUQJKaqIRdIQNoZPhbuJQrGyRqbUCPZKB/ezutvGhGJiu0Y9aOvTkfZ
YOeWIi6hkAhZgJCZe4nQlbK0f4sIzrDoBD5v8jOhC6abi66MTaMSEE4we4elHovp4M3kiHsDB5RG
PjqUzzk17N/cqL4bh108p9cIkjbP1Anbuu4aOU2D1ONa/L50hYq7nx6V+jvSeoBNOa61BTkxEIEO
eGbe9RLsdTAcsrnSz+8J1yS4eq2oPBaF2ttsXj3WOtbiFs5+IZYB8S6a6LaugvHuScKRYlwLi5Pm
kK/ugduoxhPrauszXIcsMnd+vGU4Nmw0BRzkyoSToyF/QTwjWSNE08UgZan49H0bPAlwaF9zbD61
XgqnV7TnvjLaYrrIP2jQkIn2pTUfZvCrDIDuyvDFtDwQYHdtg/7lt8n6rJYLtb30IYSHf8xBLijd
LyKCxDbOiT6zytcnpmDGGu9HmqmEII4P21l0RjLRTdUL719sO4yQNAeXxRF1wTxfdkquca2vj11e
Bi6nxYmKL65/+CmAqDq6/ZOEkjJXzlfPNww/bnYZMJI+EQt80fraEEIMK1PhnDxwSx+0eX36Frbc
nC3A8AEeSFl6dssPzyxu1M5fQJLb4Is/RhTXpzTQSUjC5cZQoLXtVnWC3TZLnvmjwjWVXuPDgRvM
ZzILItBFqGNT66xjI5LRSZMnKWc/2y7Z+3dm9NWMIWo32hbHx7hJrHMCCoz9rYPaX9Hnhey2e+rP
+L2JOKPUekTqIoPiSddVYW0u+vHNKe27jTu8tyYz1isyTC2mrYSSj5ZvO3yFXHx6tZPq0EJHlYgm
L5QATTM9Po3PrRB2zCDHZ3+bktjfE6BFyf+w1ycsU5jFAVeeMSww+3ks+46bjpdOO8kvFg0ZVBEO
b3fJfqJL8oaKK2NsilYSlgD3nhs7XA0W/A5Jx/DAGgaquJRJDg8u0PcNedTc6Eo1utCasNgLI2Vv
f8WBeXlR19POddDQFvGphkD/UgIJU8r3kw3qfcTDD+Pt699micnoTy0PWU0zvf6ELVO0eZI/dqan
XjGL+weo3ssEQCeQtmEvb7wSBflmeyfgLGJ9hrgU1OBdjRvfIhmq4lR/qznitvFYtkgEcTq3fNZF
1BrIpdlNVG2Iv5/Rrn3oye9DbPVYZ0kPwJRaYse++Ikun+vI/6FQE71Jb7kzQTbqwY7y50eOu8yv
q9pW/tlXFeW++m4/75H2kJxjbKJ/djDydg3CURvQHoItuNKLhofWYFkpCXSVZrC5tOOgdqRwnyf0
PO7ncivsEgYvKYSVpwTwv/lVmJeWI1e7NRVyzvQJp1noh6pF0QhaKLXjxGqiq04UcAs0IUa1HmL0
HFYo7tV4a/zlyVhy8nV483r4lxNSl/628kkM3efzVZMaPhDk4vfGUk16R41PtnH4LfDPpvaeJIAl
pxJkXmQAmGewio6UOWzmo555ZQuz0daPzDU6dmum1lh7F2/JRqa8fX+1AdXa0mbKBr/V33zq5gVa
tHIEUiZaCriJk6NFZQZCCVCcHZiidKPGhm+J3UYMDibWPi4Vgsbx5+z47fC0QSw+kXc2Az2XWRSv
9i20fGDAgdX2pGbPSdNhfwZBrPlypEw34/b/rnYF+J9H2w1pDh51+fc28SCruINDxLKFD9CGWRhp
aMrsq2woZEAJNiGojTZEOzcP3tkplDqKHypIqgJksr52idMSnwwVUgSnXJOu9WnBW1Xig2xVo3Oh
g1eL2FnZUAW16U0DX2R6bOFSttvT1jKNcMig7Ugb3XpMn8fFfrDv2+4BF8WYmJLfSffVWHwPgHG9
7NLShEbJMdmerL8MmE3owJffjd9aDEApz0kE5ca12a6CYkQ10XAj5WRjZH9bFd/G3MlaYCg/2MQk
j1TERapCmkIEiNC7gAhrqkOLedAZhns1Oc9Ism8PSdM/WGZsZjcuqF38hF2h41LiuF951ajo0qXl
NufwUqyvwSTKJldJ4SGNvA9fnuaahDdCx95NowL3kzxXTtkTisEvsV/o6k7CwCoGglvJPQfI8rT/
wyEgLMU4asEPE+GP4Q6ZzDyRqLu+V+M0PNo/wxahLj+kOI9jml3oX53Xt+eDi4uNBMqo47KvkgyY
ML7KW5pb7t1wRHS/+y2CL62BqxJ4vPNdsxu/2J+xPT9EemrcwggzUqftZwdvFCm1T4bYSroTAx7U
90ObOBBsy4GFaaDD8xZOUf5emp2luGtUNpndbkClIdDSb25S1KSUzWNp9/6IBpRi54y2AbAQNed1
4Q5gNOiBG7NS1oVcu6QpDSkovXddb7GFc6r51EvWSJJDUIA1St41LT6QxaXc+Q7rXREfut/zmJw5
EMSsXHuvrDsR7abNEniq4mXejU3nIIRlwg43FwGnFrGpNI9kUYsSFfUuOp9R6pnClYmLLwdITctl
/7LF3F/PuMghtI7LM/v/6SSQrlZbw4qUfj0MQo44AiZSxiMlwpi9xPcfHajrhc3gNQKEdK2YuJdh
t+YRbyui0wP0aiqNyU9xeTPIa+E5AYYat2+DNPjn6ecCSnZCa3dAcWaw/EA8BqzNt8oDg8QOwiPw
kwizGpjdoEAJeCPeBlbPRIOIXA+KMOKCvcyVfcK2Bbq/4DaG240WjAD8s0LeOMN437W0LnfkH2Nd
6rTjNyTOSjeFlhajgDaY009297r9KHZvE6+qc6Aw2hPD8yYFOBogjzeSgaEbVRM1DQgUfxFOPLUA
wkgxX30uXUFi46eo79GdEDFO0iilKLM8MrGMXHtooTrGXC8urUsXbfukCEzNZN4kIIiuTK7XRXre
tk/pqi0D+YAVQVUl+L1/0RlY7UX8PN9Dk1M5doMEP8DIwK5Bu/oI+AdLBdq+EomGYxOlnl6CVA+h
WoU88PcDNH9GlH3GgCLvdVXMrPTG0pMfiGNOi2vjRWZYqnwqy0HM4N8RQqmZuMgoxPDm2fRPX1vy
aBzG7hp0twzIpp/42onEDEh6rBVD8j5MZeUAnpuEYx6FHoAOQjyPtf3Nvo7Yw3LoXZxIBaKOPKsg
9n70STKy7eRqEwovkShW40Fhn2pzP16CBJz7xwCT1eOtl22Xp/tCTnHYAjOy28hqBez8LDcoIc5E
pmhkIFGrk0ks39TVLM7dHxT00qg4xV1XPXkPhhy7RVjP9YoriyBJE2D07dLCFhyFmnEzcecoRkKn
0QMZ8hjB36nQGQxeql1l6ZXwiSSE2R5J8nFspXPbgC9Qceq0lGBqSTAEEAILXo/gffG0bXRyfsWY
9yrfijIBrPDH0NQccubAYAA1icEUCxtWVAw0ph2geSfuBQOhj2N6FGAnXNO1phIhpMH0gRWRgBZm
t7/pDqvImFcICK9hTILrqrq+E5VM+c1OIl4MSRFYdzNNzXFrh/amfEfT35x/jGe18fLrOcAQ80HY
TDhdjN2SuLaoiFFxcaf69KQy1fk5yQ3sp+54SyRtwpzL3loyMoa/eptEpki77g6+xBMLMEYIUH7D
31w7hz9/mb1+Xu71TA9rteIYFtFhN6vwcjfXYms//p2SNXRNqgqKuiNTNxG7O+flODLwFz3f4Obk
LaxTJNhRefOOm2XLGRny7W/rcyMP1O+FIkjfTebcyDhPbEmu3SlB+JGswB5LhQJSxS+fSs5/xhjU
GuPmBUzO+epeCP3gcfQksyRkFZMFWMUBveLlFSu23fYVBK0n8Y8jGT49owxGRgGMEgJeLx/WaHUP
dQQi7g6hF76QUbHE+qVlA2kXGkNKAzzqQ8IcxcfQkjW8TL765xSWfxYIRkx4Rbf1kBV9VEOTr26i
XhSa8r2/FquTZ+Lb2vSFMCKcTiqQw/sVrzgArU0S5/vmRFTciY1xpchnn7PW5qfLCgAM/1Mv1LO9
qRi6HJC2LoZd73j6CwOb/VWp+nSu8BH+q2eI5TyUKgwDWY5lXN78rQqQ9E2q3tnbDc7nCXvk6un9
jL7F3hq3zkBzE75+RH629Ob8ZNIhnFk8Aq/ChQFmb93+y757bcKz0NLNRmGwc/+jOVcIHHlmpP12
kXiBRHjnewBSZjaARaFGU4dqSZpv6mX0SU0HSoflwlQ7/VwnIlkja5hhkjGiXuvZHQ3l7Nc6dRZs
btn4U3x+dlAAeWA8rAEjyD2fbqq4CP41stpJIo96RmHDtgnDcqMx92js2thMYG5f8jE+vPq80X1t
Jl9p88ovBrIQefYQcrBp8QsQwqmtHq5bt9khAzoHTvpBJnwrVo3N1s4TeVcS8P88eGq29SXaLSpN
rOD3HsLkGKpaEsNblg/o7u4nIXEFpLh7EJn6LY+fYswOQxm2bQHM1mhbBBpwG4FwxNUW4fgJnowq
EPkKzqny+qq1fb7PXWfqR92Re4cXq02C81AIPa4Be5144jeqJrpusPqQ7KhSeOSUWRnTlqnuMXZt
IhIvVLXCOnUTk3o/bsNRoMssuCTUyYC0FxmeZcWrees8HMvMMZ1DM/Kcqocxtws0fdBL2253t/yf
qgUD/7GNybkNt+Djaz+JzvHroTnOS6+jw5togJmdfg7jpQ2j6m6IAr6dgfrdx1xJ/kWx/j2D8JSZ
9sEbQKBf2VmDy4qFlF/rmsylmmvZkk4QvxLddf+31JhFNPsP8ivk+3oS5UtLMYFXJkkSO5hVFioX
HAvMPqHUcZkRmgtGQk9VCEjNyfhlz+zWjyiiZt8292t37S4GepIX/2nOPcnAdgwCKHW0XnWvEAZ7
fEbJQgbS1oN9ZaGlH+9s26XrOf636fo81h22f3ThpLLOQzkd7NT3ve7iwLzhSHc08c1Ehi2/g9qs
OXgUG5d2Uf0jqEnDSZwoid2N+7xdNjLoXsBbmvbz2ZCwLK308LCDCyknma+uqhRRySAWq55a5ja+
bHwLwgOBfEbOFYtXGMR+Ha2JZRzJQEn+64s7sCxwIzkkCArRrkdMpvRjWSKUqQziL+CkBc6lX700
VCDe3Z5CeBg9CrBJFLAJOKfB7wSu79HRbtwl4g2aSqVs/BlMZEILt/ueHnU5HRA1iXg4dB+QEBa8
Pqp2fbd0hDqs3+KaTzz72I7vkrUqnqXuQ79byehaNIijuVFDzXeoR8MLYIQHzYRdvinEduSqtlKL
VAjuKQwyTD7AqAUFscpSoRMkdfpONSOHSncyqZ9vQ3KfXO17ZS6NTuYHFf3boHH6Vq2e1pTmqYBv
DrGqpzfhf3EUzStt4T2pCdgZslJFQxjlaGuj+JCMRBUEkGs/FjXw8LYMzNckn+x/hp/7Lex++T6K
ocHgkeyXNZ5vbTI8tSeb5SE94GT2kZ4kAKBe85XZ2Gi5NVQdKOwLD9rhWJNknHdtkr6h2doGkbs7
lh+a41whvnFZOozILPryD4BEYkMuyYwRoAMnkFoAnd5keacxCoJBqNpVS7dVGbtQ3mzGy0RFo8gB
fYS1m2gHTacc9xZUdo07LGfi5vLqzXyMja2YeXMkbqeRoqxOFEpr89kh72JN9L0ofD39mtotZQW6
eRa2LFAlILoNVweqVAZey4/Qrqwf2feYOcguGX9TG34ZpGrKL0LdRcTUAJQZgBYKGgIS6iH6LPxK
5/bU/W1c2G83BfeGwG40fynxS5osIdzqQtHoa13sdsCiSm1GZ0RggeucaH4xw5np1epoOeZCL+GV
3z+I/XU5yS8DEiSc6SPVJwZU/9NNapeS0eb9+NRlMIcLdHOf0PWE7xy/sx9XQQOO5mwsLh3Uotfr
NTGpQO+Q3FDi9SlUGV4gglCqmhrEegiBgTwutYJ1/Nf46ygifxnrWQjtWMzN87dnn1fnxLLJ16uo
N33+FTj0qgl9wAq2cM6P0xJU50maizqzLZGEIoECe6uzrfEAihYr+yXbAF7G6Vfasq4FfJq6Zf2A
4YQXb1gXx6S7qVQvc+NhraNSGVc7FyfzOSsFra6O/0dK2TbgZjzUYoPJ1ZAAGrwJ73dpQpFWoLX9
a9ctHky4nh5ukWUFjpruHzi2x5Kn2FK8HBegO3uKgOgoSBNPsTu5j12G6kui6GSR/0l5RbyCKwWE
W2q5KbGNrnOrIfhtK8Ci911kbXHv+1XcjpjMGwuLeW1Yj91qxkrMUK6LDl8lK5bhZTkZS7/XIcVd
wM6GyMKngMlXbF8alnLeAQI6OojqbVH6v7PcigjuKnMW4r8vOUFSz/m9vtVhsxrOGaaOuKJZWwxz
BEqwUyacBs+LZJXEnY+xR70qtwNITCdV6xl/E82jqdMazIRvCB1fJlv9OwGW3/W9u7oAZrbeiKoe
woWNAzZZb9io81CHZsJhyoNeg+Z00V0eiqWPjDX1zccoMGxRykev6I5xnPepDHGp94t66/YQ3N5J
qu8a+SxC/X6c3gmH0Ck0KaCWfmsoGu7Grovyny35etUwpFvfjl+pKQnJ3RtVirxH4MaR2Dxvibts
cAbjyZueTfXatqyfZLwN+8nZchf5bSn2KKxD63az51RuW9efczaqCmiKOjgrBA16s90lhsGaO7st
Yop5a8tvPFvHWpuvWJeAbGsqsoCGF6yyzeQ6HP+KxHVR9kmJAQDTkyJU0Qmt7mrB5edYSIGyG22y
xApAOoQSeKDC58ewW266akfOSvlL9dQSknZf1imCgfeZLdLzetI+26eXv9YTL9Dcw7iSt3GnuQhr
vg9JNZwQpExDTHrQbBiPgYUL9omorTZDEfyEbYxbW2wnR5O4pEQr7GoCimPKK60V7Dm9oiH1c1W8
ptGDpheRHducMEkkqrURKRrOAvnwvWPz86jVj1TC3Wb8skd/AIQ+dTVj7J3vbf2ANfdwGX2HPQDR
uuKmgXTbq9QbiDVtJ9Jc6lE5TU9mIaiJ5E48PARcaSh+aRioaxMPSbEBHQsfQz++M4fPbVHsKtcU
sHhyN/qBfWAeXsrQtXJvtDbwmzBTw97UD0HGjucHACOVpdE7cPviUDNmVHv17somJ891f/yvhEXZ
CXtRlao1GZ/gw66lk0KxB220o2uR4jjIbNgcGldNMb0y6JyTAQR1IYMZUMLR/V6vljoik16FGlgI
df9WgQoFpBjagaa7dKZhlHH4ZLp9cDuTx9EnY5u7tcxDpGc7gMsczpR1z9CXy6LmSet5H+ALfOUS
9TOu9QpIItSdrg5wpYe0+dBUxtoc7iK9MYhiZoS1qbendKxlPz0hFY+SKKtbvTPpl6np/Hw2dLRz
k58z2+4GgJZlH8m4ttkC1uFY9VSx03tiV1hakVZpAKcK6qCJdkuwUYbi+2q/v1aTejriey2Nv0g4
0saDQpXuiZngubAZ9F3ODcS4cMi0dbG/8QAwzqSZwAmEzBhxFgMf5fl/1kd5XIgHutdpc99g4k6v
F27si4InZNhM31q4Hborwk1IPjo5t++dqse4gRB5GkihAnklMqss2UVWhZgpqeG7vWZ+2uOIEyV6
rVGlWPtnYLqoRkJ07+ymqY+rba260kSPUwUOPb1ig2/BfNG+9PcoaLJS8BTNNgSnDHptr+L1OEol
qt1GWCoa8xa43hHkbsfcZHNNAzlLkGSwsuGy1tvZUogNiY+2WoTMLAmU/HOzP7t0fSmFMPUjCd3m
CuLNwtZY6l5bkaHwE3Psr9oqqBeZqZat3bU9c5lwKGtuvv+gtSqVjZs4LmloomaxURsC3fOGleXH
9pPhQTXRVsi+BQtzW7nHV6jlnFrBBMFq1KD7sVkKp0Uu9PhOAto8boaW2GfftmVbPcYyaBV9rGJe
01jWNDOvAtaLKZ8TLRkDSWOpAapm5kXxUGZ4dULaex+e50iytjQQGPkepOTdXqU/+UkK7ZAcVHMg
+FGVDqxCi96Z60DwBFDF751hH9gEj2Hkim7LIDHoispqRFU/Zh5cVoh6WCxm6icv/6M96Y5sUV0l
/CMy750rtCp5+SV4Mf8jXoQLXkOYHWlrd8HC3C2ntBnksJV923yQZeVXIkLsPPK7kKJoHzSt9Cup
QEm1vv3QyLgM3qYUT+8X6f/z9o4um05kC27n9deWBp+DF7z8BdJjddsYkMEs3BDLT+jflshRsgI5
yaejowKNOoIpyAzCk9jhZqUpQLTjOh2MfY9mhSt5Rv979npihKJlvATEzOKI1UTyo8baxlZIUnqC
IJQOvC32x4YB0XOyjItqVsPwmG8WZCQJ1VO+QAYQNUIv7fqjJbMQDSuR3a1Cxdp/va+sxQ3E3ObX
QJY8P9sqftpDI69lFEUS4vqxe4C+hw87yUdha4YqW5OweE4zc2HfCPHYz25kq7uSWAS+1QIyPKgJ
zOaU5T/t4fh+YwHoYu0QsAruv3hWL6GoPFHk7dO5oW6uvQjxXNXENNU+8Q36v7v37HGZhEKjbsFr
9SJQN6TUwq0JZ4rbVd5jL0dtcqXbnzBywnjp5NWh+mok6KecLRdqf7FCm0fW/wdPXV02FZPRbSI/
NKiLGur06MznB+8lNf+m9lskqttrQyMqnpT0KQqQoze011CQgv9/fihdT2msGMTfF6Sy8yHZhAtq
yygRDrdbZ4k+u2P/JiMT+4jeoIKOMbwN/mw1Aj8mnMCqg8E2tTRnTuZkx51ocG4dnfTmFjU9ZrLA
jh2PDisk50tRTGKBxCbazUKzZEzL+3T5+EGLlUiTwfiQHKh0OtzTiPFdkWsjhMr3kdguwMd/FDuv
HcTsp4uIejsiFwc52c8v8+JhHD85abtO1MkiFf81rpvSMF8+WvK4IZqQmqq3Q+i9iRH1aLG1F9vi
JrcSw7InLCeUrXmc2nAz/hABEjcrndmGks2Tsiu/u662jbozzSPYxVOuKD5Di6Y/Q/xzx3wQQ3os
HHB4RINBymWm7CBf+jxSyECzXCuQ7ecDf1VlUZIu2R/9ThzxYuS1qqk6npILYmXLZ0X9ZbwFIHw7
OsTTFrGu1GAgULHS0UEO5UQbmbpAgBYU9Gk1URsKvnQAAV41iUT9SA4cirnPkkvN+4y/29isT24K
HCxkHP6AROS4HU3MBjYhamkKlf+AB4RJ+DdkmEvlGz1ANoetAQrUYvpi0BOGU2EMw5EQkdzqCqe1
1KjgzQOlTAgl1rsCGart5zLaE0805K/yrbYDX2k8v50FVSErhJe3HAwtoC/WwOAK+8q4Qsxq+zUe
prHQTg5euOhgKPmexmZoNmIjqo+YjYIXNSLfouRVa2pMjCzGGnJXGrMrQPtzWlHLDTr+a386fcEB
caVrBYNFAposPu80ytqQU4QdyNWaimO9vqCwWOREYD5n8eEPgxsvOM8/ZnpzLdv7PWce2cNDhZoV
aEl2s3BW/jrCkgrVQs7ck1zMrVuqmaZAcEBS/HKVO3vX+z/Zxh9kKWADoq3pSTndtqjBMY4B684v
N9VqWMB3zaTV/YWv7kz0Ztduv/X6corx6E28vv/xQagvoUW93rTMtgDDZYOVtgc3QGBWg1RHb7s9
SLCVwmMkQuZjQqp17iXskd17oUMwq5VanLJaneCWsYw2f6/rQUkIiaREHp8MIaq7I8ZXokeo6UNO
mDQrJ51uq2dAT+oxYqd0OMl8/GXckB7uBRnL9Qzm0HJQLTPAZIIvwku6Vds8Rvu0H8M/Smz5qPa1
PKlU6AHqgKcQ+IVNZLVPCrbKD8kBxqE9ymq7yaKiaULDaF+V4l5/mVvwaM7cQjQSju8Pms6fGg2y
2KNJDj12OtbdxcXFk+XlFWUG4M5yLW+M2JrUOBd6XMJiz6o1+pLimlm6my6ihdD5dWVke9B1puNk
Vb/LJjX1NGRTzbY/HO/tHEGq1UdFmJ76IAIyjZudTyWGwmC5poTaRt2p9WJeDywc84sCtMU+zbYx
8XRx24m1p9wo2DHVVStNz2QpXwlA4qOuNP8UT+NcuY7ctr244RrLmDDy4KOV1Ia6MCbmAyFc6s+0
kanmq2rJcfI8exRubUfRc9vPwU1NDfEJGMvBGPubObaxir3n3ig5IgBTfJd2EygozHHuH4IpgXKR
nFA6VtPiUhzykgzBjnEi6XG0s69F7IicSGJJdMJvDqzVfHgKfXUs1HrvCDT6XvKyvEO5wSxC965m
AZuwp97NTz0HkaDLvl/vDktFk0ITgOsClhhNPIRWMZCrKsayrZ41Iy+Mf/TOT/BhGJbfKym8unTs
dva7wzTVfn5mjoqQej5Aj/9nR224+q1QEVnu0AX4PlNnoyU8okTfPKdYSZMxBtyJvvyNod4Kblke
5ImIRz1tCAhxvtgNAQtkrfnYMZS6IxWc4Rv6FuZb5MPNosaRJF7QTLJ4Mmame+PuS8CxkQgtNX3c
ydF6YlITuWdygi1VCOgH3Ln1WlA0ktYLNaeTBhwUuyce7Kfxn98DZ9Om2WxcZFpo41q9iWkXhN0X
SxM93PhSQTcDzv01zvGYLCItxTqCBu5aOwDTy1p5Y/p58EPpGUru5XXJKTqXXqrKPuT026V5zmn9
MDt2I77gQH22xonWgQqsEoLzDPRu3H8hGqoE4lSXw+ck0amwIckVJE/v5git57uYhocHDnkJgx1n
akbfGaKrJMiFVDt+YumJAu/AD1QDpg7F3xMUUPgZajcnQl4yCLqS/YIh4ZQXjvNUd1kjaROYoOBr
SnP1KeJPgvpbkgSXaPlI14WAGAFBEigR/bvSkoeXRLwsHeievcf1OhH5RmPrmk9kGZCcpQHat9EX
KJCxLr7yyq6ncAu90db0HHj/Ib6DPRobMYVgBXEy4kpQQrRVsnZGQOKjQCFc3ZZav28Ib4G3HP8g
YIM/YN4KZXpSW7sNl3iKzprG5GC3VuIhhfA4iexXFcizUXhsVLZ9m3ddtfjbdQiqLotVNrrRVvk1
d+VPO392TT5mGU0QItGvzrFGYUb2YJTZ+cM/E2el07szcKGnZQW6Sm74JycTC+10PvwZuWpyuE7z
B7yjwNc2IrmSwsnEePsIWMilAShy0MQ1gabKdNlBatUTeUMmetX2CW/hEB05cHoVjyoKRtOVFY3q
PB6Unf9pEoqulFm6ZU4dQ0ww2uwVB+zLCNfvLym4m8/7Yc7bB3uL5AYjo5ppxScfzZ3BNo7zHMoB
XEgBMY2ervV3yT31QCQCzksyzuwpHr66hDum5u/9BCR3LaA07tvTymcq8zJHeS4wSqyr6yu2tlwL
NEKisHyB7a15mwNaWjNCNK5g1WDk/3+TtGzlCT5+Blpc63t3PahSneSXXU/jQ5YiVbuDNYTcvksx
kBppALJHxEfokwHriMyeSBYnzwJO4JS04j1B4nt/qd1JLw8gROkzopmo8/g0ocioEPzhMsJpY6S+
1w7yOgSsvMUTEXt1UyrHxCYATq3Wm1ULMUq98LAy3KwAQjgwpHnlFN7eUbnEpWqb0IxDs+gC+Qi6
XEHwoD6DwIUrZJmtb8g1ZOy5wPkR8vpMlTUwjvHopBaJtq0wC4eh3IwVKIRgaRl7xYZXYUni6YY2
PKkLwgJGBYD+JNYOSD2b7MHKJsNLs79aPHC5Dz7wAzf1wbD2dSmbj3Qmd0G9T2CM0hiacUnmwiIx
5wfXLx6P5SixOu9VyyRqQWO7cb47WkXNxtGpsgwmh9a1frLGYsQMdQmisXRzCKqakOpsufJy7HFa
kgVb5HW0F/KELi9ZZKApbzfqFbU7zI0R2rdMq4HXiwVJ/dxqMXgPz3rlErNEjWdJQCPEGjyBMBji
vvw+QyU8FTBtvzi1LzeuhwnnKLLxeSAGAa+EEhjGWRKbfhXP3JDh5+50ncQYC6tfpLttz6AfOJVr
tYDAjpsqP14EJbU8EfXac9wklYHeI+r6tL0sPb0Ji1VmmiwacGcie5/0Xd5MPY8/g7bcqOWUscEz
ynGPxTzV7I9DgxlqQCPYp1vOa4R+NAfMl8Yj7kq9fKqpuss2Hqk9okNcHZHAjz4nt8WmeMl2Y/iP
yMyksaIbF1LQKwU24fl7jnvPDcDjXLxKQV9pm1pKofQqllezS+opTBqLWkwwf+HnIl7Gy72NH8ti
nhHZyxd/kbeaPUIsUXNYdEWXP7e8Q4oqVb4DTIdmLxHXuyXrspsvqAPFAkSCqdBGdHsGvS2P16GC
vMpVk3BnDYsGiiq/EiNbb42H5xoP0gt415XDxg/cMOWVFCB7aEQcOACeMZHK8qyKN864ZdqDNZ3/
9K8HfSCG6h21+3JWAh45q2IK0XPc5HDRxb98R6kzA7M9biXge9xeZaFP4h80uzBHXorS9KKjbC9J
gxg9xuW1i+fKN69OLXh4NKl2JJmriwte6WTFr7TzIH0ipuYilUJ0pGPDlsmp+3OqN5ikCcO8SE9c
voOIh2b7zjhYNewy365GV/HgLVBkrwv+UG5GEaPzgfqix/Kj2Rw+59LZf5JfSyVnqGYnNbbMuJyv
Gu+9vtp1xViT0F9uSvA5t6cq2nAxjOL0ZgkeIUwkWyvbTQ3earxdx0CnEJdQliNWGBwNQWpw/MdJ
BbgC0cd5Hhxv6ccT3R3NzH2+hrdpUsSo5UqrcN6jYT15BeV/xwfCWCYh6m4kBPbXdhtFcGE5vzsu
gzilJDlIPJVWFGWo8rUN1b+tCQWzql4491cRaUaIfDzvP3Z6GefI3JMax2bfiKJab67RhAEilfuQ
bjV2UTTUU4yikbDuSQa1JheanbL/ZmRTjrMUzCUcTSaIyUr5GpMcNpFeSR4W/q53LNLgnuN4mU86
n7jF+hM21kI6/H/UpliLN4duGT9PCQe/tNbpp3Rou2FDj/ia0/oCr2pT7L44TJR8HOlLfEDbZsWN
BRkIyPK2iWdYfb6g3E7Som0Ed69pU59zjGfZsTHfszUJGHt+w7hW2cLObDGdErYajvka2NPElL85
GuyX6IFkx4EB4ywUgw9o9Yd/3irtb+GgRcEy9RsuEzq6bKpsIOteE/yZuHdQGyrWk7Nlj0Lwcx1i
o/OJ82O4OTY+r51CT62/747eC/+K/MkZgQClk+570PPz4RMg6eLDjvcXpPxOh8FoN0sOsO0Z+uCU
IKPyahE7v7pAicnLMVsiawGhZ0zEptEANavzJlKIz03zaSsJpAz1Xrv67y0diHNZr7kcZQg+KKVo
YQZUA0vSUuGY7t2yosEkpa0KYy29LM3YuCfCO9hu14vCARf0/lRaNoquSZRHU4pHlx5QKBAmdDTW
GYCKlLDnm+nHmwHrtPv5oR2NwHOg7aW/VF+vgIf1sqC5CWJ+NeIzk+RGedQ4QEBjZZYF2T/JZTWV
kIJvNSByS6kN47X4kU0zg3U6tY+d2TpWiRIwq+K6H/w5a9r69Ndsm9zD4O8On66WzZB4APDrSMDj
tLHHqVk4DoDDzy3KPGiWzg4vHiEKxNaff/AEhoJFq8U5Wk6u0CIkjSDqGf6m/M13OtkHGqwyEd2q
zQACUPMAlBLUlcb/RKxWq5QobKMWf8scEXps57dPLdk0NWpwEr7T8/dxwq9DaFReKYUuoYxM9t2s
D4bjBqJux66Xirp2B5i/pvA/bL2jsPNnnwJn9py3KQRWoNtu6mHwyyz7YWh/3xRNddfIvnUpuIAB
hUv8Q1k/+DZEnXniy/iNj6J8/hxL/rDIILV6XFkwFrfpNvoZ3iGgpelRpZeZ4SK9gP+2YjM0vyOY
x9HpopZtxG7D6en08sdufz9tGPLr7tyfLGKFvROV5eq9x13stN9s9Hxjs0nVRzur3VvWUJN4vJBV
FK3EjhXBYCooaeU0hoVtW/DjulX+FZ3psccFCK39X+1irQMFPwZekt/pb3JVK4PM039hR0NCEJwu
XgVVNXioEcmZYlTsEJJb9FNkOPG9XEuaXYI7dcljIvzdETo5o2SqJsdYZQicEM1Irm5Yq1+z1fDw
AD+bj95oDobHpHt/LKX+NHbX8+dbR9h5p+LfCmyyCuTYF+blqYriRbGDlfOXi92lgz+8ycFmX8u4
qsk3fMLK9rpT3+tD5T7iP75WC2ZlcqDkkznGvs6k5rQRAldAfJZLN9rUfmaMfs0/ifaugeV9UTvi
n2r4oH+CnpBLqv/y7/Lb/TzMoC7kkN6B1eB8sHq/WFxuH21LyJ0Bf1QqldI0UDHC5PBuxfZNDHbU
D/pkuy0LAvQXHTiu4XtRtZYhIak99YJlB/0PT8xCUgMWeZe31GxzPY1ghjydlgXRnN7AX8hLtGJz
JOr+3q5GZwpAWpIH8pBa3xKkrdZTedzEu6/W95p1XtFEQKa4OpnnAxyfoOgRibzXdVoUB6prvlqi
aqgddQTQ2MjJfvdBDiNkAmuVoVfE6cujBCAktJu+Kt/b85VQUP+aF11vHZUzPGRV/cqV/JSZ7NQj
zdenGm/9FQNDcl5UXwoCLAtOXPCtp8E2cjFdYXvLMUPyi+nMK2BqGgPkQsGXHZorpNE/DKerUNU3
yOXCmcPzreFuZuHzP0hbGsfCl1JAVsB1AAxUmuhgdnIFrVh9fprE752OLNT2/p0HP2zhZspG3l57
gV8HA//BzET1TyXJXDIQeWo3zWRZQnXzp6USRXKWAEggbHA1FyDP9eSZSwvXv7mmkPwlhgEP/oy0
+nc5SMEGxhVE2aqpKgn04oFoXFHRgWxckqQ/6ZWnFGd5Xlf5D6pwiMtdkZWdOILZ6KHrVp58FKyY
1PH1QXc7Bq8v6EywS7Q9ero89f75TlmrCGMjsi9/7zb6xvH1BFkzkue1H2xfBQTUK/OP+QuDkUuB
MDq0oBpjribZ/pEW5sg/NqTvMjZMMd15gEaK5BWWnpxc4ITsHYj+FQTqTu4wTnXIrfsAD3GtqL87
OT25E4FE2ddiH7CB462HxncmKkUVZZ9FyaCKYYlM862ncMnnC9XcrQHdRcZ1GjdTR4vyWQjrrJtV
bBwbcoQIt3vo4nsFjjS6fU4E0gyEwFKnXQO7D0a3WZtiZayoDOMlNP1Mfo0Qln56tLMV/7sWeXzb
1/4Da2p1FHKGsNk9rxwep0xvGSN1wzgGqSVw6EjcEkj14PuOH75QspmMhXB/Ujtc1dDiluYs5Mp+
kTqKaBZR29JzcdCS6h95SqhjFFE3kzDxPPt7KZYgQLRcQDlflLpM/+anqPlBNMzgTeM5UlwM25F7
8CkJqLImDpZE+s6ryo9drdGbizTtggg/xr4ftK5deqKT8FojUOHDGWPv5fZPt7DGSlvU9FI2DjLG
X0Hr5bdzm9pxpiRbOBDeKx0kuDjrRoUX8I2j/dm1JQ3SDufXSMgcmJcyJAOpSuADy4BYDh4KIUJS
5mr2yG2fNnyEuOm5PBCZNUdiUy1Fxq/JpEBKm4uo9StdyJQUyeSh48HuV4WqRaxS+Yy/e56tdf+q
i6bu2sfaiargiWFiNc8mHsEk0WUYLwqQe8jLTmlgYWbsm6gJaNmx8nVSRJasjz1vMH0QivqXsgUv
lJtcVuVUu7mZLW2tYpBbFd4qWzugI8lvgpZ+/ToU1dnB4BeMBPZfwHFCP4RhcG0d5xU66CqfbxfG
aZye5cD7NaJA2V3yYmBRJbs/lrmriTjXuhN+bkcnTwR9pGKUX4jnxCyrukMaEOsF10qnbY5iDEuq
lV60ZumzHqZ0oLhHozifr8mQ6lOEnSyshXZpb1PgiQEZHt6ywwJnMxz2vF2DvC4Sp8OH2SsA0faU
5viRgBkUwQ0yAontHZBoPLVnWpA4/EbvtTf5f5eD/iddbpq2Vjbz0EjCGIegd0mhdP0Q3ACkp9WP
on+LLtR/SBYCT2kU1oJTMVKjPJPhJ2F9p4EAP9OkvZOZGhA3ZsaD+en/aqux7BpgzU+Y9r6hrH7B
JPUEANJea+BZRRfmVf4iS+yixITDtxV5lz7ehY0C4P5URCCKZaflUzfUmlX7NtjFPw8vgJT0Gl9M
5Pe6yyJ4kKrBWjBF+RX3J6ALTeXAZtDcjQBJptdgDIyl2Um0xGD94pmrHP1f9RFvQ6Bz6kGWLXnq
mfnH/o06YwKE9V3RgJsXKLPOgM5T6qECXIh3l2kw/dkR5wFPYSXESXSYg8HvhJKvS3i1xzPpeZlg
PBZd9ottS6m65vYtV89xmJNpdSuqdZts4CBQKKCfuq9AdDBzQLQVWMDZrqIVcJEdy6OCVcMsfb04
WGfM5OUZK4AuM4LN+Ih/vC0i1rXl4m4vxNLqd/OhB4JPzhNwRq4kzMJYMxo8sPFqMrTpNkdY1Mth
iIejwbRkTe4euZ12wf11/9oVm7nZH7YWCq+8rbbYBKCXTCvTFw6LBsAnNs4op288bWTcvLfl53WO
vSHF2cCVJLgdib3jM+F1njkdObsU/QLNYfAK2H/8kJ9jhIeks8kh5x3GvYS+j1mT8TSP4VaO7UF5
HVL29E9bIau3ffb6ht+wFIyC5ICtLr8UnMz0jaPecESnGJrBze/FJX5hvRZOcjfzviHxzp7qG3gO
CvAhjUXJJt7JL8AKpsHiw9LvuasmIz9/rs1nrsD0y33BN4lCTRkNtTgvVo+U/SErpuGAk4BvAQMI
FW30qAFjs8wo4tuCBK2JsOiu/jJ4Cf09J0oSc/z3ANvwhFkwqSUyZUdiTqCiSVzv4lgHKoLoy9m7
yAHmbTUGkazqu685Ch/Bjwpk8UmOVz/8IpKfkK5jm+ry52RPvB3nVQg1Crr8sx70c5ZClLMBCoVO
N16ya9Monw/dBsbNTR7EIjLZ4vluEZl476UC/MSm5Eeq7DrUqytoW7sv5/u+6TvCE0vK9KkwoTXS
kjP2+E/Nhu7fwxOSlf2ERPrdlQxqBCbPnUQrHV//eEfx8UBWcRhif/4v3qXb4l/vSH3NUCzYY4K7
VmVq7hHZJy4mS3SkzY/+bql4B5NaV77aJxQLWKfrPQGDcQ2r5VIb++EI013jnDVBMkT+hK+h1o4D
I/gd4cnbHnf5mUxZ+7AHhJL+zXhKVYoaq+bwjG0OLmIsWckOKEQzc2ZorXfNfXfH3sGHHmzCtn8E
m0ysfXS4MmFKzF4FUW6ZJ8Q50PKNKGPlprm4tbIdQph1hMAbup10AJRM59asrZ2DYsGBUOM7IjgH
v8ZngEiVLMpj1zViqMTsme3rlc/kHUpamPOB7au86L4Bb7r+0BDCWvrL1q0bIyicAd8F3SglQtRW
yaUGVZazwgYMGhTjheZLIygNbHRfEuNQf+wvZKFY6UospiGHDTAX0IDt6lgow8ovN8pBZIEcdeOZ
Cm2PXz7eooFuaSauUuATH1B68nzsqqNBfRx3N+7L3fezqlMcRGAjlnNT70qhpNbaRnuHqN3cnAAu
940ZfkS9DYXVmD3AX6kIrD1+ctpb5wT5ANN4TT18fA7OD1fFk2LN3YqXob/q9lKTxirlxzg55CAn
y/wthHi06LM1hCMbg9k5r1ro9N6vwQIG1AVLScPD90VikZQU2Nm7VCaNiFuMxiX8Dielfow60QF4
OjVrc6yiWmq82oa4oqML97AsmubMyxeRyrTUiWSvWKZ904Apnf7sLuHUiYwUNVs1ZJnQR6tqnTa9
q9sH/xDzD0Tgdab6xujKxVOn4KcK/D+xAioG4evrjzNoGtuEf8Vk1CsOJ8rI94KWaV5sRzoDTW7u
4ypGh+6oqXRmhHXY8BzG52eQWktJidNSL3GL1+3C6Xk0IUiiOGXfxyLi1IA8G8TQx3kRp0JLx4T4
mfBDOAgVTpzxNB3WK40VXK5R1esv3Iuqe3SoT30QCwVBbgsR4CFqS9Qvq/oQcKaSx1BBMVGq8lj/
uQKANB9TaLa/fNQAkhlOrHnHePPicMKtPpR2r7JEZTlBXZPHd9hNH6VFcZdHu+VkMSQBHoLPlN6m
obOy9poTm5OtKblxLxh0tBJtM6y81nyXP6qDSiocUv/C8Ae+DfeeoWeRGk/ioDE5E3A/cDVe85NH
NRxZhYd+xPqvY4L9FzSC5LanwolSVz0R50ZO2w3F+bqaJfYM7qOIyw3IJk1HTk4XuieAKMa6o8lA
NXxzHxsHj4TYY36/aXICNBnskhDeVV/3hLdphXP2TRj62PxcBqcd2NlNLuKlj3VG16NK7CFB6YqL
s+522/HYaBNOxCRB1jFCHeKOkZyuISHoSlsMIHC2zUJJnGKC8oAmyktpJsWI2h+1zQ8gjk/yWvSs
E1UF+vq7eC4VB4fUt6a/qjzMqihHQBuOiTBfu5CWXe5RyUhRcyr8p5czh0B6hRT95wsZZM/o8zAq
HrI+fayRtemBv1WivuXIRhPTkpTOfhjo5qIZ315RPifhMN2CG17r5L2Sp/3Xc2Ag7cwM4Ysg1Xqq
ePzUuQOmbkUyMWHCZQAzWRxj6mNmimf1JUGfp3olmtEfiF+n66Ex+rS2jWf0BUP7q4/Jp8PbRjim
TNh3q/7zQgssjTzQIn8U5L7cl55Wy3O8+/yWACv9AtvggO2NtX+aBstlBi639OeG1OSz8ljtaU2T
6dibYf2m65S4G6Ly7MPyHMS0umZJgVGjlbsXjYZ5lTSb+6HB6GbG1Hd+3z1UPe/vzDVKKQzRbEkx
+5fp/blnLUzVYiPn2ist40Xsydj0XJtukoI/dghshgMrlM+e1nCCkz3eZkSqMlR7Gy2pxdFFw7tw
k6JM8YpgvSWwC/eZHmCqyd3cNkr9P2fmu4jiht6ovsh86ISnvKgNe2nGMNjcyebgvzDQ7YntxAE1
Y4ApkaT1mGZjv2DUrk6et7kB+640cIh7/YkRBOAdla8IS9vuHJ/uBuGH4oI0iWTjxBLcqBU9+RIQ
wG3P+xbE0JpjJV6m0Dm51+HModWaS0JKDJT4hsTznJvY5iXBWm+rgXnHLs1RASMVxPc11yvtnd7+
GvOrdbznG/yByJRQmWbqXmxKypOfRIav4INq6zuwcxgh52fAImOPxTdL237GSsOZc6Fbyej2kqur
bFHikWZFoJx65HmU6YHrXuvMbINlkeieBwe75xe2KFNP63azmpPpZoFtrzzk9Rl+uVA1wnmIvGkI
oqfiDTBDrOtyL9ANDH1xO7RyOk/u7mzcWwa5Kntj8piwVDBGUlYHVDw4wUJrnP3sTEc1Vrv/xnUO
GZUgWtYFOx4HsSjMbSLtUF6DHSwJ/SfUy2eDofVhZC8upFnFLKMu2sgGwCnfI7/9L+eZbWQqTQTs
sVGKsiixpZxUm8LJ3nOAyVLF9d64SQwMO4eIp9/iiAkILaqlBJpL3eYmemKYi4hAPgjgYVv7u1ux
uNFOLevB6b/cWa/vn/cnnJGBdYTT9I6d+rQEV/pOsNFdYLoCsNbVkEgngkwRYik23NWwku4yAKgA
6oyEG26xbhbRFIcSo9NVygvmZoZ4wbuU/jndEULl9IYS1FLBVyWldBgfO5n+EbAn5q1KhOGbwt1C
TeaCay8U385Fz6e75MCBnNmcNwQDCc7eeWRew26U0BT0Uwff9bIXCPTA5PVDNno5pAf7NnEsaKug
SdSotyzSkJDOhIaaAH7hoMggc8Ul6oevgEcjv2cTM0XucolQAjQ01s2qXV6GGNQr0j+M4yRWidw8
QZ2WAXZDgh7xJ4ceB1L+IcGlFc4VVaCQyDkCCXF9pEzfByrAuSZ3mQ8YvInoNIQtOvjiXjELg2JT
79DwxP9j5QqSTOXRCv8waJSBb1PtIdGfOJBDlkvevQWpg+Jv3nwzoZINsMyv/GlDYIf81Ng/0spV
hZ0Q++NK+HH9QN/+3J6upusvzWK4qWSZigzt2WLSJtsP1qQdfsN3wJU63hft1vzAhzz6iDKpnFM0
YdtqvHb/pOb3u5u0X9usM7jd6UPhRC5xWiehj4WSMoamq2iYRHJNZbf34aTKDvBLae9Qy3YM5Guv
yZiMehwPRJzGagqtn2U0P3vgBewc5s/WB2HMsgBLbex1J/ZLVjBEgrSiE4vagx9zdxLy5zaG33HL
cJyP3CwW3dKXPNXJrBe9YsEqPqt0zaqe/K40EO0yfHZpjRlS2sRIvMNbePNAHwEurQpA44XCP8AG
Haui7wK0n2zNILl2Xiyo5Ipnzr/SMZ+g7zltTcc12ZSYEw5qp9Os/l8pntHjKjP/r09EKst3OAkG
UZzcA8S8Mq1dUWWpba/hU0eQzUBvDpENlH+dwYwaIJI1tmz/LpSk+m72w6bdO2juE3mq8GvBhGWi
7WDiqD6siP0JIaVxjuvdoeRuCCcG1At+dHUMjlTQeADRa/HAirHIlcL2FNBgkPhquf0Y5mK6Nu+w
ZeZHl5EG6eH99eNN1KGjhwd3Txus08+iZWrFmJDxEd6A4ez+AS7gih8xWZeHH882nylamSDr8UCR
64/5obsp+Rb5p6SlE34fWzi1cRlc60RJGwaOxc/R1hNNmaAY1uqV7/gklLJFPYgbDECI35QBa/Yy
DabGtwKXneSuOFfLRvMVCV3EQA8Km1GRf1KWbsP7Z3QPfeg8D19a4Zxl5GoSt89apJl9DZhHmvVm
lFEZY7yijQn+jHfLn9MZcIjSo8qLeWMMZXlmJGsp8Dje6OfcyRL2AszFb8uwH2YqUKVxCxosvnh2
Nlztkk7myJ5t0DPOe5yuf48I5FS1G2VIia8lU3pdpUM76VvCrwQJxQDHVveGkGRcupt7DA0AOw2+
xULKkyvgmnRo1RMw2Wugi+xqUdJ40zt6cCfIawEvwuhHWlX1XPowqpkjIvxD0OCYGeMDXzc0/9ff
Dlq4LAqfD1rkL9Cuu/AU73EWgtLl7cNL97AouAgldfRur7MlovQ6Ikv9RpqSlX3mzrdy9nR3jQBD
PsXE/t0IPHEKZRwg6iHWNOwq6s1f5NbTjlZz7j7rKBlgVLhbxvBZJwZ6kvQ5Rwa+aoDSD7KvTVjd
35PUda1B5vzmDFTkalP6OnufHWEshRLO0ZdLNHgy1fLpltqJs7SDFGywPKkbye8BIJYffXE40u72
Q+zR10ypCZtYW5VPGTxuTxg5qLsyWVe3+gwEa2ae0BE86QUmP1YP75Y72Suwz7fiKtgSf8aibcH0
HVr+0j0+VHxrlNba7YMYQ/1I+uLz3adpAAynHrgI/uTSAsq3bnsHymn5bHqdxNlVcrtDhbTZPVVR
8PL/Db9U46wWMn6K1iTapvToKwmxUXTn9NSwf29wGurRsKJ3Jl6tZQK4waU03+CKkoaXnn7aYcw3
f8RcfwPh+tt6Rrd5Z2sTSOGuc4Ig35PnT0YOz6DtUjHVwUDj5GLqDN4MF4aBON8ryg46NrfzipJx
T7OByEakbpgV/dA6qkMX5JvT/bWBCKz1yE4M3PIo4C6+d829l45ZTaqjfVAIKojVTdfwLiNti+KY
3lmEWoqZdJLhleuK1hK1FaKIZ6f/POzWgDzxu11ZZMrStZjWndAz01er0qKaRnV4LpFOhurtacy2
cYx6tTORBUnFE9nFijO2V8lsO9O/fEtXNIsbrDqA6LXfPcO2IZHZvywDYrxzOeF1dAKBmvh1OvhN
RMlbJF0p1Yn6J1LQEX2XFORJLKEYrvcift9u1Qkz1FSrQ1BdrCXND6pR1zfsvs/Y6Di+VpLTmlXi
ArgSaeyKNcrRfVtv5/0RLjcoFFn66A6AtTOO38juMMYIpZxtwEEisFdpjzOiVfTginp3Pkp8UwYG
U+w7HYs91j7Xu1BbbAgHeDJ0p9ZT/825U8oDj8gNl7JrtTK6SIYAsFtywnYt5KJhl31US/4yokti
kNTrAVllP6AYInl91hk+M1iT0ZR0MbuwAwrpIOawP/Yy4UU+ePa6Z6ZDKQN+cfldS4CLGIKEZ8/U
+UFg/g20kh3FkIbPbhftIhpgTieWguuzpeRdT54rPKFpAfGiky4s7ffzrkYlOS8yUESbOTYiGHQf
BgbKyoQtGmCCUvDT8I4Eqc5e2su7RZiGCbL9rL/d9SwODnRbj36+i1pL6qTTNEH6h9JQElyQj9sk
Hr6n2FXuUSWZq+oPB9Jo6LZPNdOOx/hB8rMlABHafai6NYIteSUnPvGsWLX5Bj5Uf42Y3RmrQaSp
6UpasrRPqp8B2/CQvWPeLtvlqp8LgiuZ3OoOQYvNsBebuwKD7deOK0wg+6p6m/zVl0ENTpRqPr4N
t7YY8zlMwKXPzEpsiYauC10zFbDDOIBmhHgIpCoQPl8isf30zshowDIKGFCX7qGVb3CFIIlt33V5
CKX6EdMyZyc9STxKMx3KUXbO/P8oz3n6OsQaQwPU7/Ixe4n9DtUctJ2pGmKjHAMfiC9Br9QwXLGn
O0X/kbkE7Dxt6o66tVd448pV4Ewhj1EfMF9pDVzk+i42OG3stMY9ycgKSVJWbOBG7JBl5ZaXmTWi
G93Rjy5IQZ5ieXvekO2cS9XGwqB2KB/0s5WgL71pfyPzanLQ2f+7dsPaIeypoCyN1NE1Vv2uRdpD
HT6sbvPxe0BpjFS8PTsThTQtXzmIQjErTwN3LxTrI6MQlcxk/8IYxA0rAX8XZBFIacY9r8lRY3sX
97vT1vCY42hpztsJOENASygbaNhyEQ4InIS/OQ7e0vRRm/iT7SoBVqtoZnoRp90Q0heUAkS+Dh42
t1rGnk+uHhehHIfEHsahQdGLnjZUvrrfXOghBIsd4jDTYlcrBtrX6MzFfnnanzZf/dTrBD9SKXyI
n+iSHue4HqlnyuRYQrKOGGNqWPKDd/CUvqsgLfWM2WJP43It/P6pyRj7lcRCUt/3/V/CJvFAy66C
+s2DUUul+YVgwPAQo3+hmUbNcF+732qQ3ZFVLGD0gcw/4jxocf9UNxq9aTgaGfCizLZsS4hVZXiO
XKvRRL57bv6abYvzsDghGxQkFYytdz4YMIVBkmuoeu2zeQ3SpWz5ehBzpUdgNOyeVyCG2P6HZ8yI
dUBY2rzSv2TVvertaao9qdCAuHGBU/QAtsdkNMdHM6vW86SR6bFjFq21LRtAH3FazIsjxa/D7EIY
My7bFYcMBzygzjCLyJKvesDLszQ2g4dkxruEk+tM0SRn1SVs8Y721z3fuco5DF+JseofPbJn5pKG
mdeUtJpCJeMGPprsnoI76vtY5Gda9sd6yCRvLoDnk/g/ZOjq8ocszaxg17LiM0YqUM6IXDslW+Ms
cjpiaSEOcarGq9e4Nd6d1OPwStSketGJWdLoVGQ0K0O1GJ0Vxps3wc/o2XnjCmXAcChTP9s67cgk
qFWznmaDnV5Zm0kfcDRoa0ZAOOVJr85tMQ2tMtY7vJyTy9xSJTTZN3Y5uxY1NgK66E2Eq5ApBRgR
uYZWg0ky1qnqYo8I2Z22pA/dpWADPgA5Hee4wCLXveU8OGlOWx+9eXYEJ14WoXdQMqgjbgaLk0IB
joJTehfp61EcxZLbk9AlXzHJqK3VDC6DQHWhCJjKZqBMpoebooCdJiaLD3V6m90ScHjPdxnT2VVp
ZHIwKdQiCtFGeFpMdBor6kCgj8j/0BPRFgWhVnYYQscT7hOa/8C38nQXOf/AZ7BJ5RZ3jBSYBnwx
YS23fWaTMEIs0k8SKVmbhiSAuDV5oLYh7+JCT6mjTkyOfYo3GnspCFw22sHgiJfQyYQmsu5Gc+Ec
Xs5TcnDiSA/qGFXcmT2d5ChYEpZjdFbaZlLKCvE4xwhJ1JRqKw5in5GNtFX538yKO4ZI0dFBUnXf
HRYSP1HZKt0qJOEiiwrPwBeY1jo8Z9gqv+bkQBeFVdfB09ZgZYRJiJDoNEsXTdxTqa7I9nU/rTzo
QvHjAh7uK6BVbnbGrvvF2ZTkUnvi504sQknigYjEQzBLpC4o0qkKsBMrslqelPXL/F7gNOsGRBAo
HMUuTsNHTV/k9oyEu1IZgziyGfXVaOWRvzWUGc/wv7pYwxObIrtyzFrOn4HbFtI28uFn2Oc9OBqH
iMc8awPB2VovN2nIYXnzgPNuglTj6O5BQ3L/8LJMnqjpeRC69Tzsw5K+KIWUpwW5qpNB4g9s7jmt
bZglg4qQbtfX9SC+cAeEg3zZeI7OUEAjHGNtLq7dAtus+7oXjvlSWwFWfZq7SCcPmUsKF0OMuI6T
hQoQBLvefZhLOK6DyVhcXu/mgo9N5BZl3oEc2nwOan+iEzb5la4bg8rZy3ois9WIZVQQ2D91kV4T
FZWMstvi68WpZs61REY2htQMM18v4l62f9mFxydEc2Cw9DnAOUOqMY6CUgBR3WIn6J7jG0ujoc8o
vhLuuIlk7oLOD71U/SdhbZYvPlZMUZZBdjJJDKzvJpRRRmOPFxHCLI47yvaD2rHFWzhHUi3kYgKk
fkdIb6GVgACCRbZdgum8ez/N90LxiY1ivYiYoD7BfC98d3UkHrGGr/9ksUTcEZwmscb7fgerwRPf
c02yx2rNbC1x3Lb611q3fGgxE9U1nOjAOxNl6VJt68NWT5a2rC7Nx8F/6vZefBaLZhc8uTf8RjIN
vhxZapUz9iBwZQR/Em4OYljfBq24LECn9J4A9AQLL4Gjc0kY+Wr5LGbWxz1vneuQpcly7aCK+jVs
tnLlnlAxwl3DTMewiHNAGE7STnlpYn7a3fqwv9YrHiTGq2wiSL2CFpeS2lPipa9HV4jHCjJHKmMO
/hMP4Q47axW6qicyNDhelJnXOmpud8g6RBYW48DIXbmC9dTB1DIUO1U0VJ37+6uP7/uxb8h+H6Go
BAmQkUc0vbhx1dSSgSw/CoUMZN/6n50QLzZwamn5WEPb16NwAakryqfxuElCbFtOdgOwfTsrZ+nR
0reSj4kmaw5nFyWk+HRcLJzHJGomOvQ4qmndFJdjuhge2N8ZY/XDgTv0Nqo+L6OQKJ+aNe5Hvfxh
eh9wYOQ776Ayg3rq2FpDEioiIRqO+re8dSvt92oVFx76rI4GUSVvHsxBtJnY0ne7BVXlvWEaSW1z
aMRV70DHRnH2K+9sVDz4ELpV+3Mz1ApReL0D1W6g3K4M2dEjH/s2ffnKMD7yi+gHh7uwGu8V7LpZ
x/q55EQ1nq2bk5sxtCoeS/+MaW46KUrITWmivvFgmVo02ApsqhYp48x9QXyX9fBjADOeVZRSJHg6
SQ310auHwG/r9kDlHxjfQ3ARCvV1Oy6RJxw4BSMkP0EhZMFa+SOf3Q0/QhFu60RSVz1HdAksP63j
J6CG5cPcWbH5paowjNkmAKaMQDSbYDOj70h8Wc+pOhAZ11FysXzS3HL764gr5opnpamY0cf0P+Bn
vY6ciXTluGdJEtYAHdy6bQPiOfS/W+dOFGCU7+kYlOU9bKtH0Wn65T/16rPmBfOhLQ2jR12g1Erl
i5HvspreygZOu1mGg0tbTIs5HHFHOdB5xa5pGPajbr8AFbOfvZaILphm2v1fSzjclU2aR5xOPBYh
i+MMKBcI+gJuaxQExa87pnR1xJglp47AYvS1iutKWnSqUZ0GPAKnAbmAt3he7BXNxGTCbJmOPvb0
m2NU6gtrrBfd3+9GwhufrmEfP3IoHuFcM/0WN27gOB/g/5CPNTbw7/YFtWg6uJwJAOXpb67mUiRA
EyPtMMIW5x1//cR/ReyY0QWlCRSBTDkibr/3X3OalC1T18OXUXxz7xPx6Q/Zsx0nYixUCDCzq2GL
gig4x5L+Jrt64t6f9ml1LKx+c77EFV1wNei+1Tc4HWQsHdzTcldU4s+G/h94va6JEjR6+45Y3N8K
BxU5zgY6KWMtxGfhbjf5tH8uP2OQ4wfl7MqFe5jqSG5IfU4fkIfjgPTwtXx7ScfMIF3KiOu+FdI0
zLv3I2PFslJ5gBFrNGmTo2se1R99VRP/poVUZ8VQptfger3t6WF1pgZO/GBXuDk3nzvGygSiJBKU
gtbil5V/PLNXdtNnxQAEhWBRg1ZjHLaCFTX0Z3EKBqWEi8W8ThmkahWYutRXInvD5mh1MWLsXPa+
DNE6l7LabU4c6zA5VgyEbjgOYDdvrY3cVVrvNRygNmFht+hDAlPSBkPEi3S2Chy3BiHdB3CPNlc/
bLUbjuAEYwtwr57sEnpH5NlU1L8e/NtyHzN//B1L3FFrK2h1XWuHqhOO/JpWIUiqJ7eMyKfS4wcx
FEk3KLfh6R2zzTGJNFF44z2LOWDfG/vr5Ow/FTs1DaZYclnCp+mzqUnLfi9E9sSvaSMNz48f3MPB
+xvBBNcszeL3Yg6BOrs+kPxFwHeOf17rgfjhyBIO0czMw5vzhq/EuFacKQhoRXGH5R6b6uvqLQqz
VmtygvGoKXsr1oYAT7wnXSeLXYSc9WAotu/kmM4oPW5yCymScIaRDJubF5GXmR+jLqPnZLOvKY2q
zWLdL+8TsjS/af64tul8uC2nS4bXpGTryuoRILdEGHorJUIq/LzS0XfcKrjaXpfGVwLPQ0IaqOcO
mKZmSDjMjh19rtI8uTOPakrHwyF1cadBoYx+WceSTTraxiPcWy+mGqWVOOc1JbRIuyxdcB3gmORP
3bkXgQMzGzPSqtY9Hs+T4OF/qBFxavKUHaWiMra7DydZyfPbZpRAfEEbe08uNfd6W/vMNPuhDnbP
RAtv0HBV3VYFHmghlqlDKR1/5FSdINGhgiRPVHBNBYgMrNOG3M/vSXCCW8HC4y8V/yLu3zniNe3H
qW2j9d/ImXdAkoMgVGTSZYaGO53yzevDNJkDnC2mqYSoT1UJfT8SEN6ad7vPJ++/iNio+hCmcDEK
mcn4A0zIs2UJo0koxaZs/MBqjWkMrnJKWUt2cJkcWKSoV9IN1JPfU2NpFh9R42QzRuWe2JK+JKHC
u49u8iDURhFoAz9Ra2jnkhva6chxJayWXYjJ2DDUv5URug6aYO4crPd9hfq/qr/EcOUzAkM3MBj8
zjyFp3rVUHTgm/FtcDaXCl/KCnF5RLvTc+d4qVzoTGuC0/4vXA+zP46RVJ0INAPFqYkOi7ePHm/T
dldo18Z0jJGI/wDgVlMm53ik4dJgjPZZMffrU+e+zNtAVURVtnbqkMu0pUqiYujPqG60P666M7/z
3fh+pEz93Q5/OcRzSvdBAuVOkmpDU180pWawx2Ni0LYq0/3kEhqaMuiDmKFV2VufDuSqnXHCKnsF
1ASSZZ7PwF51HCvJ1mdWxQHexxsYcLaVHAhMjr8Yx3YreMQ11PUw3dilYFBSpYwZf5h6MBvmqU+O
teDv1cUAFHBPbat/IbHdeX8LMjmg52U60leC6qp8ZGrGd3rt6Tw4MszN2xPLYJgyiC+lJQY3v1s4
uNHSqnM4hk5OhkWS8av18KHw90mc29fsRzcimjxkUpreyIe/dPBPvjqkI35Y+QpABskf2eyDT945
mRoJaFtdZACW/48xJuNMobSnAOC1NnA95Csfu7Tog1J8P0A8Nx3v30k5RW7zpTBuVjVUoP9laemA
9MvsURT3EtMMsgvYHO9Z12NJhUeyiI4ggRdat8PCGm7D8JcRAfJg7AqPW58PceHVNMjHjkZ9n3EM
tPblBv7ZMyzg9PSsHCN5qjNdffnMJ9sd+YGBTF9e3R0f8XzLUTf4HBeLkaoaYOhlt0RhQdtMQ82c
Yfa6XBu3beSq7QP9u2jh2VF2xSbNKNmKw/PMyOuy2VgbYK80FvBdWm6c0yanpzuBlHtoWDe0m6zk
tN1wbssd99vI7EESWaHHiLGFDIJyIuCRB3WnP3UTv0j2KieS1dTJEJ+7pItZevd4KvUna8lE74qS
Cn7FE3iotgjXIqQ3lI6qGXyE3sBE2v36FTArF/oAPKEIE/Sz9QQcINNAdR5IgcdK3ZUxeaS0eTGQ
oOquPTVvTaYZiU/0PVUInT5uw75C5Br+Mt3LxFWNKFOjBblmG3RQGUvuEdjuNCWFrfs/Nk92nnJR
TEioRGZ3BkBRI3O5DEfoKZ2YIX0ndREm97DsIA5fDmQTbjRkRjDrmTRXq6hqfzvYM+Vafk86BU5M
bwyQ81pMC2NZzKERPIBBy8byhKn9RpIBz/0+92gUO3Dz1CrM2yp5O54klVYWIihUMYTH5HWuzMsd
LXE8YgeBj9iGNMQkWsaBzQwKcdse5mp4lih5H97xeSmYKoEOjYzVZo0eXuCxmBFMEeyZvJuWo5WX
+ARyzNXi4jFyvUpZvH9vlV7IHNgePUkQ0QbEaVPuEEleKrVPaYUcU8YZH4wWAhHiiH4wxzFCRTw3
XvW+/iJM661cz0AzJHjSdhRpcKiNONO/yJWpRkjIi8mGKl7fDDnwz7HyugpJLJdBhlPYDWOOvAXF
reca8cvtDvg0EHjFIHbInI91pIpE4iJYzq+R+0wrN6UoAlX86JJmsC6wDwfjGPaux4IEkuoE1ZYX
p4U8E8r+4nFTl1dbHELUSAfRfz0hoE5A6p4ppjMZFTBFaNxUJhNmObaWZEr/ivxvIiSa4xPZIKPW
pxWORo3j3UrWxSEuJw+5xFU2YvHWq+1AMmhoRh09YD5OVe8S6tN1WTWnviOD8mBEizekebarpQZx
zbiq34oj5iIIfEjedIu0edEZn9vc5ZQXELJsnMY3TPXvMpaqeYnaFobeGD7dTbOoqgfI18whGNvR
GNP62n29yCIPyszl5w9jQUWsCMIchzYZLgKdzpPV4sfEB/+3Qo6FcPhUf7Rl623CjI99zGTCJAa4
DO9tFKcOTmU7NvGqOAi3XINEtk4PdfUDwlVMheyb72HemPJJ4PmGd9eHKcWmjANummGnx4HNeqWN
/Y2eQ2mAL+AuQYt8w+VT/kl1kkQ0NG8xXuTZhSf0XR2OZcFF2QTqw8S8K+CIr6y8zVw2JFDuCtju
sVh2XPnrfAXwlwkb/n7dS6RB0hnaCBMPWzhmaEeBJoFoXbP7kcU3Qdfk4N5AoUA6mPbcYTYCOckv
BhmAnpK0Nhaj3IQbide4d7t+IRIr3xaAlzbXRrIP2xnkxhA6LYrBcJHh0jcKJKKnfaoFNimQpx3A
X0eIt7KyCoro1OT9qnfPOwNKKrevpES458HdjYo+/U0mhvw87xVtPaeDqwBrYGR3EMRAnLSe4kuW
yNtJHGXOA5gSyOKMNYnKHsq1iRl6CZaKoyTPjSOEWf3YWr4lmiwHktKnXSfHOWkzaj1XxhSKsBom
1kh0vst8IscZjx3IU7TYNePtN2nfk3VHDw+WLAzRtZgngPkmOIZIt5AfwRn7+Gmd2qZTpSfhieQ9
71Cy/Z69S9ADmJ3VUakGfTLv58zm7lYyNs6+p7cLnZBB8jRSaJ4pZGBvhMKXH3owB8aG0uv1phNc
UPnpdW382tsIaol4pZyDf83HKZ8MxBfBfX5ywCVrSLP6RZqNC4WiioMVfkUaDM4xSCrneAXSa6fn
kHeUE9TT2JWPvKvLN6JYr2Mmn2HaVOOQ6XZNebP6lQFlqOAU4T5SxPaCmzVirlBVTJI0ugR8tAx7
yoGLU7ObcXaIbHAacAE70FA66eD6wUMRD8j7ECZIFzkkxwUg5HkBLvXwqzy8Itkz+2DiXnye+2m2
Jx+QENRKQ5OPgeIdd1Ja6bI6Hh3usUDiaGbWsadWEkMQiWDV4clqGFXS1+Np6c4j0CCjqz8I5cMR
OAcz2y+IPODlHRvGuO70yPmELITPs4P6SUcHP6vxQKzgU2KsL4XpliUKlC6ejrpDnrHOy6ytGHzr
5ebCkHHOuOOQHbvUZRukppZqLc6YW67dI2rXyRSUU1VrzIBJMnm64013qw5Tg9ZB5k0Wt+E7iNlh
4nAmdDB/7KIijMz/Ue+7GQ+tn+4D3xEUySkZIJykgdE/ymvbtLUrouTyu0T4ANkfmfG3jHqRAURF
9pahVKWRzgib/lAS80+WRYfB5oRM27/E3P+3aDxJ8CA3a+JbQYBOPT+5QvvZCEvxoNOwLpszVJNk
gpfQZQfB0L7yTVjJSPWo2jnL01dpvMGJeCj5wcPKmSggdnl4T99AJE5XXp2bARg67ZPkSMzkTBxe
CZb3J2jkBLXdSROYtGZtSnHhyac8a2jCO0wa6A+7PZQ9XIvpxL1p0rKTSWYWdioJcpGqz3LXrH1n
g9QP5RaXPhR7cIA6UrcuqrRpYCGsbwhN3fKMV38Rt1Ug7mUcaU76dc4ieIVtgrK93A9SFUia9aCp
VM7ikhhSc7oGFw3EHjqmLi0Xcjt7HrKIE74yJtUJcO1nOTKjWB+aWCt+SD4xTPMa04GgVaqDgXes
5bKSXb75GauVN85+riUAWvgHKbdJVMCvqFJqKRVgIYYz+Vc7cW3MzM43k/cKVsqGfolB6rcL/Dnn
ZNZenK72VwiuktBcszgGLqKJvmOLEancap4IOXDqfIdW5nmPgKy7mWOvKfiQ+geM/Vb7GcfR/VG2
sseUgBATedwgWIUqmQ5kK6Nmntw2JXF2gNOuTOfDeXTZNQC5ZKvQOBR2vgQa4uu01+O+je9VtaBc
vRpxK+MizgDn+pNk+5dCSzrOVTYThJrRZ4lf2YsH/kaBSj/1rtLIFirZM305GmdW7YjMP5uQcD5l
3aKKNexF2VbJ0kG0cQHklaApoZa4wbOZ4PKp6JJ7Z9yR4TcyNRvhQ3abu6Nr7biPmZxSWrdXsuMb
G4KzEtOOYjU4CzobAnjVq1fz7QIWnNRcaloK8eF77pxUiBWEehmhSF6F/acBo0+k0wTGafjctukc
wXlNxbGIR+dxTNX15FMunQvsXwQT0wTrNVF9KII0+DmUvfG8CzM5nbXu/e8SSGp/Ua21UGCX3sgj
h9hqiQS9mhvM01Bi2Ro9W1jdEINrc3h5IVL0NsZtGDVeW2TZxfpk7Vqz2gZRPHNEBtkDDCQ5qD1j
og/qJdni5rmYCHBB6LDHnPeo1bsigtS+3flZIegZUEdJ7vDBK19mCxGsHieW9pv3kD8X107PpIyp
+BxVjHN7hITd7J12t9idTNU9vg6By2bX+fFdJIYoBjlToN4V19WPyUC2n3vhR5anQAf1a/Mxdcyu
nD4jinsIwmQ0nce0lqd0Kf0afF4Twt07wQ4wJcfEK+WFBFrBrpIJTX9SKJEQxvThFVh/ZvXkFL9+
nMX0g4+5x1Pwjn+SCe+yx5a8dz/j1+QMIPx04H2hv0hGEFJ0zJGOz6qwzE6o2geH/ZaB86y8xCyF
LgYgRV43uPB5omUJrK3g6KfbiLdM7rLU2brguTUbTcoKlCuRbtRBV8OskQiUlwVEbXz49xFYiXck
QB63zUrSNr8PrSzVUHUH5aNo/fqCVQTglmF3foGyT4kUe6EDpdcrPcDp7GXUaxmYXUt/V+G0W5bU
oQEGfFZFcM25SIIbNBnFnXiu7xzx73qNgCU3vXlGtIAKjfLS2fnzNwxjChU/QtUwN6ZxKlKmSoYx
0ET3938aQPMdRuPwCJ5N4HaVlpQdkmRYpQe3LMsirDITbme/r4G7duT1JVDTGfy7uNJo1y5OTEc/
RY2w2cLmaOdHhl/dsLlXbKUiHRNG1HgVXYfj/Us/Ix+brXQJkFo9DKSMcaUVRY27wuXk5ldWVhNl
7mC/AzDW3S7cNV5rC4tNNYA2e6Fj/5iJ4Y+nDcda72C3VM9RXs2yZHiRF+qIHKp9u3cNDZKVv9qh
8knPev7zWtYd8dFNZ6LKtAbk6pd5ROvCt61OLv6GnFEa1AYnMDi+Axz13gbEnSBi2VNGwR/DwdDM
r+KHWhNrFn82RWgLoSfKCexbNOJejP4iCc6bulqx1PjmbmlvxN+zYe5f4BDu9S049q90zAjGQXl0
bYeQxh3slxheSp/QEDkkj4SyFcscrbaFVMjlKA4lLRYSOUIgZcd93rVwpH3m7wrBSL+KaBsLUm+T
p02X7z03Vm10vQDeIbP1SgPKCrF/Py6YAWTPBaotZLVbCv5DUA5kh+UjpJzSGAn3ob7ARAJToNVh
IPWCprxVGdFk2P8xKlX55p6jwaht5iihn0xOkN9TXgaQxZJ0v/gksD6jssn99lS8hGPto+1qftlg
RDWLe89Fg7yvatgBAJMbgfU6M/WKdNEjnYBWdfA4h1R9XiGec90p40oF8pYbGZEbobHZUy2boT+j
O6YFq8VJAAQ3Liuo+ooePM1HwJrnrYWvx1mWDCiYMxQdAzyzpuDkRWD59ghqPFD6Q+ih//TMtu2L
0R0YUIUlXVcl2iz0jK1SNIQFiqPZRZWKBHm3QzxaV4w4wSRyB14e1UMaPCYwoUXWLtyKqQhsvlA/
VsXQ7uZLHKillU87+h5rR7XPqFVTNsVHlI8Va0jsaN63w/rv899P7mSYmMi+nuoIrMcFJKsSCbOL
gkgW00gT2ajilmR/xkf4QZzhn29nqYVVxm0ymGKslQF9ulS8uasEAXOrCPlskbq7xHu30pS7EMO9
Q3XwBOnbsSDdrV+Sh/d0Kf6I16cgv58ZBmdev80qZSjsQua9ym/Bbn3oWvuctOdpuuko7d5rsPUJ
xYOlGuGC6ZMUF4khMEc+L10smOZPDT1+tSfKR8QE/0KXQlKJJHxKG/tdj+/PopxwTLFQZ+SrM42r
f56grbyufpUwR8KroGjSt6UABDasT1lYlqZcE9OgPHGMnxf8Y4iFL7JJgbdv4cPKPRchlm7t++Jg
eMka3jXyYZorDNXEsVCYMPLP0CnNPFqW8Vb5s3P2Gi9Ir60Iygt74Ouog0gm5IBzpk02IDarPRdH
3k3f99ged80CjzNZvOexxRc7eKKEsZeEpYACrtnBDePNqfFNGnypP3oWjV7ddbaeswei0+dC3cfQ
8NFBZyPJpyv3F6kNjcGOhS+VnTVnJNq2ImK8zBBshD1bQ4HoPwvgr2nXDd2JOlB3bMizQlSwGj2D
FZAJ4OOLO5V6RLwJG3kDIqClvfnUlsqwCr4Eta/tZJNGwOscy3abIwwi7BZzWzUIPMBmcmRZnBcv
3EJEr2JWCMxtqGxtCaiR6pKbSRX+hC6cjICTIDJnaNvn6ft62t5qAvkZ2vyo1kWPQMcZNkFyc5Wo
LvG3rlAPasR8UgWhxDEPP3DG/jQ7uIUGxy080FGHZUStmCU4oe1k4WFZ66sv+XWeFlByAyy5JnMF
j0zyxJAphsSpSAw6tRqqsoytim5n0cMPRM2aFc96FgDKGafwAu/CtGeWe2sVk/C80FDMirGeJwBE
tVK0Z92WoRGI7n6X6CkFJTn3tfRUX+D9P4/dti6LmBW7fx4Q2L1jmNqBRNoN9mPI/oHBtOFHRVph
WgUJXPpY6x9QBDDvniKQKlZcrtvqIvJJhGj+cGe0h1LirIllWgxn4yOWh8iH/Gzd6c6dCtzCPZm/
IBrWW7bxwnDSNX7hVRgDu3JQRVazZVcuoMgAcdBUDcbwFEoIke+6UjiBzmo8Vrobgu3NAjVSb8jU
Xc3H6mfjxxBkvxo1QWS00nEw0UEpIJAMj2OAMwZFeGPaxMIJzERCFZNrL5LEx5MP8bLiPimqhyw/
WsDke8lwpmc4ygB0LikEwtzV3qusKorGKTvEstMqgL3hoMebNWowO14k03lUTl/bbkvj/RhIcodF
fTbsxKeYV9fsEGKCYL48KVF+VlOMHefT57p5FfWTivt3zJ6aHmaC0auwTSZSxETSxUAOlZhFFHET
jxl9QeD78F4BUiAejJgWdeLCrptc8ci2hUv0nsjFJPy6F65xsowWW3hdGuY78HRnIZY7t34VTHGG
ZpV7nO6ywx638Ij0YWDmHLZPyXS59Zohf26tjHK/ltoHb1jaN4QFJ7LlwU+kW9DHz/iih2YZrfTH
/8MRBLAavdWMLkOUJTCDmZ7C4Ytn+4Ce+gYyU4SohYgt5KtN1dDmvTwWUZyUwwTNVuN5q/uzMr06
rcIl4ZALw35+lcEXLnyhW2G8F8vYwbAYOOTwB7jRRHc9jvmaFoIWanccjELEgbtaEGy5sx6OjAf3
sGkPGF4G5xnVtrVks+j0nXHUzcFgVHhCoTe76vRNAWuVe9oeVlFdKuNEZ3700UaPnOG01a33L1iY
9Rkwlfbpsyrayk0r9EQGvXqU+kvDjff0Mh8fPyVNmmy/S19tdPQLiXvHqcVtwq47Hm3HSuH0vFkr
J2T8w9ENdCIPIz0ItxeyQ5D8x4sFu6m0/htzxpkyHMcju/1IlwRtfm3AhI/D+xbTmodjQVqiW7jX
n/opjHwS7U0iFhuxCkzE65HwGoSChnkg3X2xQQNUdZFAepy6K7zg0b4mUJH4kNImcm1Fix0jEFep
1y8aabgSlTYYWFnY3/T+4WLYv+ivHMoLPAlGhiuBUdln249gu/FZPczquua/nDQ3TNtx5Kmvr4Lk
4ofA4y3UeIbTZx2+OulVhrKr3NaGIj13owezN3GjrR49FH+BTjckI0FA4P7F47o38uGZi0oKjAh8
irePqmlEGEuoPGJ4JQo2AIEIyIu0HNKRonTRT+DwaBDzKHvIaqQDFb3FHjn/x6eopa8XXKAvMYNo
cpjC/itTBz/trZQ3bcetpUjetYXAEMyjZUZfT+iPweyeeA56eXkUei1FbzCs3U3T9aTPYQUE7xvT
zze2jVWpxODb2dZbod47ti/SrgFB+X3/gykovlNgGSb95uFQiOXMA6DGAdlX+fYs71MVIJP2PwNh
EGnQQ/ax+AAycF2TWiuLjyuYvW1tJfi1vSjJx2w7F2/9Fw9gGxZEr6Y9Qdu+Jlt7iD/7dmkqB332
KHmj4J/OhPaSKaOPB09n5vUvJFX3h6ZKcjHlO62f/SIG9cJFOLQl7HUy81RjQqJTUJzpXCqR0VXi
J1Zejr6wB2Ngx8AluZLRa01X4sqBf5sJFkPTqOfiVvm+R5SLBSx2brBbAp3MpbLxpwAt0X1xrtMy
3GLIv2BdtLjZ6N4lYofxf/A7I/0YRrCqs7EO2Mjh2KP61BSghHIwOxsi7+fM3edjlSHH+mRpm+2Y
C7yFxhsuxTawk/jovPRtQL6XvFzQptheLIpR58pSypM4l+eh7hD66lGuESkWctgFLjqgaDbp2r0P
Ql2EMQge0DHzHNZA3lg7u6Hvg8k8gQ8CyMb2NSnoQQJ6hsHmv/lTvcaq5DsvDeelcdfc81AAdw9E
yT/WHv2CphIak4vhZwEoa5Bc7g8x07HR1K5pMrl/9TEXW5nGjKtAt0v/dcPHb36bPZXBPwxYj6io
Ue8szqRR7uYX6co+qm/bKvJgLNYmNmAsM0aV4ivLp+Qczce9PBb3owZobItWoBEQhOmjL99LErGP
d/sxHoSTRhRejpa2LtsDXoWA+7vTeOe0vPR/HQIGa80qT7/sp7vsPoDqiNUtcqJPYzLPJTunzrsG
WIy857x88K1tU6mrzhsGQBvYUG6s+bdljT60El77ef40JnfzQOH1sqU+DB5e2pPSTumQdPiJ7oP9
lVK3+hHb37hfXVPlu3aYLspKa+sQyZa81WUEIyleVRQHufGrdUVSyb2Zlm/W8L+QGhcOlNGgP2KJ
yEYf1qDTmT3cEKNWWspAI4KUznVNK75B4ScZtjl0w5/GVIgdafbHXkunDj6YYQnNJ3slhXDXEE4m
XamSRhKEljb8XXf/SN/4JDLNwShX9eBvEDQcAwfbRSpbnbn731e04edXN0Ay9nyZe314CtekCHSo
W2q96CzePm9bRcRkmHKxud0QEtUtqCCQXqf8WXLfwixhcttHG3CoMRm2cQcVvB8ENi6InbgBfW1F
tFlgfb4P+a2ijWJB48cQgS5xhVRabgHg6D5gjXZGfopWptEM8dsQ6v6/pAa5FowIFjo5eYtfApCW
JtPlK/PHNbdEmQzg1EPCObJWPgGbiP3xJ/EnVpEoopfHd8WWuNnFHzjSh0Z3LCIotpaKwXzY9zS2
iJKCv4Ybm5w0dlQoAIV3WS6WeWkltmJbFByZdB92N2U8kWjzCj1HuY5pSjqPPtam2SS+Om/LBn5t
cOIg5rlLYEQyg8HwbPP8tgJil6bOjRI//VTAwQwldu96Ndr3OsGPOJpmsR7wgqO5s+LogMVGF1va
Qo562S1qHfLW41RU/9/IxO/d2wgWYymrjjPRldEjXz4eZM4763kbQkHSrsclixfuHIF4ieWV24gO
L3jSVsJQ/Y/sQbYbX1LRo5tUTdlItMXo9Mz0hR0DjCh4/7FoIh/LCBnnjMfyf8OuH0FitW9d81CV
rp9fK78FzaKmcY8CVMDgmaqp3xuPoP98D65OvEsgCMFGe902lF8BvQOLQzy+4iwfy0orYs97ZbSd
gPMpINGYuT+4nM2v5Tdm/YljLmH/DHccwtaeErHPoY/skEbcd+Osk8ACLXZJTKvLWan8ONfRTPk1
a7Qlxg8eysKxKXskIBOdZ8QWPHvp7TzLGY2RF+pNbQKpH/d3YdHCnmhJLR/qFxRk7BmI+PF8CM78
TwnrCcIap3ksgOdS8+LDKRzAfChKHa0hSnFZvw6YGExc91NQxmu+oahp95WwxUj9WrADzmC9aip8
keUlEcrBDp58XcEtp0jhtmrpvbuG+pfcmh1QZlNtbk3VR0AFM2TsyHeybSBNSCNe8Dlkq94FjaUQ
wfTBKO2UhavlxZKU6L6e/TJA0H+9Me6jypjpoGcns2hHGwB469rQaUlk4R70zHMDnFrEN0cr2lxF
DaCvuXbbWWbR9rzPz+6BvtRk+p3qrwFgzz+B1Gi5sGIy/AlODb0viM3JDmJQH3E51e7ggZAkFkA6
G6cgcjRYrlhvcJd6bOzy9FNRYWDn4hvyudg6vE0lsnaV+N/RkDv/P/ph4xvSuZomFPMPjXf7b5KL
EqytUy6X5e6dLVAWkmEQxfjgv9JjPcLQ0AkGgtWvz1p92zU4ax5NSg5QDlmFaR1kD4vPYJG/iWmw
PNuRaAhUJJeMUtin40uQVpyZcMaXILapMhQk1LYdvpTiiV781GJYUigZoJ7usQerMPu8rcEOla7K
khpjCFQ9VM5BGHRe3CRzfdxdDtKr1n6iEHjDjaIOlBf59ns8Y+tkhV7JzxW0CpAOOTl6thOVaRmN
wSywrzqQJKm06Kdc7uO11v9eT8qpz0VK7NRJPvq4CyarP4M/Oj6a8Mbz6+BxOHsB351D7AeABwFR
UvnlZk3uG1yFfMvkkeZdX2cg0u29Qyy/Z8d1lvAUXrlNeVnwdJMotKwjUVKlRzWsXCkvbvB/VhrN
M0S9acq18oIaU6fJ36S5LraP31E7Kh04KenY/KtjyOxflPonale/99APmYbAVPQwzJbdvrD9RKWu
VUwvdX/J1c2zj/IZrfpO6nz/oZqoJ5WuUZuka153Coy6TR1ZrYavoFWIQxa0LqahwNKfpVdAZySa
QMO1DM1Gr0/LvX2GmxChjzKLGvNXue+sgIE5sIQLamlR2vUkbDsf8tUwUKPlnemPG5ljSIGRDL72
tAuez7YM4EoszLtQzDId7f3nARbAlCSLpVlKSsNHRA7kEFETqL4Tu2EPmVPqx7Ux7V2bcM0ETPLl
uEnnCYphjutuJ2aw0fiDAxlkptuvi1C99rhGFOftyWLBGJqbCw6JpppplrXvxAq9kGCz4A3NJfid
Wsh47DgfTlUbrWUB2qcO9QseJtGIguJmAiTliBS8RidatV7hOIt7pfAcvJNSIm3pT3bW1a0+vmZq
Y7KjPPp/O00O9LsIjrkTSNkegnnhnnm3nRRYUCyDxKuqksJMrKneMutpi7NEjil+KgF0pg3imOAE
SPCM+5vZmhc0JJ5dehZ9NAndTBJ9nud9Ku9pJ11fS4uBj+x6wKps+tMzHxhGyF/UeSeg3xKDQvv/
UveIn+Qz9rrfrtLJMvMPM7D4R1IkOXwiyNIAg8BjmZT3VYpIL+O/GLa5UX9cg1Nn4sLwx2FwtzLk
FobeHe+MdmkSdV3FqPz2APz8DOqDyKkUfsvLL2PzbkQNueTFRpW72Y/t6PrAZt2+HSxjDFz+CVAl
q8djZMfQpxTho2kuPYhfBFXsqW6fFD07ZD9aELK4rFiWIPAwhENax1XrKnewFr5AXPr/wQntoE+T
/TFvoC8sLYWeDShxPLwX7lhc6j3i9PaM+NFL+7gMJng2908RbxzgJzZXVUOZPP3hjR/ln+j7NwAb
csaJsl3Ii7qZlkGWvdlNhfHunC3BJ/gnlH3N/QLSPJ3D9jYPAh3G3yaOR6psDYSVIfKOrlT2VnBv
XNKuZeDAg0yS6PWI3hEyyf7HzB9az4LoAYUiqj+QMlKdq9/dxgNX0YNRAKacQKzekMWxxLm9WFW4
wHQ6Uy2H/zj886R+6vIFjvPyoWnFlltVXkFV1LaKWEquyZ5EewKuT+gK5GtwODiuUurkkZNP+7Im
DJwkHS4YKHaWCqNpaOwHecAS9rqGrq7rSahWbtFisgsbPUJpcfhBDQdMZHO0KqJEu9BFtpuDUM8h
aM1TlJJHsKDuwY4Q/dZMBY557P1k73DzWjVkS7sU/VayIj22yvff42hNOQdiO/CFgR5FN0F3Mjaa
XZtDnQhPZpUguKOe8Fq4Xj4NCIAXYhPnK7s4NwYihxvsPpubBkC1iBpTg5C5ia2rP01b0uKDrtyK
sN4CKC2O+tKHJYJzmJ9so2mZCj1VDomoTGini319JmLpIU8bg+HaiNoKmc/FkGJ+HSofLvaVJ3Pm
nlA3kxk3l8y+c8+x1P+qTcE+nUgVdUO8isc7NbPp2TokceK5ahwIv5cQb0ezoAax/3GPkJXKVoFj
VIrCq4C+GmOjPPUif4p+kefi9xsyWiMNbqkNXv+5rK2OkGoHcVZdetc8Q/UF4tDStelsoIHblidG
pnN6M2OzcAfHem9I92KiEr+AbnhUYeRhtLv0DNH5r4V6kLRN0wqfJ9Tad3mO1u9Rpe8mhupp6YqT
I6ox+1LNQG66Rgn3NodUDSxh2ZlsRA80xPSux9BAkOR7cL04su3GDbgL3RxgPdVUYvXDay4AI1+r
KUQlmDOWKSKhjV7IhSQyDZ+x+SNh+dEBF3kaxxb9oCSxSzcMM6Ez+QhRUZ/KXsGKUu4iszKlzmsR
ZQxwpnIMX64DUx8qetmyuF3ipRj7pVw/eaRRqoR8nvjoMwGODjlX4qC0MIadkOl6yxbsB6085hcG
glfQ4B5GsF8SeVSuEt36pgcQOIa32uylp6DrQyf1aSb49X4oEnUPZAwZLVNOhCHskPv85tNYsnYY
x4kGo/4Rc3IqMTo3rqGyShVQzbQaUeq0ZphGbx8xkFB6ie+FOrUqF3aWe3Xq4IkGXKDPZzWCX+8d
vDdTBKtJgzVolZ0An4FuKaUMz4xHizCTl08LfKG5AWWIYEG5L0uvYhKg9Qs22JXg05XJN9tx6faT
qfH4TcDxz/Ie3Vdq191OZIg2Y9pK3LeG/NZz4Hcp5pJjuoMRGCgz+YqYoAROlhRYwTLpWUbwGZvT
gx99WIFJ+jdPnQTgZOXtdmjIhpNSbqhBOMlDwKCxLWVaHiH9LV46ntbq8BtQC2XhnDF/3snNCa4f
zirGPBOm29y3lbz36C4DseWSfbBvHVFmc60n7DWHs9nI4eUR+BYH8rYTf1MNKwElm1CsqUq2YcvK
+UH1LSv1LlH8TDvy0xKm0tZVYK5x3uRZuldL/sGCqZFxAq4dv3La6bpts4tmU0nu+WaTws5H8th6
nicyTVemRVehp57tnkBBS9BqmSiyhvooyvRSwvYjmhIhpA2J55u5GqwmLeXqVZRPIAIUhzQ33aU8
/jwX3r1ZVOmAcRytglEV+ix3UQqANaAYqcL9CUkGDtkuM7rj3WBY9DTkbxr6/farj/BKx5D6fmpJ
V+C1Tu+WZU8nQ2Ejb4zGyvcD6dLmRRC6JYHs1vpVfTSUNH0Y8x74AjrTtDs1umzUL+C/sfo9IlCy
ZIUVwfackRSimf2csfSK70/q8nQqhUBsvCLRVz3w7Bx2Xneev39/WhJzqQH4xRDysHB1QJ2/ilSC
ucuJf9/ar630QMJfF/uPAowbGOl/QFAtO/VQX+vworVmVeYTo8ONO6s4nGukkrQmlMbrG30com7E
HiAIubznsYvfDqkQSg8Q6huSd7HsXPvbOCdJHzQ1h8YyWt5r2/dvqtOQkHHBWcGffVPltFfTf8tL
2nSS8pZhY23Rhwe4NmjaZmDDaa1QECvuFtPNa3R/T0lqg6sRZi5z2tmiWNvH4XAaitC4WZ0a2iMw
MtZ5QDaN5IMRYmptf4mkIvsjYxFAD3JbVfme1ivilkHENIfpHPM2lDsdiLqKCf+MFAAW43ewu2TX
atfTIGIYmIm9HMtvwuTTH33coCtRU0Z6hfG7eEnIU1vU+v8w8OaEDJ4XT207EdcquNlbTr+DzJx8
TVd+avS1qEETojFy66J8yDljD19z8QXwyfpS9FBaHU9zbMQVxkqd6on1F6w3eSgHEgGEVyIVyagC
FwyzOStKGcIsgF0zxQn/4hsnEF+XRn7bNEgRBwZikiRcc6KOssuLUdZuv6RTgIqKbUZ440UsoIer
5twfsHJ+OVxZ8w5PbrKgqkM5HqbZkh+XdB6b1sJQyFurn9X3LftRxsq3qVvLiJbH6L+bH34V0FzS
PoCmYE7vdDRvbOJGytbzKeMJpK3lsjYfQ9DPfxfakUiJKltZ21+wQMMurS6Sfkvc5NPFlbN2KuB8
gw1mbrG2bEai9i6RgpCz7897uMNiwL4pv0RrDicKaG1TAgPPgugAsU8vUmGLkMYJ2h2oq8eQGztC
wybmYwcDOjc70I7TRPda36mOZaVpT5Ry2TfoIeYbLl9zMCpFr6ro2whLfB/ivJJntSlD1b6WTwSY
KmLUTGrI1PShyodGvtM1roiF6AWsdw416vRDkmCAitl6LJ8P6tMGuk484IL6vqLDf1hnzVds4Swh
9bWukUqGy3juOzk+ynkPUdFVLFeMtAN3esAUgihd59m7o96r8Gmad/Ep1ZFlm/Krt3PXi9RtO/+t
rVDJAO5G6kLeLclpO2uRrPrJkPQ3BhySS0ENnZLPv4f60ZHNit/343PzKRH/jT2/FmA6nEu3fgUv
I7SFn1lqBc+KlOB3xphCITy2fanYi65XohP3aQlBp+aKdRd7grhLKgqDuH4utZTYjBecgAqKNGgH
5PcTooa5wPsuG79ORNBA47B+n9fijhZxLLbPq2V8DSZ8o4jHBbhNLC3XTfdJbjTNLcm3kLmDrZiE
iBE0fnRtD49AtAhcgMJkEtIs0xxllcN5T9Hd6r8VS76h8tj65Cb+7bjO7/0/2yiWgUNdyZYknqQf
J56pIPspfpUPHdMuW2aPhJeExb+bJjsgNXqqnF4H06ou3f7kx7rL6nEl5VcZg0lsRAkOKLDnhbzm
koL5qG69hA+nbn8WQqgRXgZ142dVgYXmLL7Ow1sScWbQGA9Le5QJjvcbtIOB49aWB+kEhgy5B2hK
HH+LTzIg5FR4V6qPsS+fZSZtdGysJVGzvjMMMQingAESJsQtIORc2oiUQgjqhKl0CWGMoFEDsqLa
utnDLLOASCAlDDnTAR+FmlIOyO9qHLeLNqbv4h9qXA4cW+jYns4J3T7zgwysFi/KsFZG2J+h6va+
OFA66c2uNZJQj6yGsvMV12382JFZahkb2h0pHcEoxe2YvszlfUlY6xpauuY+PLCIvjhjGtFfh16m
3ZYfxL8QNZHSNuFCYIFV03tulZIBGIuzt6BsZ8rUY7do1PutX4IdAZRW4Cn6wOP3JgZaeUr50sPx
KSW/5UcTJaWJO4l9nCjyeIH9ZYrra+8/RJ4Opt+Tk0v32F0S3pQxVXpbZDKCC674t8F+qQMJ77iS
AU964WrwkP+FIWIQXgvxmBp5+RDWA4QvjruLzVQfu02LRJOrdhzt2BZiGtxoOjN+jT+SnHG3XMCN
zIubnJJUv6xEAd+3RX7ZnzIkZDOCiBVXf2lKiuvRSIUt36CaA2sJ4Offz/1MubSps9TdZUTJ6m9k
+ZvbOQec4R7aw8BDzsYTAs+igfDNPRWYaZ6j2sMXNeIHxP+Bfmre+HYkSiZdIW4My+3/ny2AjPC3
MABll67WUnXpVxgqIfIILgXn82HoRlPajVzrfso5KPbH9yPW3mp5+MDghIslAFCRDw0rllhwZ7C+
AqqgmaB+ioedku/y19ul5v7BDFXZomnNKTs46YC+dVYG1J2S1kr4bpCZ6keTkqdlZAm/ZAPKrHii
N7DyiiPbUC1E1bcRpxB7xiaDmt/+ENGnWmjMDQpIpy8vCbp7LJF8LamsOwVygSKg/BL1sou1CtHa
PbtxYc1mjVK5h3WwhhwGKEh4/orOm4FBYAiNBEi5L5XlOeFEApoA5gxLpbhR0cdwkzGNPukeDbDa
yLrAY+mwvzofeJton5c0t8o0vQQKrWMML7OmP8/osHZldSPxdDDPi+LDW7qVEG6c9bnR8cfptH1P
6z1eHuqIzUOZTF90BMSq1r3CzMyrFXa0zurLoA8kXz2Q6eRTSryfKM24ThnA8oGqwBvfvbO+cNa8
bXvHxd6C1lo0atGic2+WE9M2TB6BSqtNBSMlHKQ12B25f6UIL4KCIRsKYWGytHkbaOrx1Lcgqp67
fjXVSNrh1p00XG4Oua8l4kfxFq4gVrNVXaOR4oz2Ui808i/BcSOK3zZzDi1FgXJdrhC9fHBEwo7W
UlKZlqPnVHn8afGAZRlTIrHBkrGC8U3bi9l3eLqvBBgQtEZ/s7sB6JQ/6gS6JwnakhlTCpoV/eL/
fACljYo3FVq65PEeoeFlDMeYJzDew+Uqg7xZvefeXgXJxA1aTVFCZKlveeKPEnDqIapqH0hn6lEg
oDI7DcHiXjp/VDrxg5sFCfz56JxuZff7z3moFt3p78kztDqh2s9H1jNX13MWLsUNJ+ZIf6EzhNOn
ULy0zo+IZCiZRGfCi2ukfQRXJVKhSRKSYr47jE7AjK8++KNqavAxdhPIHCBC2mWyZkyUtYablQ3K
mYrKg3uViozRKSyH/3q4KgZ/mHKZ23ooh7TLalUscj6GSiQZoncEPEiQvoAVgvuq0RVyklSRTxZV
WiQuiXrf9g1PwoW9tIXzcDFsMs7yLxF7hlaauylDtJlJ7PugTqVXNuum2Vg9t5S/uA1IflcQvIea
MSQmvVEDEMIxbv0y3icNVSoP4Lx7nCdSKyrDJmb6xZheU+Vi20PepNjtTOojwsTKQJY2KoI8fg84
BodaX7w67aEg5upaFK4lyfdsoNUU2ipdIKlMlHmTCy9YpaGL0ntoLa3waRrfHF7OWYmEuicyqC46
XDGaYHjpeIb0njoiH5q4SNA+rpdiGOzPqXzRPYhHUBH00Avvg4/asJi/mPC2FZcTReCkcCFE8bzL
72CxZ/IojtE9kWbWvoslxwBcpyptedjqUr+xcdocH/XYzzeSiTESgB3S/k9VMc2Y5na2IiZnVZ8X
myqMabm5gapANMWAVdcAW5YxJYrngs5vOnU4v2Hzhp1mhRp5kWaKSsAqkZ4Aj6kzElmqJ5vHiues
hBbHwbO9GDEIt4IOPMd7qcUijjQkX7QPw19/jP19ZwUoH7deu8q0VUVArpd0Xu59ziyAj6+80pXb
mxqn7uGJHmYFeu3521Z/s7kRVfhTpGTdLBh9eLXR2y3d/YLEHeMFn6qj4lbpj/apGbfeTNRxR14L
3HoYlzXluuYWnfwex9Cb7/qHtifcSgVEmr0SwEBiR+1qPW0Z+796FcBtv96rNePGLd+veshL89uI
Yt32Ja5HYG9nyXPh1dR/ouScqZVUKosJLelNNP7jSuPJtQt9uLEs/i/upVDbc0CsD10A0mY9A5Pi
I0QEVGEEHfS0ADPw7Gu0ab5aJKmg9oRFODV7yfPaT9p4SGE2TGWPagL++c7ms6uBpt4LxoS+cCNA
3ctB3vWkk/iBp9EICf8KIhesp6lz0UExIeu9qI4yrMgI+WOKeJrr+4ox2toup5MJuJch/cKsL50r
qXK/b8XCQ9mDzgIdMQmYzy+aKM8emSrd6gEqWWxyw+uCaV4bkCJ9Hsac9GHwFp6LJu7aEQ/K1/A1
uk2joPn7UVE/3DFVRyQI6I4kdBlJiOgxuYRgmm3CAMjtjHpFN/giUGY0L6jBvWCeyR+KYvxfkqrw
nqzW1FGI+zokdupucRDdHLXZnxjcc9xgBa6a7/x8b2IUAy7NFb8YPXMCkIICJRxlyuZrRzSXEwyY
xYUJeFY1oo+P9O+mCy9maqJOCoJd2eV2+ksWindVXhrCl3A1loSTNqj5LAfwmO96CIj5RBYwrUns
O7JkyvHu0NCgfbWqwee+VA+RExaTgjRsBgzOmWiAfWnM8Hy9WWHSR70RCiDLbG01KXMQwm/Zalud
sFIag9ay3+WkX4ShKtuWHxO1NkYtI7tviOdDeUuCF/IygsAO1w9zvOaDBkJnu2yRS1A5yv+rwFxf
Tdw3lHQjUUWL0VxbOw0pTdX3+8RFwk/T0vrhluQtvhIha3LElMLo5Q/Xq3qp/DPpcBzBACn1dCI0
keY0nTQhELu+uwGfOa7Emr4DJJDsyjkL65J75LBus/bgsC3UUCMyhQjq8avs0Tv/Ltfkyzt+y5q8
QSOBRRenIMe2sOwWHG4h1ZcUFFNWdRy/7F16AGgHrDkL8y0l9IovDBYhhU1pWU4ywLfuPIiheAnt
Jl+/Rc7ZwE7HgWTxzLBwfEMbdNshIx/jzcYCwkZXUPiuF5F2UbEXCKjdqPxW17qyqVzyRuXssG3O
D3bzM96GvcCknGFTzBMGGAiYWSubB4KYONP+Hey3d1pk3rxRgg/f33oChILODi7EWYZEa837I8fE
lsprPDgO6XHiDcUlflu5diepB4cTT9wetT2nfdQbLIXhOktdMIEUwPQAlRn87FteM62IJc97CbYL
IzxW5n3KOXoldKRW0y/C8aoDL1P/urBzrZ3r48mFHgTOH5pJOJuymhw/1TpNCJw6GMJmuv3kT+qU
dxbsu98y4kQ6dCe501eggFOQL3najBDDIstW1+f9PZ69uZza4Lz1AhW4HgUDE2PNZuWdSzZrZAuw
Iw5rNqsFHh0vwYytS4Ts0YT+rJNz4PBqoVZssYcn1LHT/Hf4skCwPT2HMXzjFeZKhq7tIoQQG1JK
/xNGl0UmmvyJ81ye0Twxodr8GbVkaHKjEomZfR/gg0AromHt1pN3VrSkRZ/K1C5BMrbGfTerSaX4
0tpkZffYjhJjRJTvphBtdnGHYM1gT34bObL9u9VPHvpay+uK+hs5gvgVCj2EjTuD7L+ErKnqBAG+
93dxbRrT524qYIUhh50qXKxqW5pSb9mfzla/+9zG5hvaZkcrkV1J6g+IrYsAYKcYCKEAnCqfWd69
o+wBvgwCWotHItYhYMrOrF20EyPTQqPc1dJ7QP0MwNUpx5T9wIFyUEMgEcP48R711GdKQV/w2Tnw
gjOE4EScfwz10LUBLdFdZYVimHgxB9cn3xHFMwpA9iKiKqNy43MM0L17PDiJn8T6oEC0T7AAuZfa
rDGYDEgHY4WjGxk3w2o8WvorYQnfUnvRM1XywGpV0fTBBEVPp9pqT5KTZ6Yj2Zj/jxepMKSwQJNr
ivCpniumTJ+2s5l8iGRzvJeqGs4MYMGh4kOEtjtYUd13dLjDnSLwFEpgXOF8+imN5YELL0FBGgpf
mUQw0T+XqOjX8Hcf4DQ0+0TgOjLdxmQ51aKXJnkFNb5Kys0qxzwGSGKOSijKEx1kWXxo610RrTYO
mvkmeuhartHxjp2Xj8xs9AgFxHatgbNylOOq0IzgvfSJhvqkw+/XAuX/zvshyTAREljMZchLUPhR
7uwV5W4XEfJiEf3OdhXw4t8bHPr9CRcmYqAiHDrsE8Wljh0yWqBTCO6kqN+2zqAJB8xoeRBvTD5g
xsgNCWLBnCHKVSc5naD/HBz7g+ciCksa4P5SVl2/ndwmDE3yyc4ITP/K0ZsDEph++9flo6wD8OFq
ilPLGOoNuvci3H6ylCjhT8neTi/LDAz9iDZpXzD2CbOsmGPR8ptXeL7aSBL8yH6YCXSzm7O0IzFZ
Jtgk8t0a6GY81UaRT16Kif8VA34kgFul6goddd0PKRUjUUs4/Hd7dHi2+BWbVtz3eqwpRadupAoO
bwq1cowqDYylE1EaWpY9uJtYWAv7uFBNaraKzkb2s5KN9fPuA4yMyjKGQ/hpOzKUqmbB7GysJFyK
Z8/CQn0outGAivYDgE9kj6sO5GvSZjPUyinuE7RmIyINteyFcBQxeUda2BsfL3ITr7tBupq48raX
pZ9vD067egyb6Lyj/rmiPLPBQo5LLhH6DyKEYTDHNCiVtkKytd5HVcKDniQXsH6xkp6PmIdoioTs
absD3tcGBpohe//8ypV+vKJeDdDN5COS0yaiMBUVrZkG97HRBsCsM5NMIJyzw7LBNuUcMzwjGCFs
faWhJKyIuh0Kj0GMwglcJZtuQT7EJSbOXMcoJbKwSARmGTzamvo1jgrBjO5OUq9hLGbc1uMlCkAH
zB0e0Cj8vfeaIO31ADg/gjS0KSRZiX18qfwaayx/zqsGx8BpxJ2aRZuCooNkSll/+sxeSZNDtuuR
X6LP5AJ+qo0FCoVtQ5xAY/pb0W2Bcy0v2ELcgQoIqhCNgvix2D9mKYli1mbq9Lwr8ebeGlZ6nuFV
a4Kms/Il6i16v6G9RQ+3Cmgbjhqk+K7iUeQZhjsjDfocyy2zwHW3nsTHBaWY6n7UbeGxe8kP3h2w
OqCUPjWGOioHhM6gzH8SflFJRhHcNXMF5T7CHNt8khrdulflt9g7x3vqoUtJC8lylsXWOsrZ15j0
dupIP+8IyybF90f29vT3CgcG7CwyIdw/TNjeRQmdWPP7ARBcA3QA6/BPJJL00AhOCxpwZ4QJCIcJ
NYBcbHLMLqo0rlkMVKGFdIIYQ7EE9mYoc4NjVQJnsAToQeofkYrLBX2nCs7lT1AMpRXFBcSecZDN
6UM9hJ1k9RR+iQp2jZHiTgkglu+t7EVhnmtOi9JANHfmssfX1mnGJmofEb+ZuD1mSbFfi6lDuG0K
UoKHpyONyUdqT+iPwO/lUUuc3PTJNtb9PGHasmfnQo7Tp3FizmEhzmfrHNERrKUrYR/5jZYBq341
28h6m0PaXlO+i2l6ANlf9tjE8+DmGQY+AsC199PcrgL+kllmym+OR/FvWTMEjscfqGuzttZk7j6b
u/19RZ7aW80YApP2U/OdgSCFYUqoZRcfQltuD2KpsIHRREJkF1NEjnVkfSvLb7fXQ5evNlKtkwAl
YOfxhnrfosjzhGSM3QTfGNu/3xobWvUQToyTix/Q4s7gx36uiH/tyfaYqxvP12JNuvC5ouYyAW5Q
fkVyPFNyFzQiEl8hBFWs72uHspAR/F0yos2sbXkquw6k4fJ95WFA9RYSDOQedPf09vO/wE/nvKBA
GeC9mMxpKc8UarN03K9x24fAFEAIqeMWkR88QKOpzwyhUOXtPg+9UEiOGIZmjA+9p9bVOZHylQ2q
SFd0KUS33PLdO4/GAUGmMS/sXQluw1TdvTf1DTEHKvfB0C4YkfL+OvnLn4yMpiectJJUXsY5PXrx
qWhsSUnYJbHWKDAK+xpyJHPCHSrHQ89WVtp4ch7JzgF5MhS38aZHtGEJAF5i0HExadAi7y05W9Hq
QSPAAwlpNTxLSlZ4T3g9I4ZYrXqah1qk8Z9+40PA1L+OiA+KH5h3bTh58uoqIOrMC/+3wb+HFkJ3
MbdtetRpVMxYm63ZB4U3xrrOwKgbLFZQYG5qvW3AAKUsDE7+kxc3eZVrvIK37YR/cwq4X0iun7eY
GNSVkZwbGitamOZ6qcXx54WbYN8AeXHzQTSIEIEvbtTLUMsuYyhkF9zvWnnE8sLMAZgH/awC3L5G
wjSD5ST3XjOlcs2OsKTQSpiSM6hIRLhQjTT0fSuvWtZiOoRYG+JE9DQb66j6ArVwPZYp/oZlE2uV
d2lZ5xoKa6mdbL3EJOzMCFIk54XKfyJHBUl22HOLksR6378nPgHb3+XU9ujhIyqsevDrvvQ/QBxH
zbqp7GkszeClTnFXtaIZkdF4LOgV6DSaBlg2IipYR7cosv98dYLpgIdF8wW51Sg6b0PowuCKHLHC
y3o/WTwS6Au/srZNHrHa6lZQTU/Drl5O3930r+G39eBSJhGjzmiWtkUgjabYn9+S+trtULbDdUqd
zG5tYtDGhZ5yAsoR7RzizVUyEtEgcVRYMEVp5d8R0UYefIejUaHe+x/sigPkpVfPOg98HNaLe5Un
qKRvialYlm741Gamr4BTRlChJibz/4XkKfLSNLPx2vmbycTMEGZ7F/CcLm1pSsEgDDOfPrCrzNT/
l25ZBkpcf++44put8fYkuY/JZOeQDI2zQF+CBUO5DXudbhBw+Mxz4tKAVaIuex8RnnDq91LjSt4f
osfbjNksTND8wToJis+/l1AlVAHtvP+pobQkgdgDC0JEM0zxamJH7nCKe5jnpsicKtzPU6bHV4L+
co0/I/gd/tg4YJY1Jdx+wDKN7p8KJkkjmKGjbPlCDfR5IqTAq15g9IZo3k01ZZfTCoSu3c0jNF03
iL6oHz6rPslm9QMTHYRsoxD5tH41PAV/RaFUq1kMtrabw/Dn3X/EwI5/HYik8qS0vTeJTBwL6PVQ
i+tBRL2UxXCOq9Hkh8pD47vWt8MaZcYNQbMGNoFqzx/dDfX4OkDFeIgjFVAnxUFhEDuHopfD6mG/
VE3zOtNzd3FpZDkhHJwAWrR5Ycypuz4RTh9SqSO/sWdcLsWXIvXug345sGtK3FaPxazLUL6pwbt+
AoHJfvA1+Hdd0Y8rxSWTm0OuqYMXdT0hEIzL/O4iu6Qxq9tKoqqd8s1H6/fyiZXVlxRRGHI2OvzB
8AyHQcCWBGI7A72bPtFlv51ToR/0HDWyHBsmPzHGo+M+c7mglkvbJo5xzw7P/X/cKuqwTcpXM+QZ
LQSW63W+9J62/83oX/mGUu6hSru3xVDw4a48/Xogms193X3MGXEW9LX21MIvIDrU3EnDDkTHDEWp
S2PM9JhJYkAImPZ4Kkje/yZ1Ulu1sKhT9n8RCSp/j3zlgG1WURIaeiKw0QRchGP8wqKikzhI6RMU
PztPRuu7CSYpoR1+Emiw8Zt49VypXmhD5P2SY+EhOidlg4h0aDA0foyepdnaelrF7MlZVbAwSnRY
QQ8fSsVx8oLA9BQ4fJhEDlJJLK72iTLfLqOnGgNRiStSHVFTBwVaSldWxcaHoM2OP8elV/ygFHPM
HMhndPx9RGsKPA2lEakDBQN4YxDpWxukEi7xbVjf45Os9oHBksuCWS1+1mUWIZq1EQsOpGaxVs8K
UPjP8S/yUYZrtnlNUjUE+HpaH9sMrPImoexg8vvHvuh3HLKSVlfhFuKXKpAA3mpHZ6qkgbFLl/1k
MxATe+HWqzo4FCpnIJuAKsIO1tqbXWD0qhMyIB5P68vtZzwAUIAPqChiMNoVjZuaA/LE4Mh5isJu
4/WcZweBtsiGMptKXmlovR35rihaqisihdhaoponm3iNbnfXWaRc3lDryAKggnCbiy30TUVce+gK
e4R6Vmfmjon/HGRAHwuyu/IBgSLx5ULYAlRpt1RXsTNXCihrl3KSwdcf6rejOR8SUZTrvMCR/KY+
CAEWPJA+JN4YLZgQrnbzDfXv0e/RC938DQkiiSa7x4SnpiflE3ClOtptICDo87LjDoNA+fhTrT06
o7ytTJaJbUgIAzRqJ8Y4vjxsIw9XRNpX/oaVU4GBGXgAnK+WgQZvhKhGmujuEixmQSVvIA63cmcp
vgNN4GeiuPeWB2A/duzvDSSeyVi4btN5WMEBopQ3Q+8G6D2tPI7wLqGgE7cy8WpdWTx3D/CtBinY
SWHqZaINELFc/5YFRoZHC0aQOfJewUdBb4Q3HfbtFgIryl0HhMH5erDRrH5bbQrYLp2oWKRiUE4a
fXT9xFLXmBajdMWMxJDMy8ohWhn8vFSXMd0XJe+MoIjTxJidbtjpypl4wJir4TwLZGIZdGpQvEJj
2Ol95/O2MU1y5UARnAMRtrL7/tpqxfn+6MfgbEF7fatErA2jp8X/gYlNPZbQD5H657Kq21yGbdeR
gGtxW5qi/SF0WgWSmGmCvbuIyU2Fw8xwQcSUAyHLVkJAixybdHGbDN2pQHLc3dBCwpVQrpImdoE9
3TvCaRiFGxgHlz/GvSt1QuAYfbX4NmYL21bM/i6Fs6u/hZMJ7HsD4XyO+5/wN3ACCcsIE+zn0Dea
Trit32pbYiCtUrXbmG7lxCDFWXIRo6JnilRMlJKq6uwCA7gsbrXkeilqwXtHp8sdmQWF31bFvfwf
LysXQi7iWrnBy+eVJRSfo8LcM1Y09S8meQtqlKzOrdLY+HtGecMbat1ViK4CY9BhlgRP0XMGn4tr
aRd6TNLOL66YPUafwLvPsZiWsCMav5IwYSagvgplBd0q312r1u0G/XNoFrLrPhQBCBIIrwGVuEc8
6nCpDRx1ToOrGHBn7gPNHpKp65LtTu9xjQTLhjafDiwANdX6aPX94BL7Nw1idvIa5d5yA1ohgb0p
oqaNW/fN6dC8RV1XPOw5R0fIdOU3EtnSfsGHN7K1T0ibdUdqZI/uJAgUodrfb0y+3DxLW5P/n23r
KbJMeQ9eH+GavWOYWuFXrPT0zkk/nNZwpo1lB8+TCtX8rq44zlTE0vUy4FB1ILs4iPedgq91Uyl9
11HTN0spkiY5687LIP+hgY6yA7HGkPgn9ERjCeyIDkeksiaTXoE+sOgT6LLf6oU0Z0tQs18V3wDt
2XNHuE26km7cxii+gPiCd9+wtb8TAd0vvmq3dh1UJNqwzBVEU3/hQZnBk22tQsul4JUeRLpLePcz
JBh/w6K+MT0m+ltslNXwfrZcq+tXHM+8/6qsj0+SwFMOojGPfriBgAih3HNvBh8ewv/OXClBlk1Z
/C6F5ZtTQpEhuWxFT5fLtyZyRaF0FFVqyLqjQrBIlxh7815m+qf9Qs1TvhpL1tHJ1G4cQ4Ce0s6J
7LMXcrpxlkQlLeQvAhdjIrVCELSjB/M26k1KAwbpzz0uS3yegN8b+nRn/CcCGZ4bHFc6uLoRHWpl
pUyUMqBRRLg8aIZftAUQq2nF50vXJQQ9bM0amz1kkVBefGjNsKMWPCYayDfAYxZjGV7HGSSbPrwl
rK6ZiiLVP1+FD4Na22K9QxOGntasmDC8Vq/vUwMEpVleco86Ese8W3l7sesJlA20xT+Lqxb0RFXl
/6m6U2QeDcD4/5bYPIOZ9+pxZc0WwtuZHMJCRz6Ge+Pneo88jgSahIGm+j9fhxJ0sH3N4i6xQVdA
WgcFPmgWAT1t1ilAdz1HtX1JToudvzt9p8KkxnGSEmhf3mf2XteNsERgZ5dTXuGCmY9CptnuqKAk
LwuM0t5aZ+yJBb45tw3bZDvWxGZdjKhOYiNETz4R9sIaokMfogYviyKPtG+Uzj9cQ9/Y0YQL9fGH
zgbAk+/Bn810uLT5DmRgf3H6Uf5VVTPo449qAJpf3qfy+EsTBfydk02xbngOHVhhzCBQ5ZNzATr8
8z8KiiBiaIZuD9riE54HfVeMWaaEUGG9wdVRRlLLhGZF+dFhJPvxKhQ45jPo8f+lLl2PaT0h3MV8
6uJnxa1jgjKKtzry56vtgrlMMe3Jyf401dn/BHx6sh/dx+W3ZGLjlFnr3b7gf1tSc9ZXZhy/k2SF
rUx/bpJzgI4Q+YhjHVicEV2eWE9AXL2B52Kra9riVPu3ULJHkY5smcTlr7x7aYEC78fRtDKz01+M
NOpO0rAzgl/6k+1HM6/sDyVGxHe6l98FXhDt+Vm0Ln8ta/8N+bzs5CQpdgGL/S156VlSYb69S84N
J3egN98kmhUeBFCYo/o1tJrGKivImv+si5Vvejh9FnJ2bCJ7c/11IuudI5fwTLpzvJCiBKfB9dNs
LzW71RfG5cvW0K/3lt3LKiWVbGzKsBbh7Y6vxn0OUnaw2wIBMMC79xMtX7/ISXXRvMsO5r5nDpmo
A+/aSIfR9cVpnt6ZmXLotfPes+P8DP0PeYYQ45nlJilBRuZaNbW0hc/ODct5wOykgg+8h+0owMj0
K0cv/S1auhelg3+kuf7or8WcsSpQ+RAuyjpsoh2ING3ohiAAognOE5MikTTUMHbG5N3PTGd3ASSC
ub74+QzchNSGGpM3KjP8JoK5KAhu7AZffyDODawzeYWTWtUuVTYA/xsbfU0IbANzPpCF+omt/8pj
mZKYR27Jk7WMzupKsXutpWTOk7yEeS7p+QftpHmSo1vSypJIO1v3JdWFVB/NdM1ythBKNIr40yT0
zQIjZi7bvuxXKANyP7Af2+0zFLOd/EUzqPcOOLq4Wkod5UlVOqkZncyvtmLlNOpyadJx1tVuzNld
Xsg6Z3a+EVp8u+o5MLQxPsMsfeA1ur8adn1v7F5MS5gcgsozW5gMWBMDXNIqjVS4IsetYLtaiqLz
SAYgOf5cMPCaL/DhXQY0Pu45CZW4aLSbbpwSWSPbYaDmOGbw1PYWla9dYZVLOWcyr/WK7QQBst8z
DXICo5RuE6LWHRBkEbi5kIUm8waU9B/qc1wZvNk0rHegTLvqp6ApkQRirn6BkFovnCig6WyTxeMQ
PTTXMvzxhaUxUcrsrFA49WnMLPrCOgTmoNCrY2KLvilHZeJ96vzsLWga1HZXtJoUl6EASg69hCSG
UU0oDwmTZZiMsumgch6DUtwiCHdTWAUXiKCen6AW7MXXmREkzRHm8VFxy9LDEhoxAghDF2jJA2fX
P3bBhvv+mqrt3HfenbIUrQyzSv7pyZykwy1tlQTiSD5MO/DE2fPagg9FP93Wxp6hJHZP3Vz/hkpT
eM9zTfUzYAg28DqcqlwjOzdSCcgsZMDKLubipVEk7g1xfsXUhIwxS1rB6y4rQOtJOPLhAsKRuvkG
MqOIIaoJZLpZ2FDIYz10qX3X+deEz0w1g/mzsu65e7Ipg0JX2gfPW5SeVEEFOqr8KYvj0RmTYxIh
2N/Dl35MTAxHvvXEm5vD0itfYQojFV1HaOv4mqvEGp/Oj0NkYU95T68FMLbJFZgeDJyHKdLniig1
DIMV8bFyKYC5p/MKar6Otg0hQ246kdrxOUCskGzzSdDBzhFAL/QArZ+t2f4HbipchMnfTyR+KEvC
ZLXDSIh2ESCczCWp65/g3/S1sz0rmLFYuHYfZyB+AFgXzle4kDlNAwOmgxSx9e8G3PE8tLYdwG+y
xSZcMErv4aN13dt2yFar1p23V+ixY4EGV58mFCAu5o81ZzjXNj6s55K2AJb4NUmgAongW0zSuZHw
DPYfPq2ijo70L97/5dnvTUR5/lJSjTWFoq8NCd8ccNPOXzjXC9L7KaFBqnJKMSqNY0/yInXnENzY
P8LM1s13MQ5JI21LVoMFuhzWpyk/MGMxreFvY99I5yFDlAna5gyJEv6/PoRLoPDPHS/WA+HokStH
VxikW9mPu1lALoP+TMQTCK5zfWNdtiqhEpwcrskWuy+KaQ8qMo/tU5LMB1SJEQHAny7Xw7ajqR7I
0fzZUFSuPyVBzd/54Q29wBXARfGP1Vz91d2MHod3UdH3/D7V9AyBfEQCWva19BME9JXMJzVeWxA5
keX9Lpg/Fxt+3+Kbqr6PcPPlNuHTlTmOPzOwffpEfjpFbWUy4DyEhuCfBhDkRRgryt2c++Ku5axX
vyzBSwPOIYDhmAe2nqf00rkeRgWqESMwRc7uNUS4KTvuvDiribsbq3I0zqfQ+Cc9vJkcsCjAMt3x
KGosq7LJHqeT05Degr+KDpDX+6jQ7aWr9CHiGlMAFV//kDKd2OQ6CsHRwzlZ4X/lcEOXAiJ1ECj/
i5aopeqiwz1l4hziCbhdaM0BUvlccSPTSzZ0ZChaMSuFFGeW4AoQaoLV4IvdmIq1tmpwVxyMscFZ
iHa+9J5Jradfivz1oVE30/Sr+IKpbThyBS3TjKC3UA19vfqnCtMfJ1X32yTRNW0M15vcyI+VJpAf
NG2tkagYoULDZesp48HngyVL2mnbQJ82SUi+pUfTwmichmDyxBFhVAVdTtas6PDC9Js0JfmC/Sxe
Z2AXn7rRQ/tIqYV/q/3i/huQDYlc04YVndIWCBhtnGjWdnwAuU7jHUpBo2JHZseiV4fDYUKi+9v6
itbVsychzhQEha6a1LuhFscc8l8WFhG7oVsO+1f7gfoODUGSnka0AvpRdk5y8qMf2svMvTw+tqLI
oVze5wImsYfFF8SknP4s40kcXw9x2YYwn0m3obczjc1OoLblFJouD+Prlhh/UDtJQaBpihnYpid/
Q/Pa71BC358tRJoCeLkZbgMj+UhQLMjZZZm1zQdA0HJxDlChCPdGnk9cPCtMd8vNcDEPwVaSOezL
7h781vwkSsSteGkl9MAksAE2o8VycybNmCMlEc4bZ92HRVW2Gy8hvXOme/zFFWw/wUCjFfA3s2PU
i2s9mHm4Z9suqyM/dahByXm0/FhV5nGo5pJMryywSVGd7c0vma04d40+agLlNONUM88i+vnCvP4T
O9f13R70HjKFKpiNJZT3lRUcYT/dKgTpZssol2L0NEO8S1dVk/l7mFkLR9HzzQSPEa+ZZXayvlOH
WO2C4xHB0NnhVURzX/Wi0oomCkLNp7icpHinRo/IwHsULrRRCS74WxQ59V1gtP2EmLZtt7tr007l
pLDlfJ0Z9axCaxlS54nG2JkM1g8KKer1znbZLSbI061BcgvjbCtGqPcoCq2wVaI93o6LxhnKqNDc
vY1rkaaKVPk2UX7hcsgITplwu8PjzmiZY7xHT9XgcpBQnNE+comF/H0ocLIg4fgVeypoJoblfEVJ
MPwgXu9qA1g5pdkTR8x6o9TGaujRZh9RlMGmBCgkQckU4/Z4h2Y4tjO+qfWK1KtImK70Ze9tR4hf
+SBcp5nI7I+jo+bHgTNmNKRuKXmJAxmwZiE4u2wV3lMARHIOF+WIqL7oA1e+sRO9wfC+HyIuoGnc
QGekvgOgi9d4ae6tK5AhSb+ZTQJfR6Rp6Qc5kErVL9QdiGd86gMYrS0juRjEbbvpk/3657br+OJK
BNtOtrksODpfHH2RT//Rc1ccrghB5M9vrkqVYSvNq52BRD36QYo34O6bKEqqUcr0UHAMfrPlpw7v
/wPbxwnE9STlQAeZFroqd7uyFJKzAI4k9EFONROhUoOQcEAd1tOHQ+9oAwieIcdDCvHYE510ZzBh
ciEwxkBhrUeduH/p/w3DMW2wqmhgpEPcIv5nlHYchn7MMh4DcnCtermg70QglXmAp4Of56jJztMJ
iqFXqyN2NKqvQNqq1nXHuapvyad2Pgc9cT9VmXnKHtJrtb4ylgAGza1BsyM1qVHro8DuK7NsPsmc
2033F14Hkgtq3UVaG6GLYDwZyzctoG4YYWbLNwu5tTm1smjrx2a4lJfAexhoPqj/Xd7DvFNGZymC
uR4EJVvRNxB7jk4ZZQ4VQ7NGDNnX9fTN/amiPlF+Pr9/FNSOfHLRHdqbKPwVdKiWk+BAejtr/Rfi
r1ntSLqlgYwWCgKLZlZg4R1idQ/HpzacukxRMQ+GYhyVOsVxKbV4CP1tQ4FmGsQT2klCGpyNm/9e
RoIjYTqyBt6LC38zkwSRp0XMiq1ez3+QjUqwrXn2nmXg6l61PQCdPFvbsfBFtGv/Y6FQXqFUIUx/
6um13SRmJ0ljqRauaL+XsD+HWVPVfASwey1jcgCikeZN2oKAzEwt020t5dSH8r0CrchIoxmnmQ3w
OPpd2d99gqIn9hPKlHDvJpmJLO27N01oHjIMC6rppiGQONZb+l8AokIZW52qeVSKy/9ov2n618e5
19x6XpZFxM1NflbOy+aAdOxgvKuLWqqo30gDU/EV921HQDeE5OKi57i+IM5DQwDtK98RNCxqCtJp
93zPOBSXFzcr531WkiFAxO6jrdMzSZLMtGqx8rgZL7eHonloyAcOOPZKzYK47kZhYpFTWFEpNvFv
B+GdeQFKEyuKS+ZdBBdjcsrfKpeBcKvMjZV5WomLEmuBmrkhT7ujJUsgvtsz/opzDnoh/5TLq23T
9yClOXErTcUCTRWY4fjhNbpGhib6pDkClA5dag21WEd8V0615RJ+8nJFsr63bhpaLaj8x5uGxVDD
+7gzQJpL/Rws5/F7WFT2kgeYarKV3nwcFNBtHfg3s4ShQ7pj9TG+YBbVVl2QUVkLmGVnPmbv+2AJ
OGrL9mTd9WbS7M7cLMFKJWyFudVbzFnXnF45EB0zrds06Uof6Lm+L6/9WIhwOISygOQ5vsws4I2K
56GG/zyg291zaEOM66xaBAYnCGkXcjRPu1w6k47bpCqV4Qm5KAW+G5s0ZECKpSQ97IB4swgaFJqo
D75T1Ac3xZS4mMJTcsqXO9+QXP45rNlx1KJj3hB9auGNcgC2fUL6nOl5m2qeR7h8327A37wYGDWR
hjYmVM+ehBOhLKHScOyag9aPh1b5QUXd39uviYI/yddx2mIllV3fl59I+PLbCS5gCR6oFEbwDjD1
GcZqKzoJNGByUzS/fN1qe8UhX8GzrDYD4FtGzik2OtajQGhvM0M9TeF/JpiJtcHd9OksMHSYBAqp
YJRTX/m6BJ6/UH/0BRFJjrHsa8F4GtZpt95B/+ueK/EMzgMeep7tyEHd7rPOtmcbSC/hqJJY+1BB
M4Nseudkr+Ct5sDuinVsCsMz3mtTfg/uuU7xxL0DLsvx9Lm7tIS5BG/sf2RYAmGjD861KwOSIuRn
rAUha2lv5V6PNj3Rmwf854mNc7EiwCu2gt7aHwdtKO0tp1u/yWAduwyKjZxcu/i9ITxnPtcHn82j
SxXlDeW/v7oSgKQCTcXu8FKl5XzjALE/wKUXTOlIrtDbP9Pc4TDCoxsFqmiw/1hwCeYLFHh3FN1b
zGpKkiOZm0tJd8XYaS7l280K3dB1yakU+Mg2VZOj4Ye0PRQkkVqoMLqOHc9GglO3Y8k8Xl3mt4Q4
ULd9f4R6tgH4/0343mwZKtPxWqNjzqGK4MGpEMFmKldBS5JzGYCv9Gx6j1jIOEKMAmfVBw8xMyoP
n95eHpySF2tP6FmSjypGX2I9E0Ayk4ZsdOy9Xvl0mOPt+YCtmLWCyoxq4jGI3yTO9x1SNiQdznMh
BaywpKZxYh190AvVfAP2KjxPjIEit3NZIIPLRIiE+Ph7bttDdNmbaBNc1IqmooOjLWMe9jmsWYCN
x9hA/v+/GFClw+gja1xCmH/ppi0alKMY7oy8a/ZF5FfZSt+8VFk9JMOu6Fi06sEih87uk2SwA72L
49Ja8wDm/Jd24WvIh0G+nVZ6eCjhlvQfxETX7A58d1Wvqvo38UZj9bHJLc+qq4k1We5/09yKVJu1
1uJQLLSM054lLU9/V+7CGIpGIH4pmdNUZylZxxtDxourfe8AqNoQJDlkm6Gw9NhHd8fHVylk2e/d
kzy30Fq2vF8V+ebofDeKGmiTKvfFuh2F/3Y2iJ3rvEotjbJawwhdWKEqQ1JOvqp5qdQxG0+QlIGy
Lf05zdbm/Bo7DQp42uWsWvbOSqnLqG2bjZiQQNPoGTPmKBQD7jkfJsgq8nlb4Symzm/0LQybitd4
94njyUo/oafd+N3J/il7z450CrZBfJZWlwvO6QFfMrPlJWcL8tXBamQp2UtJK4jzXCgU0IHz0Gnk
bZBT7RXd1vnTxDgernunpAQEF8WMaw44qyWV4c21VN0Ixy9WOJr9YrFuLb9VhSq2odEARNuInjQO
vrAv0MmrLYQaO7HrYYD37/ui6jzEFEGNIcg3dp+vHgbTNbvRb0E2RD4tTHXqRUi8F1lsmcq7G/E7
57/94ehOomfZWMBErVEAGQMHN2tGw5idx/XUFWV2+a9tYvfLil4npjdPiang69p/4+SvRY7Bqm7U
Qb3QSfytbKQZffOOBJY28hD23RO6LeuLfCUmMN+bGYypeCSXm+A3IPDZJYbsZRNR9F7p7Jv7Km98
QH+NkeBPr3rHxZAQAiJMXkIP0rw9UKRoXGP0uVdV4FuzxWNlfp3qACM+5njHEVD4oJ9zK8K0y/EC
yDDWbwbkdPrBbBQ2UZOte0z0KFbXuNL/bjyUEuEJXCHQU9kiQhX9B2liUHFNH9sglz2PrB01Yw0j
78uXHiY81Zm0om88NcJXI5k50mVaFCkt/p3mlWbmMz+Bjt3PEpUX/SNwiX1k0mPTKTzUyhW/s/wm
ESRjnBHw4JStSO1Q3A1CCemgYBVj8lXSEMhQ8shN/Ex6bXb3efAmaABqPs0vA1FH/hBC/MdIsIA/
s4MSWb3yIHhLBRAXU0H4G9jve/dxlKv3qNRmvb4DTkGP+DkuXyMvVAKO51LZsS9SmW3DXxEGk5VZ
YnPhdxqclqTEVpZJ9Fw4bao+uN6NHEevCC42RJUgknSZJgSMul4DAl9CT2VWgml1YUfdm4AxMCcs
lPCr09vxp3POJAmM0w37OPjhCf9DOKQxL7RTbfVp7RrtcISPwjCp5f+ZpFaeO+XqU/N/LqyC+pUi
I2aOcW8TuDUOvWgvTl3HligdwpzV2uPvGQX6ujQs8uwCvSdS79VorIte3DnFv6gxrqZSYd9wF4UN
D5uoWWA64w5sFUpH6UMLRFD+wuE3HyG858f1Y7f+62Pg3rSzrFsce5lr0TLEt9zZEuDXl4UhEnBq
mF118e1fTnt5LDGeIqsvZ/BvCztQ22c2vuAR26V6rQtPabFe9bMoP9mKU2O+AoK8J/8lHAuq6UVB
g1YYsAKpQArHTDZ1zOWZkMYL2LL8PfPqQiRiFiN5Fj4Rjt2NWyTB8/9eDFonyKhzv1sSAwumvC0d
VbdFnRWmDMeklVhffRoVHjtmis7FHKOzmvv6A952BNIshNXuGKNjNasjA6IsU/RquE6quVTiDC8M
osn+qHuptRSM4/SzyEJZfAKKX0zGxOcki0Lsoqf7BGmQq4hNZG+BVyN+UJvd8Fr7n4Dr1zuWFaca
IgJYPYJ5i6whaRbgeKCOBvLK4RC9aWLnXZSznbHbuCuEHoS/JSMvcFMU7WtHypuWu6HB1cRp3K95
qZqRuzhAm+I8YeagNa7gH9Ixk9xUdfidzEDcxyqzyaa5ZJE/pVI08+Fap8HsF6PKdTfzY9yKBmzJ
bU4oVumb54QOx/h5Gr5Yx2iYxt4GJB6yr2M6bE8ODz/svsEVhpUz6kinsdLWZHy/D5osJAMKMUfz
YLTP2KDiWYfxEic2fg7/VSaUWxX/cgMKRVTzN5d+cJtwAEx8IyITvCjkL+XUEoCCLoFJ4QvcmxnP
p7hz7VrKqJZS/t3EDpAn+pT5a3tc8XY+ubm/tXqnLKGApfcp3LQxSorJ9hreHZA0NcJv8AYhZWj8
mgwnqy53UZK32R3AC94kJEkTIiZf5Kj4QncvoYfjuwmpRA5Lu1Nd7Wn/X6Pvy3CSNJN2z7Y7Lhm1
faj+ESbsHzgXfpkH5GrT8hcQgY9dRwwkdr9ZqjJRHA5rBG899VRt9p5Dsmi6T/uFEbfPBWBm9VQk
dPSE+t+2R9E0lpR9pTmkWkoQGU70nC7wmkhJvJNPxIROmbPgbx1aTE6hD3B1U8dccCf6OpI/uJTi
nNeF/gZRRyFLAuO0j9KbwU6I5ahPqUkvVcIx2K/PCfqFm0Vf/s5vmnXgijNmhoM5VrnF9TYNsWg4
AAvGisf80wwBLgwj3P6lBjgPO872fZkklh509ba311BHXMVcVovLEbfS3MXfZWVCPE8SyazyVy9Y
jS/xY0u1eVcSPjzXEygmirG5Tn3nVAKuq+PQRvDNYpLPOidYhZ3VvxKEQRGglWzSBdCGlKxpBMFj
BWzRcLQolq3toRGjiO6BWI8+L5F6GhIOOz9hLUtYVOhb0I3ZiCQQF/SkU35LeYPq6k9GJjBS9yTl
O16D8YYeuAgBHXefgEKemJRQ2RJhhHeZ62w+kpqH9sXoELWzKDCcxY6bTAk7gpHBPMYnE2GPTAXA
tmvQvLh7GXePKoYlU13N6f1Wn5xP0HT/iu047p4u1Ltg8BzkfTSK362ln7PEUeKByGmxYYhmJk9y
Q6SHTFX/mTmCpZHNxXhZyLUr/KGLjwKDEIzWgz/I8t8WRlcpwdMlVG3RFvAbPjixKQR1xv8exWR3
h0fvx7fejEhacXQAK/J5Wuuonsn9AvIzT0zzKriYnr7EZLf2smxlwDMIZUHrGYtlpW2GyxYbqw7D
D7nRAyLFqenb3Ffq0DAnr+gTjtknIpTUXww9GhAyhDGsBSFMMAtf92p8CjDuHXJhHotdnWNKwrj2
6l/dQGXbxFPqB+MYe1geKz+FycF5Qc7ywRvledCu4bVGjhN1aVaeMBr/vYG9K4/P7qWdkA7bCf5B
4QkWzCgDBCDXJv6tdl+to4XjI42CkCj6WeEVoi2jNcvS0bTdzgceZzbBFow7bXLwKQAwzNmd9OgI
PQoyWp0XyTKH44KKhHApQ62El5eb3nYVZZK9YFNpwSO/aDvZ5QJU5epo0qcrrYMYx/NGdLLE3w3/
P6WIoV+BIm6HNKt5BwPkrwg0OGbEOYaZ70taJaIph5+kbOk5YOnt8QKGGEmox+QS28beZZk+T23V
filaC1clyaQsVe3nQ2uHSB46Wy/oCOYjNI39JmsjK5zCeC9YXpGXq3AP/Pf20dFgE2pdwGNHZWz9
9CRxU+b/ts1uyd8W4F0dpw3Yj88BTQW/ZhOYONdFePA5QuxEdCz7f51fy94XsziGfNki7rC/np0z
qpniBOuemcvkIA2uQZMAAd0WFcPGct1FI3sAUU/aZj0RJ+dOxhg4VdoQ+Sd+EFuMTnx129UV8WtE
uwjlJSQBTTbvzZI99bQPPV7kay9oDfypsNCQR/3NrRDm0ANRY4AQFLMcynCsd9LXCm7wMis3S10v
xn2LeBwmFmmH2YZRo5YhL/o4nsweF/wPOIkHLwtc93Ud8yG0iTzrV5atwwNykAbFj9DtJAb0ypXr
LHD5ww+5A1ayZiZmtkwn+V2pCGJvfAjP5h0b3/NpU5nEcXrrkNQsl6sixncqRCI5cVJsdzjn2+k3
SyEkq2e6PeUlHC1KjyDS/W2LiUbNMyZrCrX0x4p2OWlfIfB2G1TXwHWGz57uU0dS8buQAKM51w/e
4mYhI1CK0YSswV8C7YgllmWGYQlPemCQ94gJvaBlOjdQ1rO+bFIEv9vnuf0B3CmIxAiLRzZ0nu/2
LIT9IiAi/vAwRAFPvrlq5QsP+/mpqADru4sMbMm6bSHX/WHJT8X8MBx09YTz0U/B/hVUt2ObtCoK
shmbdC498Q+qfPvd7VdZER9v7+EfyOr61xpzALm1Od/wqlA3FipqZqoKpgRpuXk6+fxrAagPWDBc
MRK1a+l3HUl+o4k1sHg5sVgrLlxgyN8TMvN1AeMTHa2djMy4PcCqZ2nLgIr4IpHaZGEOAO8+S2hc
bcjqUwSG3UF040QhP2ROZLQ379gT0iQl3JwqLZ4e0Vk7WP8bHDB6MXThUHAqJ/+qckhic+hyVexn
n4Ab6A84UIPo8roJxeHPAQeYJfjSczKhKblacUyTaO2oZgqlVB1QAtQARrdmFWGAlYNqwZkNeoEI
qcjW3UoafHVdqqMXqFz1G1WzskWMTqFT/U4jBcmpqfrIsbpNajYluC2el5nSLMZ6CAXmEfkH3vrB
ss4oxt0nApRuI/emz/EDk/iZXf9GNly7GTvDUc/xOUYu+qfRDYyGU91FsjOIQsVMzQuT30YBYbQj
DkszxUb5ja/oKLnnbVad12eglxAhmyDHFn1bivhfkiWm8SCe5CPpWNRaVwqzia+5DJtShAy6XIet
jIrKIk+aRLPwEY+lnvR2Ikyo7pD6KilWbfN6j/axxJWetdEqCKTQJZ+VcUWKjVoWEbNVhcaA9yy4
50VjBnVkkOLoVcfWe0gwXSG1KwUlVNzTIFAHtNIt2P0jyFuWT8ih0udOiekD2edpy9i/OSdFwyz0
k1atehCD1ych0xipaiFjPnyb/kYJKWG6FTvNtMOF7Dqwp4gHEwMKFK50Ylw+O1yofVqYRG3G7F5x
v6u1nxy9elHCuh+ATxhcx4/lGo2JnifvHws5uxhLlk9D/ZsAjtfXOiMVgwKnAX2ymuEarPOHhlNn
BrrkZrIsjhhivQXeG0Xw8FCTg1wcPD2YdjakoXCZ1ECPFfRBL1MHhFxRTR08v1YMe1MOSzCNNSl7
D3A85ZiSlUqaGRdskFNtC8J79OX8v2oo+6nYElBvxzxPVVZ7qpxAk+vibS5Hy7KfFN2SAV34bRQU
U4Ft18H42/n//5Mir1dIPfH/375QeDOAPmTQpiEaiuQmJ7oGtlZbBojTARsAFFoPBHlq4ytrarof
zb1VwWuTfglQtLJTK4tTL3R/KVKzsgWZoNUCkW/8hrG0kDk+Btkxdo+tp7LbmGnkt9CWvdBJxulw
VKyDz1PvSJKKaDsxNi4u83xlVc6xAITrhasgetklw7XOZ3YAZDghbf/bARrwAHm5gqn46VFwmDQp
65CBRJIcVx+MH8BLJ688xpv9fyXDN1vT7ME9SCo0xMpGwP+vQ7hMDxlpFlkGPNffOhb7vUqyJZrc
0vLxWwVjZeoWNz3h0Tx/v1YFdnjEnaeohXqfGBxK2KmyE6mBvbgCY19v9C/q0eeAIRNbPmq08/WD
suMDdC0N2qjd3Ji0aqTYQ9Yh+TyVGGdFqdHs/aOFzoI+qq81WpxLxNw/Wz6Je0V/pEGo6s/rtXgN
JusI2rvDta3Aw5OUoabw4KE3ebxJkwZLb8fKJIfIp9+TyAciUT/rEOrpykh3WEOgQuYRaQPGhlNp
s9BVOlHINk3ryH0+GYxW3rLLtCPt5mmgAwqHkkGm0dxZqJ7NqZLS3ncQAOYw4cgcD9hGT9Bom84U
lM5lmkoXmZT6JsEDVw7ficiqLFBfcqzCsVJCAgGRjMuKcKKdnTdyImwlqqpqhtK5dELK4x1ysetu
0+VQ242RId4mEcJ+VCIhQ4aRbAWbXJEVGfH8CDfV6ZVZjN04G9uUJ7yQZTUiV4d7h0TZryzAyGWo
6jWxJi8gYRVXodmUgbOSaAG1CBd8y4znocg7Up9ci/BZz4GfHvT88XGBQVRTcaYJAHGKUzRt1fO8
Civ9qwt4owhLmo/AZilcWmMQyTE7S3kEF4BI69SkuQCFONSKvElv3IUWz2T81ehiUz3pynP4Mcj7
zV1hE5emaHswtlrVIOnPIkSPyXq1EkBQWEz7goTtOMweAlEEkCnuFwl1pqdnJ5YHibUt2XJjo2qE
/QdpIo/60osnOcDE9Vx/AGBvRavYANcLDbpLMB9MZ+fvTqSEDlJvCGiOPMN5o8iZ/x+nyid+h4eH
c67UR/wZDIfH7TecR3udLtbG6WUYN6o+Hem3eQEnhzMDVaeAXEj8Ryv/K7IkCGfOO6OXj5/mC7Lh
kB6mf8v2CK+cjK+Rv9J9slHD3vis3USN9K7S4ZJoftncPCaaay3il5iD/CpKobEAWDDO98ggvTg4
RZbqUCv7B3jJJ7xQiKmyioXoAlm7//2vlbLASWQaIr22eWahjyh078thq/wtC1JtATi94qDFqOQA
8fCf7dyev+0sPyhDtYDGXqdoxBaVNejpV3v6HQDdr8IV1abYgKhnGOAmjwJSlDjAfeON1HQ3PaE6
vM2GS0k6ejyDzM1WySLvxtpWJ6VO8x2jmgOv0AV1A5htzkgI8fJzXjaSgUF2k5yqbF7H21cZmWHm
W8ZgUBuiT7TRmCrqYqovhoSGA3gbtVLjwGx3RKRT6my5PTkfek1qxosjQy4iXW8oPPsvwz9CslnJ
cxJaJavSV2YBWKBzG1Kz0tgX5lVhokAUOqm50Go+NpZhuZ+qjCLytBdPh66XNIovtWT2MZXHtqZR
kC3Nm0Pk8U94nyMQQchsgC/QahY9dVw/awMPeUARyMz+x24AY01+NwYJccERXkIa6CEeb+zxLrz7
q/Acx87Eu34rNB2ogKEGkOVhEnTarcNjc0Yf9vJeAWVVTIjcFpdcv1Ns1Q9kGPgP7Jx1/VnCZmRY
dj39lWv9D3iWET8FvdRhpUy4b1DSVQRsJ4VLctCdXb2JMl0ImH4y2OiFTQ9iiyBF3iqp3qY9A8yu
eh1k7uGFm5+evD7g+Q+bTRvTcdXIDX1jnfrZr2Dwxt8UwM684cKTIawwK21L1vXsWOdVihq08eYJ
del974kd4n1Uo3c9mbXG5hSls1XdHaIfhfW9PIXWq0MfSKC9GxU+vmUcn49s10VSJg482V/qmZeb
VXsRBoUzOM/BEfDBg6ngqlHaYi1Iats0UwDSUt3n1VAJfP2OXuUZtk25NORE6eJ3Cfvmluak4F/r
0rr9YEI8Rn5EuSYxkpj9H53oL2irS94Q/c4SBNJ5dEi8OXEZeta1fjEkF3scw2Oh0lHa6unXvoLc
Zcl6ZCGpVY9AfB6eAhRk09NTQSGOWZoGWFoddkOJ9+lSon0rkJi6GAYXxuAlnKZSPvDcHjVNojYV
yYCy9ab0z48mv6FrRqgBLVh6dQgbTlzw/sW2QMj7WYOrRkfE+QTN+ASMU4MjEqZW+ayfjd+YkhLu
FLrUXKBWqPl8nvZwevXyRoqmkM4IDi2TpCESLLXfPOg6+HOv5zZ1R/uhZcYBEyndgBO/pzLEPtbb
I9k79azTQqgCjyeSqz9xEpgEmt+VQQk2QW7vKzSPXMWIyKmtzmsZWU1xSM7NadI4rpmJvLMVHrpk
2ogVN2Rkr/v99EH/bny9SXhofAZaNpu4trCeMh6c84/ZeZvvoG2k00gV4gD4v4JTd5TQhZU+g8R1
YHNry2/9OPK1Y0AyyczyvI7p4Gde/CzKl9W4TRf97e06dOSKqC1bhZyA9BOiblpiWo8KEz9inyg9
3J09495h60F76ljbBQwD6zmd7gpgvgejYiH0TeJzAWE5/PQzrUvvuy+/iLBBiBxoMV9pxcHSuS8z
pYZAXXJPbslo8paKAnpN8ji0laJYDbKqjQ27H+nrF0W19hDxCxhU11oqkABeooz5NMDF6K0cAMa6
iSxm0dmhBy5OLkO90AIJZRAO34ztmkWVXvibYU/1UcamN0fpXsIdaQ+Ld9nh/LVb5ZRkOX99AqIF
CRJMBLPfyTmOJYKZx81+ikfStIw5elhTfjg35qKGnHDpc32offvLEKFbXodAIwRG5RaX+4geB9xa
CrxfB15QSpo3Z2EcLPuJ35hRe0vXBkfvghuyEl24YMiweIHmKdOlq8YEBpN2Vm1/VWYtjRvAmBw7
rfuqqMMYDEbXx+2mUmT53iLYRtlmS2FMf3KkE1fwkr3tPNheIsV7dwPBAFE9MgaWRv35Ku/qmN2e
5nBfRW5Jjxz8BFlSCjbmwUxacX26Th+JQ0dRge5jpaqQOWKo1NvZEySh+nX8CpqW2mzrDsgWrcAX
TMYWBUgBFFrUOwsT9ckcKjz3X6Pwr8cSln+9PWkNwCkteGDvNyfSCe59uomQeSvkuUd8Xhd+oLml
JMjz3grng18NgZQYa+mybO5x6pD81ymfIel2V7RRbGYsEQwVaqj4KzZQv3hJqvA5fpAZvvxJGeAR
wJg6icSaLOtGcwV37c+ZbosrTGDBeZMzTzfdKKMZ1K+Nw+/eUny4NTLN1H2i5YQP2CSrNyTjUM/r
hqOIVCvMb/cdmYStRG3uqmsSpuPZTgvpfKPm8LKl4SGF51/YFjhEDgkrWh0ZNsQ91m+//LyA/0MI
ciOSeYJ3IfBOGA6CPML3K8cM0SvMKgfQzxS+AI9BTVfEptPXPAJhWOoYSrn4q5FfANj2dnmYnojE
gxdSLOUOe26t2i1yuptJhi3BF5XF97r5vwv8JYjvniOFrbAHyK4ZemQ1BX54DhRXd4BVPBotanXj
AB8ZMonP9xhMgfdHg+h1o1fPKQwizelMtBHkv7UT2OUMk3znfTEplXMaoepwH73kENlu9LtDgfEE
Zxs13UIfrXGmMb+9IkkebHQ0PixQYKN4/3vYBIyVOfl4Q68qU6nK1bUZuSaTPEx6DNNLtHMdOtPq
Et+sE+b7d6J3s2UZoAFrLwC9qIwAlXCahCpq6MTLiGocGCN19RbFUFKvccPeGoCp+c5cBQPLaT2x
HW3772cGsaX5a4Sd2TX/fozMBV44rPz82am8P1ZDCCxoJksusMOgQQ18vj96J/fs8Xx2ibn6sFXF
4kV72PkhTy/3RnlTEpMlm7JOomngnJ/lkMumlTuOsG3PR7uxBjCS4b48BBYXLIMmlW8rHRs9CPXx
29voTCsFdgjnxPzGL6ese7AoYwbWUSYTIm8gxLz/G8pSnVQh1x3UyVq8ZF3eAZAKovnpSsn+BZ1K
v7asNTdbTIJ4475sxw+eCrPnV2BsSzJ3MdrZ5N/2aXSi9WCaVImmYWvLaG/OyAt8qm6LMJ8xgabg
imr5WnM8n5EK0I/wFms1zIYyPwXaIp6gB9KNliLtT7Eku21zx8mHMvkE3ueEzmhz2Qvd6GwgbglV
IdPuiezAbM3cY36LYe4ti2h3cP+BmOvKHT0es+OKpVPWyF1mJoP6fhvJvRrz80UlpLMUCVdf2ynn
V9pHjtDjod7JaVkxoGma65xiagzWuE0s8ZIQAxbm0Vfl5eqIctbJ+PJ51G+2SHjYgG08Bs0n5x6W
J4eNcN7yURrfzRJW4sh0nLhYrKXi+VYlyWHoy/HRDrWw3PUuBxjMaget1IRg/F+UK5DozOHoecuP
CJbsUXx88myTkx8juCTk0Ol/waN7C2dQ13Qf88m6zw8nN+bCS8mUixYFERON0SM7HgwJCaQph9ls
tSdktJ4SozA2eBcmIdBeSkejJMaqMg8tEW/4fI5QTKXlZTLJ+jfh+T6kPjieweFPe4IabQUQ3YCF
8+p2DbD3dwpThx0OQKDNDLKkifCJmdSilUbCpbvc4SwAenF/nSLm8fJl6vQEDO1JiK58IGQR4ync
0biDZ8WzIDOxRbPAQvkb8GsGiFDa0V8k/AMqObxg5CaNUlRAM7M1A1D605FgCzIM1lw9n9h3Eg5T
G4MRNb56247YhDpExrvPcpzvI3UzsFU8U8xuK+w5DPZiwxicNc+vlP0exG72kxJhCNDQdnVoQ0rS
PTfklw1/Z7opHoeA7g/Z+0ZZnA+HCRUTa0WbRBqvOdPK4kipJa66RD5+iLXrr5GCm4dSJ4jelnSR
ff6yVeZZmVQbxEvvXI8SoXJJA00fdaZuIg1+1RoncxkbIT2s4NYs3icFaiImEorOU/1RbJzVyjGH
hY9SUkqIK7Ym9VchRFEN1ybpSEklWlpJDC8dYlTqnaQLOLQffvke0Nlyn59ihvER/z0RC7ve4utN
3V9z+2iKKpAJCEAx1YTEgERDh6w62Evga13bT8zBESVrJpMsSwnVWerbyIoqioxbeb3wVlDMVnZ2
WYHXUFxGMZD48WjiDsT+2yz80kpQan67nPWwuGNa3OXQ5UWL0rVeLuQcLaBLbXXsf63zpPiO8lsM
7cQ+Uiw2xe2tQe0JnqdiGapmF+N757bsurW5gtr/Qx+CkWgVWo2Ej3wua6v1jtnG9BzOXh4bxsD3
bCKzf+9pB6R6YT56tpX7raT6Mc9+gHFmVM6lM2t4hqd1sEW/iUZqfOxsDzEu5WlwGoJpQiC85lYV
RbLqRFQ0ilOe1r85GIns/N/27O7uoiNBGl6eEKZNNNHaz43oLDtUKySPChRfnkCQKJ/LVrghxW22
Dz8CnovjH5csHWAhv8uzoZNmbmo9q9DDlhrIMrdpq91Z5WeOQBB0XhfxFm5EP4+eu6l5Q4vboOSu
kYNsf5xmiS2St8Va+kHd31m/tFRnfpb8amQrb+WyqRwypp87Q6I6OG8znKum2TdsoEBfViFuAMwS
rzuutdroQClOqyzT+bUzzfxS8S/fIbI9owZc6wEoUerEMmggxLhP4ARSME+NvBIJ+/ZBraPX4NY/
82CNjH9ZX2nz6ZnsqevRH/MV5IWBy6wLlq1qDMhfrcoM2x8tZmi4BBdbXROr2DRZ4foTAEvaOIX2
oVJ9T5iwXSkV6LxuklkloJ7S6bnjthauAeRKm7QVWqBRDI6zPUCPcK4LoJUDOOLtebAYhNz0knrJ
dOzYXCsiqjXylayXlLHXKpzUNssTNbI+aXat/rED+G7Kxoqyj93tZd3SVqHTmP0u8PNlfyC1toRG
UfefyIP9fylfxwDCTg00MasFX7IG6nIMOeZDZ88Ti228DcTNBl4tIpAGqlO7UlI55kdFHgujiTOP
196XFMfbZG07t0sgJ6Dh5OejjCIZKCJJ4nN8DANHsdtCChc7tOZI8NKryZcVMfxXPIdlc0CPh1kM
NlUpytt3o3Qjg/dNf2HDkeSkUhBV0PDPKB7q3JfQeInH+3K6rysVDxfRN4sRjhBlEI+c+3EyVLG1
ibtK63Nq6HoTQCcnQMtmTcKKIFPNjGiWx7dAicEh6BBQ+f5hJiuF8m4OkmD7qwFQcubX9fAXdnbg
e0eLg9R/0ps/FvOlK/NxXY/fXmplieeVjopLT7q1ccpxj+bwx53mUrhA4XqUJrU+pAfxUP+ZClf8
mpk+qywGAtTnFl454fxwlTmln7TPnwvnCxaQ2dffahlRiHY8VtTdBd3kyaAcJKNicVKgof3AOg8f
EzgbgllxeTlXIqD9Rl40zNiBSMK1h3ffIc8DfRx583CcccQOLjMQiL7g38Y7S8OprJMEhCzZb7wf
2ZERD8uid8BvyBooY1Hd/E5tCJXnGMuCz7YprqcAn+nRrtLPSulkdeWLyBhL27oiK+6bsUXmtD/7
crkUcfqZGMqDTVTmxUX/ttn4FasT8eN/rXWXbVcP+97eDyX5Mo1E51tdUGwF70qEdPMx4gclqWPS
ShvwmNgXi9yaYeIL9EaNzi79Xi5D5N9oJmB3P6sp4PQ/jxRZGUJsXRMzwsg5shAuPbeozZ9anyu8
iF/DZDripOQDnM7zmT3PSCenKNRyLTAXVT1LXTrkrBwLl5+QU+lxgYlpLUlrbR967zXTwxNZBpRa
X9xlCxTe9I8+mY9cnn7VPfIcUbV73d74lyR6hwI7rpKs4gA+s993mChbucR9Kf6ON9YWCXeAX3BT
tTDO2lahGMG+XKl4UuJcpUp1Y2ZOpm+Mxu/CwPyQ9+KrntdFg4l0SoJ6pp8BZDiSy/pkiDVhJcQT
RNP06Jf4lhU94O1isR4tvNIETdINt2BMHWdJD5iCMgEI5F4NXGTm+D9ARP0o6p1ySmAWHa4FJhQ+
pRhlKEDW0G5RhMQLfAvhV8LUIahs5XNoyKsMfszURxLWoNZKdfaTpLYLx8PY/Nw+gnWB1KPjzeRw
lYhjm7FDRyqgjONxz0hVeXUZNlyQahSy/8H8Z8Ugh2sac+zJYDdF5VMfBJ6dIlMscpW+OTkjnuZt
yO+lx4vZOEMnIYSxXwG+vhKGBMZIJquTS/pXrM/kS++/1DrhEMUju5r+cq1KP4PqM0Uzb0iNRMzi
UY1nX9VkSfGMjZxF92Rla8ViQvnfuKLlrELFpCDlgwcHplFyPFqbBTKy2qmUisieSw50nu2ayirw
85Rr56nC3Oj7mOx+Plcn39euUjFjFxdlRCfKBAIFMelOHbhhXNl3SNDN8Jkj631vRpw8jKkIuxiS
HoOH61hTIiV2ksj1hdXmI7UunmMbCVG0Bp2Jnd0j0lC+iLJict5oLCv65IAvTgmHJxIvfd7r7ieA
wJdeV+4NTo6t7aRriqkBy5p+2Voz0oA46fQ+tKbN4I0RjQDP8v6ziMFf8cVo+00XASifBCZdrC4T
tRXp4kouz6H/5eIUilDg3Wb/q0GTdWBB84QvgUEIPuar0oGlDdNNTuNer6jvP31n8sNXQzfHphdX
a2rRi2pEBxi2OgOWsSh7B3f5S2dJpmuoWzJ3ea5QQOXyTBUO4vxsbFYMd5QVOxL7C3C/uaJY300l
FE1gBR045jyAlNfP9f6jCz9tx2LE/bYYWTkDJkG5hmPwx5XPO0E9wQZd1usU9eJgLH8VVEKjjKTK
uGNNoiZyb8SrX19VPOTqkr3bwOd0ZiibvtRKmvHmeDcadeQyzJ5N53u7RQVhOzsI+tdGlfWe8t18
4Tqql/Mo7aombJxUmM/s5S/FqMbSv472yTm0Ia4QxTsVBMLon6uyu6Wzl2Cv1RRTzJs5Vglm/etu
YXOboYIfjE0aJMdBevPsAQgyLyUsxKSt5wNMvot+AVbnS3O+2ThlpOelgsmgsHBvKFU0wrM3C6mU
ScIs7NvZumoT/qA8/JK0cDeCWo+5lrHt+q3ofrdmyj3/dxufTKlft0xly+T49av71GwVS4L5IaBO
3O9pvQ34XV/x0XOssZs9LFBe/T8szrz3+nHQtQCfZSBuLnWOcnEjNMiPHiSV28iTuHOnSRihmtog
NqV3OIrpu3X0PwLvJcOP2IYnGINw8/T/IiE0EMvSzYI5F8zkR8HzcTZ+Vet6yaGZpWcprT0J0AHS
2VczjLr0N85dhhHFd0kjOZbr+sjSG1pFKDVcUr+1ii2oeS6VVIalF1rmPtfZFpeoT1VoV1lJj78y
KmR3fiqpp4DAyjd5j3rziWWSrhFGZHb+Q2aVWoH3EpKphGWoABfio1Eu75zjuT2yimizPS620LVw
oqDx9grUqLDW4vCrBZQ+e5Hc8ib3fJsX8PJJM1F04AJJ+B5hL7knbbreOQaDm12m/jnxP38O2QGg
TtwumD9GpaMkF2GoblDr8n2S21hgzHvH4FkpTUFdCI5zxfJUTKXoM4/GcofKrXIntXcqnInswEGQ
9HlxVx17aK/YG7A/vco/2a97CWqtuuppsHh0qCLGIyjMzV7Eugsen8cx8cev5q1AI/8G9AJ1VG/h
DWRseNtEKfOKwUGjc5bPzKl9R1csFfjj3GHIZNgevr9O4Gw6qKT3hTljGNgXdbznBxlhRw95iaCV
kvUgGp6ep3266tMLcJpfD/9E/ElvDE9WZ38vjs+LM++i4B5Gqrlv82bQYq1OKtLTlb1V2XC5jP2p
Now4UFTTHgn5n3zZwPq/PNEn12Ni2Qsak666Fwa78qzOn8rOlnNI4E02l/bkogMWevVQwheJU81U
q8EhkyWPDzrsR7d/XMZ3RjB3uyRSXa7oinSRyOg5UdkdtEI5GskEed9ucuddltzDN3sIoOV7dUpY
EiJelRzP0ok6PuIm6KejR6G4ltAxOzAIm9Cw0q3T6VAIdh91PuvO6zm3cPXQx6NBb6PmHbwwAemW
M/eQoDzF1NSeCVbOnjLSWZJgulpmPV1+O0nzu4CT0dQF9qG0veb+M0aoBBgD1DG79Qmr4xHs3v2Y
Ixsokqsc/viOfWnULdWCFfAm/ObNaesVyrpycJGTR4MVKPWmHCIn/H/bMQEOblIy2Q9HEEStd65m
MyWiHMUch8V+oan7r3R5ZnwTKoIQRMKvQUCyHnAZOTtYXX8o9DtN3GXBkkP3gThRHVvHBOtU+sbg
xHV05gMHU9bmjuP3gG31FElDr0xxuCNDSOz7i+LtlvHnUFfLt+bGxIL2pN2+QR/Cf6ghWwPdhlpY
8zTDMIgASfAvf6LkEtKiqlGOH3Cmuf0zDOA7PqTyyJ/DeKEAiuIjZHaoUhElFfGUqayL5pYstCeq
fIgg/zideRXanIWN2HctMd0t2xPcdfdsU5YpFcx03zIJl10SCZ4HifSe7Bl7Xhwae2nc9WA6eA5P
E3aLRMY1eCPzBTJ808dl0auLhdMmEK9Sr0zb87cSYG08rNTwI7m7zXzGfJ7IOcgXC/HhzmxB3FnB
N/pGxtMDqnUez6b8bP1iZ4tNV30jWrEYxij/CQn70W2SF9yIJj/ZIQ2pQOQwuK3t7l2S3t1ZfJeg
gyUtnF6K4DuMJ574SA2jWjVwR7aBcHxmKHyHv3SZI3MrCmo2S0/WjaLuj9wqs0VdmCgeS5TJdyBE
C7WPvCMMg4DlJbHVCodHcgKqIpmn/dplEWhp1iWFk1zYsFNRLkAnc5/4KP7LD2RRnWvYMyfAWz78
KzwEg16dJx8Inws/JjfR08VkDUctM3JyRZGSHwFvAlDNigNjjJm/q6Wl62m5qflsG7SzX1J7GJqZ
B9O8K447M+LmDQXvfudQwkWygMg1za/YCfOunTWur3tjOHvyyPCuUUcwScs1UJfcMh7HDgm7UZrP
NJxqMhGUoxGbfL5AsVwJ+7f0JZB9lQbc10mywVzDMyMi3uMk11R06T8jGhcFuDX34n3RrN2LLft9
A0X9zOjooWlh5Vnugn/AJ/xIQhOb/N/miuyY3NR5zGx290NLIEJXxggvYZl9lEfH38Zv4Xm/wvwF
YKkbOEC+aGtDkrT3vbANScNdqQquOGv6y+kB6z9Qz4vXmzD1NSREdSIJc09v4kp0r6Wl0yd1tq47
gZeQQvXFOLRkbSmY7CpLfX6XMWA8dHCP9hUKQdm+4F2+2VUNiw23Hh4CIgox8i9UlcLDIonn7oC6
wY2N8Om5Ztn1e/XgCEtcpRlC+yxzvPOJJyEkxTQ2H9ow7wWjaeZC3lrI1hDEu9osxxSwFC41PQWF
jUu4iUhaMu0q2j1mxGjdMQqlUjt2sMYWz1m34wctI9JNkoOmFejTQQTtpvwUYgWRfeUbWhLE697i
j/F0trERTZVNSQXok13XwCkXsyPZI/ZFXfptBo3ifFkOBQ0yfY/1BkelH3JBoesWQ6FK8nsn6vS5
xPVWEO2XaHO9/d3tHtIS7gbcld/VgeYQ2voT4EBt+rdasojGEssQFlr/fmXGXtgU4EMCJB/T/JQ2
IeGUbxP0rRYy9nxRyUs9W5gD8gH/41XpER0scfAf1z6knO7hxn7i4mSyu2fAWt2mwtBKw408OpX/
8nGUW/JrARiLJobG5BM9parwhr/vylwtZ1YFjPNHQL4Ey4HXd62fCNAt4cmhI+T9Pb1hFMN2GtUe
CX3oy5tcCsQCVkv8OyC/eKj5NMzHEOpsgtXdBlTqfGUh2aTYmzjZ1cLaVRpLoVebsQzCVNFn3z8q
p523DheA14ijbtzMREJx9Wx6a//fakCN47i+ZFFymwHBvuZEzOxrzLA3eKakR6VuM7CguXCX9Jg1
ceVXxapPcls4sXraxv0OmOJW1ft9lTzC8kewihpUsY9G07mGvPDlx6oND4AoaU/XAB6bDYeB3C0S
YPZGLRMCnxmJ9XqjzJJTICq3WmP1poQxTnp+H6JYa3bkqAMwKnAKdPfnuOInnQwhFmQ+9vWOZ4qc
QHHZ3bKoO8r9sUy6+kCel64uYXnjulWaSXJ7SY96sWIfSLRJR3L3C5/2zzjMEluSF02jJu7psP7I
vsoaqKISat2FZzcSuGLMZKZD9Sw+5U0aeVTo0IiWQRl8cnsA8KUIBgh3BSLMkH+37ro16fxCHGOR
dVt0oYBdxhRCMzRX0xMhzRvUunG5AprU9Of8igD/nsqblYVm75O3WBocCpoPQjjpMkneLrwbsbmC
jBK+Y9/U3/HCsZ86rAGxfSaWlt7EkKu+AzkGoog2nYKCPeauEhoidpO7o39YqanKU07bC5o3ih7r
PiMFjuMqhyx398rSh/Szsbgoq2ITKuXPN8IhU27gKz/XYFpEV0gjwhCnLW7IJkA+x2H5XoddXqDi
LhW6pkqa7IDGi7i61JQATo/glljsr/xcpN0ik0kia/BUlpUFDxFb6ppuRABvbGgFuQ5N53+S12Jb
W9IYWV/2EkCBumue/ms/B2xqtrMlv+nUf/mQIE8syYQFM/Em3Man4oZjJcGl/gI3w+p3qK6w5QYV
IKB3r+y1zo8hLJsc2TLfHuDDDB/M1qrF2rBYHMTMqE7C8FANTsHl/1bZdzIrBh0NoxwmgFMQtMqa
d7Jp6Cxd9AVEeFTqsYUQ5f4rUjbvQ1d6A+LmyNdeBg/KCyOwIK7UZGCavNn+eDRe77yGMHcON4qH
zCKAC2y+r73+3iqCm9K2FJ/2OcvupTEwwKIwfD9Pbr7J5Ww82OjkoOvU77zwQdE4HbsS1BWJZdG5
bJ/unH3Lo3eBMY52CHTk4JMmTPDcuUSG1n8qhjlyRHL5mRZWnOchQaCMX0WQEexj/ZSOAWnyu1N5
dfyVpxAGOvifMzWD+xnP8FdJE9tAYm29DVsu8gzUMTryjQvIqFLGKpTcrixLNhprhX34rxDpOqSD
/g+bG3F470pPQd5ByluhrcMkW5xj2jGx8zCv6f0e8OpkLKWCdWRFrqdzPLY0lHlcbp++RRG9hWQl
FaiYbloK+0Cs/hByn3KhjR3dgS3QmxKQXPiLxlf99vzDwePRo19ytudeJQOvJtXSnEEii0jjQTdW
St2XKEJEfQ1Czb4pI4iXu8tMjulaKDqjm/ZCsjy/wbZQTB6XwgzDNwUEH+VVf+esLTL3Yo4z9f8Z
cUR2a4JdNcNPv7zClE8Prd7GCVpjbB1hNb88ZfTZVvJo/P+BJ7lK3v5UwqI622Qg1RjiDXtgyzgN
0tj1SFDvz66r8IXULSj/P41cHzCY9HZr1fM1o3mIhxPTecOL2gYbM5gC3Xd8dNRGE/0cLdgWGyc3
TViUGSnI44aSIgzsZiRdEtDvSAwb45UDwarrEGp+n9QB1OD/gNoJwH338NKH8x77gH8cXEllqSwN
MuHu5kApzBbv3Nstqd+PfhsnYeRJdwkkbnLtWxiTUuTxh02OOEULFVTH61QlQqFRHScvtiYkhYFL
BstS/CE1LZ/nc186DL7lsH0gW4VWV76Y/zY4BepHH0dijX8Z7y143npaXp81tgg3xkt2XPYe+vzH
MaXJVuJ71aetJaqfW0hZTkY1noLbDBzbs0QxBnM4cURoroQnQ9I+xPVA1aSTicmE5H5Jnr4t2hfd
u45bqEAsct6qfgw2r7yNGyTyXWa7UpIdAmZWgdlmBHtNoMDsqxt183L9NOC8obxPQZX6ov8OZjjb
15urJJWAYc2fKjfX69di67zw+hlOXlLbx+cEDARtlWXX9is5qcj6LoiXE3/pqhu0+I26BkxyjEa9
9ksJPBLhrHRHROEaF0Cg02qzd5vas+0G7KecuWxnXpT9l+6i/nMDVbRRIesW/P7mnfCYmCZZEVAE
fTUuZrFYfTY2m+8vjkZmZajfwGrObzY7Kp9RMk/EZNIG6hwLKvZ2zlaphDFUkkM9yzm6V2jKfmhp
mOoA5WkKZoxJsk+/EYr9XwC5kt6Q+1WPSUW7Nvj3Lrir5EskbzHeLm9poUQ30P8M9zlwPUyx1gdt
rK9eBeO+xaQ2WKVIJwE3YPJvq4ooVmvaw8PMzjcgn9Ctk7mxOW546sIdkONBxJiRqftEesisItMv
kpL+g+xEMNioWZGBh2LHdywqSMNzlFv3BcXt6cA1bcJPgSZtdQsIcFg7/SB8PugCkGkaB6vz1I98
eK4L0DNzGuegyGK9TFnAn15E115HPQCfiGkQ1UIGP0uANrfi/LEiJ2rnYnVinb0+Wf5lbInLidwT
hvfTZWPoaGbIL040C8q6puR9E02821RKpf5OEi/pzbK6LFIYIkDk8jZqx+IVPTfukFDV3ac6Cjg9
I+viY0TppuJ3fM5NZ2c6UMEdv4X9tD+reebboXIDOjmdoHSAaXRGtqV8wJa9I9BoewkFsZQ449fs
yeWK5l4LZYGfT2JE6a6mvF5YjQhNRCj7SUK5nqH6nE6tv4WLBGWMgT/c5jvTbc0Aw9+ojbZBwtWi
2zPp9Z5k7bc7Ah8CP6P4pRCjEzWBl5o8QK0dW50xzbHfNV687f6vdQTgkAlUcQMEEMvDPYjeuk9i
9XZ9nVwZSiL8J9BFmWxeWbJjpwgdl/D3mnTORLfmr6XTz8aF853YwSC+JS/cS/bRA415IF6X8oPY
Uo6qKNGi8tcsseb9vtPthnUbAJnnY6fl6wtu1aWP/rzdiGVn72lEt0/AEfqBQYMBspztNA4PhxK4
re1IFSxFT3swMPHn5+vAyr3iVGJdXHbroVvXgEyQmirLr2P6Ojmv0/lFLekfj1yUjv3tlxBGRXOI
tYYHMllrmegJH5K19BzG3q05TqlL0l+2eiOX7vLT0322MhAxjUM1lkKzsxbm7ipuZuLclDyAKHOs
9pON4OyQvLLMp8DUnX+jzQedlKfAlrZt1uORHYEjLTbYvtHWbcEX627VQ909wFEUWhPJ6eB9V+y2
EVv7uOAyb9s1kjBh3ew4rCS1KLJcachziT5/Ayak/II+atp24A6JGUdvywMMT3d/+uea2e4S/RcU
XbvcebwQjLo5K3nvHaSrSazEDMtqTOjEdvkn6rzBDgBbiaCyZzuSEhWV9QX87QAz2JTUrFu0MTpL
FFbgq6Mmwoi8ezQjOjVdAke5c3w2hAwJu0eSCk0/2xrbmNZz0QqyExxb6mdBAHju28YI0co9woBW
OZ/5PjvKZRsfvz3OjwP6NvqyxA8y1SsUe5ESv3hd1kMHLCDyFSAUTx0sjHE4y0aPX0kQpOQ1Esg2
tATc8GPs87KWTqwaqKnr1pjbWBzQGa8fZW82pKrgjFnlQ1LsRmD6Pd3+OJAz0GBc/m7STwugiFIi
tEZ470tiiJEyvXUOQ51ADCFgdV7eCseMBVcXpgsuQAUWIQX7lm9UyeSuBJR83yOtyQxdR7zU2h8X
hI3Z6ECjVzkbA+/h4yxImTrQuth6jdTiK9kCRUA5MNPHzF9yYy5oXGCTVeES9HVAiU3P6TXcsgGf
Ta/9RrrKw7Z/zakhIu2eyLywtcb65OdB6t9A300X0EZo6YgesU84Sxp915iap1WGDD0OucmvOPDH
FHuc0zxJK6axQx7d71frIzx/GhBTXEwJ3zSFondAXAzMUv4pzl+8r/3QJlFMOCZs5tg4PYNpBN9I
QoOJbDQKgR4Zpg29ZemidLto3WKKlr0yfuCIkmDKJRjBy9SyvdXK9bMl8TOtnq4WS0UljG3BS/E7
WcokhjEn9zIHkzPBCXBjLMCjId4Yh8hCVcDT3dI8V2OwBT8KK+uaP2etPbQmbaREyXHgyf4VyAYR
wzj506R/8T8hQCXp47myTUqeJxphIxJbR5wEUvCQ/u+iS1+7kSpwKklglPaIv42KksBQA9gnGPKb
/LjSsZPcMoZa44CDUc5R8vyvXwvHc6Ysl4SkZGGiR2vQXgiRukg5v6QB9h/8c4d1YtX5HHSgVDEm
oWDnH7Q6Vx0FJxcLXP0uNi5ZJxOUAst4rX12ncZS8Ph88NbUFNngykCGnWbB0eOZzpgKyb/yOx1M
Lfs1OriGwH7A04X6KIi4MQ/QsNmMgcquxh8Puwr2xdXXJH5mCx140es1bdvl3s92mVidBNr6R17J
vG8+y58vdZ79I6L3o1ilKRmr+7tsU9W25Z8wvBJosJgTgSgcp/6p03oE16J+N9rqEAUBiYC5Vvfi
6xrcfICz2Aomrwu0VJRYI/L2IM83mFV1sK4OOl/jzV51bL8zv86AKY9lGW1ZelSJMDe0ebVSstmF
sKLW3y1uHg1jB5Pyxe9oMZREugN6BHlEqD6W+74nbeEMbIDJM3PnQ4ThcKRs9wKjaz3Mf1xTlllR
8AmLjtzLRjN0OTlmfqgRJ4eH8WDPStUcao4UWwHn4jIaUqU7OVYcrrv7JsXO0iv9TD6W0vEwR/ih
Fs0cZk0jhNavVozjhK2I3dAq3gFtASF3cKdKeMnfpWMdFDj7IzhFfiwAgU1gOoI5hsseEOKkK7wc
Q5bVs1zZ12UrbewQkqAECnL7H2WSERcocduN7Oa8PGPvmQi0Ba4ja1sCUqY1CFCKKqxtiEjpU9pm
ZNrV6rcAImIs4eH5JI7a7mpCWfh49zdH35wiWB7I0mBt+v312oyMutprxCstC9zhMDBP8HTtukLe
GDeLpTXk824E0ucNeTYU2p9LyG1E8Z7o9Bpcv6bo+MtiSZu7zMFEP90wuooKjVzlxZJmqU2uDx/l
ZGG9M5bFgsgtAvPtAnl4TvNiUJHb8E1RLsspMFpBBzEBM9NIPWROXAHOxaGkAYgsE8kqdXRqLavY
c3TqCDxl472LPYkGwXRNQgg46vtUBBvPjEll20tkq/KXgUVTlFjoMDRaU+KnK5jjFLodGx7YQ21O
rIl87aLd95Vk5hXTo3qOMFzTHXuaeoKSe9lxBdoY1QMpYuDaZWHKtjElvQyJlGf0c+YY1ETk4JUw
vaGrd93e9UG5ajr7kScNZUDiSOd84bbuMNyx3MPybJsleowk3pt5d9d3TuV635C4uyXloFbCGQsI
k+VyzSmXi1cYaqs84SIh2vltAJqig5soZxUMzTwiYnCzBtKqjR+5q3wHhQNzUnAlKmjvb8AfqNe3
0LzsQXbvAJv/JUP6AeLbjM5aWOBIX4XIMNPC1JnBsdpEqvYXQy+HLgJruDBwb0INb8zHd+9M/2f2
obrmhUh/KSkZ3KOrbiMzdGuR+FtPj6qd1ggtnVApJOZYIy2KbH1JkykOUx07FVIVi09Qeeyz+EhU
2iivrVzeHmyuUhKuOcfHXrOBJIFDdG6bExddCMMAcD3m1mjBy3KoZ91A8syhtlp0nXTA1Vqs6Kyx
IgidHFcDffr4vaQrZRzktJuFaOQxOnAJ26Nr9TQimD0falNUpRXUjKkhIBNJYWPexkzXRLd7piCN
3JguuoHDX+cKkliW7DwiCfQEH1IgTSK1bRUIM5WwNwrO4ogv547sISb7zbAH+gwLSX0JqevBOIci
ZaF49iiH/Fob7mnE/mJLLDstJGUtk+7uHN3c/VGID0Y7/bXNGBeOmOfCpEs8a/fk+bxm8Z4lDS5J
GWuHn8Pbu+0jUsR7P6W1CdAFI9/lFCOEFFStH1TaBGCGrR+fg5ZeIKt/SMxUveF26hknYUY2ikIl
89xSL8+CsXdbBJNv4wK+S+aycQGyxSCN6GIuIO563vCf1u3F4HbBkoYDxmKiScdgkUXfoC9jRO/X
9B34EDy7bc0nJksut9hSEAhOTKEp+Bf7mYvsnx9a6GdsHsN41XGK0E+jDZbdCp1Pn0Xa6BKP374U
x/b27i1phlq0GXuu5RL7cBV5eCYZ9PaPcKxf8sFDz7L0RLG0QQVP9MYQslVjS7swKJlFVadKwk/c
QzzUqumAKsuyvoPYCTzHmGP7iDWzjqy4IE1Dz8uVOZaammouwltL3oZ8B6ZiBMktUVSoU77uC2zy
SqYTAkctWfXlhRT/6C3X8LHZUq72bldJc2wokkHjs4nInNSCU+dgEEBwvIODYv7/j/UgdmV51wHe
TOjgp8Ua5VZ8QJrCTLolXm2QN/zgTVJjD1XDg2lqGKdu45RW1xpXKtDYxmpnyveGRwTWPOfQwmrs
NqxYrrlOwtNFSVHSS0/6fa0UTLjlUQXz4rag1F7B1pO6FyyYso8DRT22O8rhMCeHqc9Mp9ha28uR
jQUy7ywer3PkrCN99u9z9lwuta/oKaRo0fmpmsD8YORLxGAoTjPeQ516XxSTniLNnWMUhMQm5oX5
sdKKNVx1561j3qTilO3G13zn6McYn8CnrsXJTbfnHlpksrBiXqCbOKExLhFAYoxboC2gX6AC7/Yv
CVHoqqKR9akY+c10xTdvFRRmm2yWZ6zjN3xpcFMS+hWivhIJVovAgOl1GAi3kY/vhGMAIaBJ0ZjP
srYNJ34ogJrAgabYZto8Rcq3m8PekRX69r4QLVDe9VjflI0rmPmfpJ6inMkPGnuU3cF9IgMlTFxC
6TPoZYIoSJXWNIlsrxp7/+3Vy7LIsoitwyd0vycRpC3iMNO11lnKc+Ozi9QgT+lxW+Tige2AYyRc
oHqK6rMTe42rpE/RwujeSa8S0R/yN6/7m/ApcntAdsJ1xE3at4KCreJMpiiX4ahiS1zysQLzuEg1
7zeBg7UZDlhoeI1VDwuxt4Y0VWxtARUOourtXA5pRsThZagFX8igM0+vIgwYuC/2RZ0rImfBApfP
4W3hNfb9aXSFYd2D6dgbZTUlgwIOzSpqQaMyA4BNShd/AVs2mdlrWbCe2DlCbcz+eLaLsS1yAzV6
JDgNUKqfZGjB9X61KcRXFzwNuiusiVqsQ2eq+3ynEaHNQggSLOxEYd6mzj82MS9vNq1pwouDLaon
wASJOZNC9WsxDjjP9QIlUsVmrxjHm1FkO1znARMpKbj9TISV3cYxMQuYYa9HlsAm2SmHag2SgwF5
Eb70cW7vSi3DZITlo8Hjp00I+8BjjjAQmpZyrW74FXzmUVGgAycogBpnu6UmUVEk3H0NqGFNrGRX
eeUGFZJrdXt7Mgtk29Aw+WjVF0a+kgpHLBZLI9RqDBFWaQ9XDRi+Wdky41QdZbXSs9lmpnzwNb3F
t8UZCZquz048qrNJfKXGgt61giiiKefFpTD7vf6QgFmMaM6L6GXK7TdXYFVFut4uvJHxvWx5DDee
uPN8EaIwKqNutQ2eH1F4cedD38jhKwkqqG1iESNMUZXBlOFtIgpZZWXOuJEs5XI5dx00f8iJV2Ja
zSulm9bO1GMiJYop8Ffy4kDO/il4QjmX6UWmxHiIUdNMCyn3M0FxBs8jOq4regPkIm8C37UEKwU4
WaxmvQ8dy2mZW2V2Ua6jWBQ0jLW+GMATzpwIYJ6KmHUmqrVHCG+bF9NxVZtf/8IUokZg5fVotRn9
IVTmqeFnU5CH0WDoUKVgs2rKZKKrBPvqFPrSERErdom4mr2NdEHIhNHeOUgqInV06/6bIYyZJg+T
QISQuwMFSFN2elJwZWWR/bHpH32xgxtLkDxcOxfQ22eo1K2s+dBPVf3VdZnKMDwQ2QF9P4vpH0br
0tF2dxLbYjH1WLLlh6/5AjSCRqf+8clk6dzD20cqnw9ONfexaiVIu6/k7G8ovOieJATNKlthM+Ox
2r+b4e8viP/Zy4fJqQ3/1nEzSjY4USDb36ZARXnebhRH4fAGd+9/nvWAyVUAAl6VcGgpEH3JtAIM
+oyJ+4CC54wa4CIiQGjVgriDK3Jl3uoh0+m7wTe9c4+bNMbSTKHXSJGNWL+k8RV5Xb8KBghSGJeW
Y+6BcCd4+pXMhCrn3nYHsKqjv3rmf8K/Tb5InaCBDrJjCMwI7yGMly2R34T7KJd1qCxypFusRa6B
HdXsFm7sWVSgpagNXsML8Vu0ZmykX8EkI82Qi95JGQNwneJjB6gpcZhBbmWFSlAqVeKEEGZDiKA7
PvgE7WnnX567ulAjj0+YuU9ooJ0K/kUHxqMyK2m2osK3PSuJTqKmhs1G94ALvVm0Q7qIgyh4s0Vq
NGBM7XaJWMNEMP8T0omfCsKM/rcqJPMQ8Bvd1tKiJY2oyzdwO0l2cLQ679TfGXvm+QffKGpc8pUf
SXD2uzJddwv5Ky6UFgsAYBjkzFqaFvLYbIwRHfZ2PV+qbbYS/Zag/pU/S73FtMWpUZJxpWEgZvvd
tiNd9guPRs0mP9XS4tzKgxvVA/DSVdAaIttFcTmmE3LicAYIgmdVFOggzLygy8ue2Mk7CIsaIBUO
pkXDU36X6fFZUZBapd7lOYiv9h6T5kfOFVCyEzXXBY7IsD6EaOyzgHWw8wu5oNQyssyerPiRMvfR
ilD0boEE0EQpE4DtnpygFM1OmQLAZaq45F8ThqWPY+EPukITW5kAuHOJuTvTKYZ090EaAb7oBGoK
74Y+zC1K84Ro5nZpnLE/zND5Tq335frjp5SDpcnb5bkwBxjkafxPrilNeFHKnXPrgKg5iMbEP4DV
/Weaf+q7DsMrBPjIKxuR7wVpNx7IZjpQJc/dYFgUqcAoGv2QZuhwwcJQ3AYYGCJYZEKtXqU4l4zk
JmD7fULGGuz18pEzRvh+XPIYXYfH3ClJpvfKG34bLObCiSxVNVjHsdU9TahN2kKcGMIeRxl8ZHk8
CCYuEZkkFOwxczIytx1me1omNeZPMnRKf8OCEaInA5eN8y7j4w5E7OCiaIiJfYOigprRWz9FrNVo
rcBA7/JACC6qbLkWdKi1eu7psQaxiOeLKWbGUJCYNTmAAhz54qxPbFj7LghexC1WiNqxLxRQWcq0
z3sbVDOHqYR9ybG2aU/To3KMYa6jPix9ZWnBF3VJO/sKXePVhFYeJngEtjSnNNm4pdOZr9HSWtkB
+fv4sQNjMSNxN5eGikCYIFeK3RllEcYgSz+LU9afbfUKtmWTplDApC06DKfiWh6WnvqXxx3L+arz
z+6YcI3lsdPUh+7uypCms1ly5303LXys8LQiQVO7yJSpfS4RQ6FFsSGyCAgxirng72NUkwC+e4XJ
Y5OcF0/stFcjvUfmsRl13EoDBgmoBXRoQxuPTySuGpw0xegnxq8Jc7fTZk9NW0VbX6FH5gbnyVm/
YbvlEhN+vSPg3LnwRGg01DFDvYz3vggsSYUsYrtLnGaJ6dHe9vHGrK71UX75/D0RE5dXNI95mabX
n/TpEKcOZQy+IAHLkIG9JoIQzmq3E3Hktiz/rqxM0Bf/zu105F0QnsDQ/YRewkvmPPqxj9RkRM8x
yIhHYJo8GxXkxTTtCGRENPeuRcmql6RfO6wbvSwtqd+2I1sxwziQr7L5f4fut6W/5vcmGWpRNzhd
6PchXTRMitel8knnx5kZJutVQlQTLhn6qhzoEkCSjQAAw3ixlrCNLHFvbyncw8tcDJs3iPuk09le
oHZsYa07vUAma6HybX9MIydvwtiio9bfSTupc1GCI0ysbYJgo/wMzei+o0IiPhC1tr7P+XT/59Fw
2lWv5Cv/XsvaKOMnhB09I1HXaVeqa8EZhQEQl9unkXxIJjGmcYqI23F+1M/tB7In63RBvoKiUx1Q
8k3KAx3+6GMD1FL7W53GvblDiXHSvtpP9KHkOK9+Z+T9CC82xtUguMv5uHnuuQmXn6FF7Zr3YTfh
z6O56FAbumSyEZM9NNSNwf+717Nb6joxj1w0YITGEmroZVmzw21vQWs9BW+t14xmm74//Qh8IlVU
J/x6Luq8EiZOoPl4VDzLWaxibJTm7ADwbmTgNdIOc/ixCkAP4HfMbMoC9kVoebpt4YgoeTXZwAE1
PoPLT6W056tGs0NNqbovyf2sK6YaTQR5fKGsr5WPr5BqpVOMXxoQhAB7WGJO1K6rf8gg53xia5IV
j3kO1ctQLwGsc+iwE9Qg9uiXe0NKI9p+y7bE18a8so4inUmi2a7Kt7Z9sqog8WgFjxTpBGQDc7R/
rnrySOvSsVWD0iLSAV9dSlX65Gza6RjWYCBWXS1ywgnE30kMpR/5xVDspniKtuSD2aL39Kk++HXn
h8PqDJ55ORQ1UTxriCV1u2YKZV3/BZjuL6mirFRzwmgYL4+Y5eTIVig58nOlEpwnv1e6n7hWoGFK
WN8vwpDqjpy/ASHvFglTyIFLPbRrI9Wp8qXbVgZpCWVnT7ZroF7L+keRnndr9hEs5kvHUyRGzIwS
QEYuOWMe0SZ4XnUicHyey88HwWa2j8dTx4iV0FBUJeWiwgsu7NKxq1J5nIDF5SpIsY4LRwIhrPRT
P/NR/0JsRLF2OasMlM2oTeVtRg3MMILZmtidKQDqfTXZMESafm0t+gplk9JWcgJiHNQ86wGMgmnE
uzHrDLnqb7uQCfFW6/UiIKwjzKmkFnOWCKENZ2GbZ+vUYUzdTsH8tDpflZdnu68APHsp0v1wJkff
7/jl0RV7i9k6yfpOO5fOSt0XeMw2eBf8TYLJ0WYdRijQyUMGeqQyltdZFAXap1uIXukLYlsb09os
1GdCY0a/1ZT0sQ4AmLpnJES3dQOSOR7O+/vINVGF1sFzONZH10NXsGF4fqdzRUXUwQb36Lfuqelo
PrOuuz3XAAJrF3UT93kgX7FtYH5TL/6pppeQFdzDgsnp7hh0ldLi1j1AwoQW3lP74Wcn+tndqm21
gcd9KrkA2g/YrBUfyVuOUCPS3YwPMiemrqsTpJSk1Ollrs+O1vFp+wJ8SLX/RDZds8QTDXG6wI35
qfIJf2qwpzd6+rjltD9UOcyAiKz7AojnbGESvkINumLOLIAPJUm7XVj6dzXroT8U6q3TVvt3nwNT
AnPaTOcAQSfSGKkCL+njRTYfFsfyj0k/DFxk8XITC+3LXnugSYDrL7u35iptluZxLX9lbDsAyKtg
pQFoPLaqa8mJuTXUITG1yGVjz4QKY9ms56jp2dKBEGhBDT8ffJMIjrUnLEZoM+6w5f1QyPhki6q8
C8EkDHwcTKy21/erJUM7dibFKcHczXLRgZAb3kiu2KJYxqn6QG40AXLPf1wDmCAAuEq8rctr2WyB
xUhFb1h/nsuext2UttWBmUaPcCztRyi5I99rA78hCJrUzEufpNg6qlGhD4GRwFcV+2rBAq1lN2nF
uEzNpSTLpniStumZoXZJ5UuBt7mYn83mOykMN7AxiCBeyZgmWhz1f32z/khGp1dkCfFgIcgB35O6
GqLKeVxK4IisTuxiMgq8goheYbo8uEKNqG7bIg1tt959CNrRRDi/E9ijSam72kgRJplvzsubNjlx
ADhAppZ3kbVsCpCvFu6Tr14XU6c9WWZX16MHwR01qdLddcnJhodT7dpok1wGeS6fM1eKrLVgUtJg
owId9f9NsFu6T+is/hhGyMdmSS9Y/vs7zn5h+tQYVMiVNeaMXnMUCG+PnjoetUETEhyCpGVzlJas
q83onQzqCp24ZbWADl03o50SiMdKIT0K43mwjsDyCrLgh3p11YCGwhv2Bin0ZQDjokM2CkdXavIs
hKSx8dV9ZQIWFYCxLW6lTRgfrNtErDyp98I41+fht6Toh2/avnqXaMteY85VFVsn8h2dZCRM0Phi
EHvaU0ovRSXU3kvWu8UB8gxbNv7LFUyZBuvHQ1wFDP91UaABaLZfYiRstlRtD4Q/Ok2vItybR0+2
jyozAcuwpLYRDYJus0Ry1J/dPzCOM0fI2oA4ciPNzCB85VbsQ/n5Xc1v/VJKbKwWxFUjRzzX0kSv
ntPXEHYercFjlqGDahBvdkIHguNBjtsPNVCMTLIttwmGUKdANurbMRXjrJ5GVML0lSQ6ZLpnFnhq
2tjCuy+425wpc+4YL2eGF9wu/CQ70S2/YF8nLKSxRCUzn8b+p/YeHJcW5mMG8eUVXX9Gg8hV4ARm
CB0xbo0tKMZhrNjV05bj7/IlKNXaTje6XsK2t/2PcA9xwYgLukP0v4F3HM/vw33ZkPHKsKawrnpD
E0kAxrXf/4PERiYeEBNu7AKp1WBO/gmqSH4qL1ZqRqYqUMx4ioJlhmlnmD4H9BMc2940r6wVTkW1
KXClMNa0+iNLHnzdlwTn1Kyn12xCUY7BsA+SK06bKLmu1wryav4B2CpF6mGF8BuhoM5aWp1K1Yqx
EFs1KkLEaWQuMAwIhKoUTKA0wM5boeD3aFGDPRAQSA3OlYJ1MuqMEkRRqj/U0erX/gaO/tVROdja
SqKE5MvAH6QtO1Ms6EBx3lu79ar80VrMSVrs718jEmZnafX1sb6l7z/eZwYUZcm5kr8jp0XoneEA
YtU0nZJZzA/qequpCBrhbtHAU13ZuxrndxlO16Nx0S7Hxc/WhgESu/1rqf1cj/3BkYIs+8OYmWW+
YZPVrQdXiGLTHKMPem/TVzhcPi/6DKw5mX+1Fa/3eCxD80DhC6Ii3H1g6RO+nxNO5yH4IiUcLqfP
rv2rPUFX+h2FHYKxigym2Zvv7Wpto1J1c6dpqfZHaHWOzhYDqIn9d7t0iiId3oNQ8Ecfogay3wwB
OKxvbgSf0rgQTyKNBQ5SkelAAYsSvUc6XoaML12Wy5iRR+u2apGMYNFH/4KrMnIMIySBqn78YTbr
RmUX/utVBA278oIsU0B4Wzffrpof/CKuDe6q6oLjGDTCQGs4MkFAgEOkqSkSNIkCH4b/Ay4AT4rN
iHpH3X54q/dS6PE1L5LENWisd8JuoFlKAD+LwCqdd4gKjji0lrByG5Y3JVjd0qJzEKkkqUYlRI9f
AKTz1hwIwLICZhqHd1MTUOg7PiE3gzCHJzZmh8Mi7Fj8p65vkwAZmR3GS3ofDqfyaFn/lPJeuSpM
5BaYUkXpEfDYVI0IIm1sozZq7hEprBcWCnDzvS+1iLfpNGd2TSGvFwpTNpuPhxqd5P1xXGScoNmN
p/L0M/mnSC4L5NfFG8hXn2qgZFo+tQGSd4101EQiMr7l4GRQEZGDfW7XlJn6yUoCRUBD+ZShnwO0
aK+5eXcMPBwLFyjrgItIdoLlkgLrRrR1vb0gGynNaJ0oTNRi3jdLoNZZnJlaeFvWy1kEkppiHcHK
TlgrXM9TT8EvFlfNw3v0snuXYDGdjlkoYVpZ1KLjBruPd6mBgudIylwTsolCUwpf8lMTSXFuf+in
H4L2H7UejE6nNpcW6lvy0Xq+sn/OafujsEtg4v7NcdRTm7W3lXPcTBIuqOZgGncLocUkYABmjjDI
tOnUiMcDtTsIDbJDOR6e0BfEmNneh+qi1Kkz7PzmSTP9ak0bcMFWeWxdLi9fGXkO2TehU/rfkwuo
62s16RBfEeuSSx5IILWViaaE2Yut7nQowRw/IzFqTU8/9dM6rLjkrzANlDeACYUiQeHlVVQOoMkv
0UqxYdciDkuCAbnxEOS1x+oPxzE+SXd3/HLaJ6BaPqNml2MncQr61nkEGsvoFGDyi5F9B7tPDayc
lppenD6cv9BJSUBqbuN8rAlItUPCzWoP9b5IUgl1U2ghUE7ez0Ba4nkXDxzHezNsOYqyWGHuJxk6
Tv6frbuTJ4PzYb34TrEZe/D5BdWHRyx65i05THJ2JzgEvMzEjYFBsISXzk4gMXY0vJpbgzSZNEOu
w/qx+vXQJGdISuYKDC0sQk1mMW4Ha6K56u9SRBvsn+EU12JG/DwdhdKKmdcdVItGFW/WoquWbaM6
Y75s+FtJLOC0t0EA2xVaw6C8bk3vvMDgnR2XIAj1ZSxbUY17lq/IU07N8NqYIoNk00SIrIXNCGpv
AWeFmlv6ogyxhPurWw2nKN4inbeWiMYPEM60zKMSr2mcP0cYUdXMH2FpA4XCXuSZw1Rz6/ABLNou
eGaaLP53Zfdh5P6o36TW3Wwu/V0YihPRxWMPBqOGbEO2epK7GpnNOMa/q8dJgFliJxyJ56k3AsSu
c0GqWW/mu+mhENGKAFYoBHyzzbkmmdyOfLGuO9AbbHMBwxfAIOwR8KojQMrgI6zyyqgkVuXqIPDb
2+39/JLtv1yOXfFjjy4ayzf2ZLU7IWdhbO1JQPUFjoZn5GBfBHA6eGfuewElm+4mfDdEx5oES+R3
CUQrcPQtHNMY3tLOyvJQO+9Zka1u7ZJ/Gbh59YJzzHjPRmfmoZpcjTwvuaY+vzbvNATvfbR590Kg
LiqT7P6VB7UZdviVm96zf+q/jxraoHWOV7fxXmnFS/rP2pvoStUCCMzFvAKhIxZXrhjj0YDP4/Q0
sef2HMHj3cuJBhk+H3Voz0wK2whnc9SfE36AkWCfcY1x9Vk9CHqmtgRiwWXyrqViGnCBesSHFaJV
5ErUNNpayqEMv+CGKqZJ3z2+RDc8db/tCuGU5sFUL6ctwIXdalsxWc2jMep1Wc8Ip2GeDzvpiCMp
r5GcriUKRhEN4Ro1z7fbw3op55zgcjSus0Emn0skfMezBwf07Ki/qWK1EEDFyOa4lkbXI+vrysPr
3J3oJ8PfU6iC8n6dVOEvueofErMzGNphtZVzgvD1veX2d2GEFeQ5UPOF24lugoWlCaRT5nx4YIRp
Fmt8SX75bvQ8GT1hvw4ZcIAEfIMLIMVT2cfntXIogSyv85QtD1++vWen1sGUS2oJ4m/wkMV0P09i
Wzg2BKM0ghH8+LTHpKqIhsM0RPs26TGmgLSmmH72DYg25I3qkurc+7SEjb5CyQsx7dwO9FKDwFKE
4VpbDcYT5zz+n57L45kRK6rNpRySOmYHEpBDsHPwJ722AtDfTtQh5RO3IVeXwSJs9SMVAScMefQI
VAb8zpywfsW6TsTYuf5E1sr2vyVv8fRvAwm1xtmnpFDjVhu3WIfbOsnO0nbNNNMPziXDyuOaPfOu
0Cck4dm8aySWrgGSAqZgt8t38j17sVDP1qLZnsRQpDac+IA30hSpwZxES6lBM448vzr8TkVvRd7Y
Zr40tJtssNvS72beNxlDSsixlcCA8j1IBNXQS++vZLb63SYt0Wl1I0voHbsIQIXxsKpEMeVq6XX8
33Z7fnqRpBt2qXg7w0bLK3Dke3tLekGY4LcWcxrMP1/2Id29UHkjNdXEE2k4IWa7JuPNt6Nu8w7P
xM1tmj1Guv3pEVC6s9Z78hInZCth7Mno75WjMWkZzN7mt+H+uo41TffDqvipuUZQymuEYA6fpdlJ
umFKeJzfars8oM9QjXE5oBCyvhqRg8d0wW3d0wzqFHYm3+GFOJjYEgrWbf2tunrrZXn04mdNBsun
iPbWFYnxeGErTbSBZBLnGkWALCqWhlzlvqquy127Am9qPvcdenQ9wJmi8JlMB3sOJIgMLe+KoPtr
CkjS8Nt+Bt3MXmWjcdEna5HWID2UaSNpeNAS0JY2R5RPvdp93QFxVzvn75E73YmuXHixFmxPp3vA
NMgfT6GFYLVktKvJlDa5n6KuA/uZoZkiKXkPPFyZtNVRNdsrCmqSFWmX7iAJlhjH1zifCPQ1ww5C
3F6YE9kPdQsEyVyQkJUWr/bZVi5yj0GoUjStKjTN3ZXaTzx/7qjk9uVePaFedYPqPC1gKTV3GpeD
jE5X7mjp/u/gfryv08GnoQm3fAHAjo4mk0k6GxeSbhX7SAmg2AGWfvasws8X0ZO4DSkFfrg/WmRn
s7MqZ50YIOq9W3C7vL2YJ3xpkSJNm8LjVxbWh49IXtLUJSAFvv/cY2BHMB9udAotcw/ZVByf/5Z3
2bpI8JeR+AO6p/HRBIRM9OLm7ZqWj50faG1MkvSPtVuWVd2W3YfNToJUaOFTu09Rc0HCB1GR6Xfs
pdzBjn5/NMNzhlYpUEnsYosFnijcGnKJxUhtfA2HwAX9P9hJgqd3qPtsgEV0H1OHHA6IHKKNQnAL
AFPN0sy4gNEF362TaSCNfzB++seJgn6+S1CYRbvZ1YsgqFnOY7gFGsnJsAP6gSRzEXPoja3GiMri
GNm7z2ZJOF3dBWidE09VPiTHbrYgvJRCwxKZU9SJ+WWbDyO6CANNl9uXCsC0rmEBGmhQyy1bQJcs
jNWscHwGqL3b2Sqnx7D0e2Cmt0Rfb9gX46n+gASUHajl42nF8WFKCdrM4wLdej7puWXL1gAHOSA9
a3RORhlr69xkPHD1dyTDYDpmEB9/70DAPBmBpJyuOnCGyQz7/dBeIlLy1VIe8W5cp2e62hGXCuCe
pKXZIoWNbYmb+AVdJX8VoISacxX3F5RSjIngclJg7CVbDjZxq7g9+DPBmeBZMmkGlDBBMTGjUsEE
0x7Hbn2NxFs0dZQG4/mdTl8+DL2qAhPqZ5HcB4Ci9N9S1fAQgjbmUbRQUC7plTgkvrjMX4AqsMjV
Gf04mSEvOCSblCbYeavvFlzKKwT5eLs6IVyFc9dzdu34Ffxzvy2dj6E8ZI1KI+NOXV33OsSnMTkI
A+feVJx1wW0BlcGXtVWC2WmiLbJGIC/gRD23iUKb2/mXvlHQCpWuY+8f+fu/jdIuxTxHDENQ6+9r
2uK8mtyjx/IKpm6I1ARFp3XySb9ZhoKODyMxTXXsyFxRrzcAkbwm59wQJfVjBI8oeT7MOX8+bS3M
MHK5Ys6kuu2b6j8UQJTkuzZC/QjSiGed8nwP0jnvtL+3in2sFrbUPS9Lm441zvlY7L6KW5YE9LRu
ikxmEzPtR4VLQ0ai2yov0hZ4GMXti/3ajtshAku5wJDhpEm9J6vTuKRbcWBjmkeMwvOIGcXDj/ba
9Rs74MmnGmkE4ysfTYTu05fy1+fSb0LfJGd7ESa9XOxrV3yWHoIuKbu4tw6MOEc1Z9r/S3nznLXG
ZjDywSzw+jMqg9USc6B8SLOBSJ5rqmJUK7KcW8lnt9tyMVkHOmSuCmOA4ul9A9e3ML9fZXqohjxB
0o5ngMQJ1yuCP9/PyPLug10hZBNxfV5Y5cTJFjPACaZxHskhcff7+JPtifKqeBnLln38zWFAqxbG
uKp6iCNmgkfvo7hhNv4Mc6tkqJKAChoTV9Nu2P+UZAaPrq1mqdP3gVvg3/zGD9GhFZs6ce9f53pm
sMfTjCVuFH672g+NmXklbiwNvPbKEE4rmYtQVvwRr3XYctAdBtyB0ACUK8rqgYJIY06TsULg6biv
902iMg9NOlWt4w2BkdXr/u5GwA3x42s9B798YtVAar641GolYft26JYY3nhbNGPOLoCjeTZfmtLT
qmrKHVgOyBuoRKmowA3SLvLBEBoeWWm8PkM+6uIK5D8dWnNwOb6+Lr3CCgFTbw2wUkzAF4w9vjre
0ovD7ucQG5ql6Y/V6x/yonDPZS+4ayXvZtP/2W3ASFEDE8QFmrZBT9TbAxSAfznW9K5vxyDdQlKn
BrBIsCD08Zd/KOr5o02kc0wM08ZsUNDhQf3euOI+v3kjAW+sd7OpC5XuZWbSOElL9tjU8NDoM/Nb
1Npx9t62ZVbXKuporIrFpw2f6IbOvtqZSdZcgegEXEQxRc8A7uKTMlwimGunvXMoncWSqb3P8oTY
p5OdPgb52FPlvOFv9Qr1bQS7PQO8A9KzaC9M3SF5mNgzdWSe2LHaRjOZelSgl/SJZxvvfnxa1v2E
K3NmJtd/WX9CfxFfC6AsEdy//Aj1leRi00Nu+7u1IweA7UXnct1cF17Dw+SpxXCpcrQteNoeSx1n
sg3qE/HKbGpknQdb4HJVdAFaps2DTrdw8V3a07+j1RvmmmWylVtas18tAcApn6tsSbcn844J5QYV
2VkND6n/JX6bUmhesXWUsr2otZDF46mwVnkMknW6nedfwnXWpjHqe3qY0svZCylG1rICtzkAh5oC
WuNYeoufUvZA22yiHAfBSXJ2GpZaj1HmmX+zj/5bhI48l3sIG4KIOwLFjD/StQDT9c9eKTWj8Q8s
hutgXme6ayxaqvodd1u2kI6s4w/oWFXdA49itrLcM05owOTEwkyknKygCWPibox7pTCiZCcq5bua
F5mUMQoPPDYxXXALxu8V/h+F3vADi1MznQvdb6vj5rR5AZNjlB3+RbgGf8+u6hwObtuKWxcvdNQM
p8B2ZFIkGjlXe6K5xz+HmXefzO/dsYokEy+6t5Xm8hxVhi7BGNE3GI/KC8kjhzl0Gmqx9xZJ9nqt
r9wRKsUaBwGlIZorOULPqjSizhfSW+tcbwBSjjerAa7HF9dUKtfXdW0oV6Og68rmPIUlhtDUS6jq
t+zkgw36APa663WH6GpbJx8mEAxte/NYy0qKzl9jjU50Jh6/dmWGelLw32dJ9SRVhKeEogu6PM7C
o3L2AbxVzNZWc6c8XQ/CSp7+EODt+GBg2ZCv271yb3S3s0LhE0UYVokWhRb7VBYfKMdyUL4ySFBm
6oTG119SsMGcjVbKDkhYnzb7VDi6pRbpRcQA4q5M90iMLoAyhjvqcg8A+GicrfdfnDMe8jFQEFxG
SoOXk2tl2puP+5srZVS8fJr2Gzn+1fjQbIU0U/AN6RgpjtNxCGkrxCfnFhvIgWrnzrTG0XNgkZ6I
lPzYlMWZsWn27NYAhE758N1jpUe6ZyZ/doI3k9AC91Zw4ZxuQj+0LlQ+8a/S+KXBJ4h904EfGnW3
nvwtO7ZVsokVEJR9gdwouZ5UVysMrRhU32X2j3biR8JfkQ/ir4JRd8DQfOcPAjizJVVTi6Y4Hey0
tRkt1aDMxLAXxi83nsGFt1UvXjtiHEwZykOzvpShk6+zBDS1n5IUPbwjx/+Ymb80BIaWtKDGuTpi
eT97+exJGdWRzzBvNqft5IigNVg/AAYCZHxg0m8eZf4y58PgpN8xvrT9+za/HICiT8gH4DR0f2pd
lHkoIcj+qzYp+yvgSIUtDw+iV7m0i1HTH9AOrsr+WKe2l7uPWNHdueslCO+ARYU0TOf4p+j2G4N3
2zf/u/LvssukBAx8q9os6hFTRNmDzahI3qnR7J9JzNPy+gs98Vd68SDCOF1tUPCh84Q1lFZO3Iwz
zl+YaUXrbGEb8WqiZWhhxQOKeU4T/L8P48hADe4qp7r/NigyPuPfCSQwHGUhf0yIMQmdi5WYeH9X
wYaXkIOk3HQbIf30bWjNGjL4dh0IUCU6V7bkFj4/JMdsBpKz0CtxJ5dAhtlvxmCWOv+dVJazVVrK
IAPoZi1/LJc2g9cE3IATsaMs8YApcgZjk5uzxh5th7hK6r+Rm22SuUu0dufxbdUeVKykcRB+k6lc
SdSSUMwbgew1c/GVS4d+KkiRbhyd9ROOweuSHw/dqIUKK0+5Fvf2jAaKQi8S0mlCekCWtqaZYzB0
Gyof8GlmaUZUaY5lTkM6Ac72LF++5ZY3km2N2Hxy8xwbuoXodZ7BLJ4GmlDg3b3haELhlPOfuxrF
TOgu8P7DManoAhvRpC06wimQiZhL50tDQmq0QpNdhFQo69IGzgrTtlm1XkdwxLFr/DP5Gt3598UL
aqxkjWaOCs3RIhkuPESbK80W/8AXRt5JavMnOpnVuTV16qBN2MaXsf4vFihX2pCZPkGmZyv3efke
wC0S+H310KmNqRNlidFugpvRlyvX4CZnRw3rJ60zxX/tI4XDOlVyBHqkuMIPO7mZuM0wRgsOj4ur
dzgkdRvTf6+ZcA3UrescIvkHbxGGQvpWWAAZanyf9RaXye6x1mWLUu4XuCacbquRrGxzn1XMRWUM
MSrrPv+DmqeP0rOpdtCz7Gy0sgUrLsYWDeXrOAt9y0zuNJQQMktt72I6la4y4rYfksFRPyxKj6em
yEWPn7miPEsYZRpz2HcFWRAoQLiLiExOg67S88vfFYCjTJVp/zLYfwyKh11bm26udTw/jr634NN4
t7hbSVvQDe1JyV1jINb7Q8ETmbWlWdjZxG97mJ2scMaDsonu+EgjVk8OIvEYcQEkD1Hb8a/TRR1l
yE5r5JGt6IgKcI0frDTRJcoKBGl+rvqMx6lWG51xJ9svFg6OGmBS+/xnLYytCtPCb2Rs9En4bsnZ
7xLGY9Hi7ddXjKd85oB5MyvT14hYU6xxO+HFp421pindIoW/+4rQHr5DmX+S5Gj03BZ3aGSmdpc6
+TAg/QQncMPdDpMh5CNAdCtjELpE4A/powJhFStzL4kNKRj8SENJ0X0rbNv5HVwlTylpxtPP6I2s
+53YZE8wPSUN3Jw0AyWojmlhDDuyVDytohAI0Yk/mjRoPWD4r6MJbBa2NArOg/uDPrFAdtI5co2d
pOF3PsaQ1Sr9PVYtIbRkBKFmXZUhT/Gdl2JS9qQJC4g3Cc8W9m9XZymu3MXOcIDmOzSwJWrNtbh6
U3AWerqAtpOCdHhhIt+ShetrcOdgKtl43B45D13jc3Nt3FjrJ5KRxd6uL8czhz18ycn3zyZoi6O9
TDlW3BgFXivlpUvNsgTtxcQVxvND+Zkgw4kyIZeYanxNu0wGfTUHZNXi86mfz1Q8P3QkjO9uzsaa
8XoeM0NTqKc+ahieF4Uzfll/6rcMUww+2l+wQsbXUgMwPxo8BcFQU6XOyJOYhStbtwLT8RXSW7FE
KRlbL/bixrU9Mx9BkqNTmfLW8njnq8AIcNaxUOi2SUiarLPS81M32KPo02+/ccfhKrV2Ym6VQzKe
7aDVj7KH4OY1IhspEmoKRBFhYWshRDjTbYjUxbj9UthEEBGQEMPiuMhU7UsHO15DQBbIuk+QWQCr
oyc23G84IMjx+FxkSd2JEqCsfqstQxhpvTmcAcsymZQXNCJFs+INGSLxcZufBWKMYunZTrozoE4R
Gp1It30Ou7PDi8iPMinnEHCbCXsCw1WPv1y3iwO/JU69/Sj3DNQgg0HVq+WlhODkt2AbPKitWc9d
//XPWmX8ICxkY6jOAbCB1gwMm9fM/GHcRltFlsp0Q3q8N7NAJiEG8NNkvFlOUPtVL8drBD7SEhxu
R2BRAaMStProYg+UPW6GLi3dtWNP2AvMwmLRw4fs1uOi7gJfj039KJfVFNiRMyu5l3oZX3ezznR/
9HF2YFfZerLuZI52ZeQXrm6wNCVPtjokmnw2pxxDUm2yJbujcI17CV4hF/fDSAnnUSQ+uvRfFBf0
JlHUR1seQx5THWgiaCZXGojTdTkl0gp7ZSme3FZxRkM4LAvEeXQLWAVPNzMGZq4T+kZwbDJDHYXM
5JJCGEb/DQToV2mRKDB04d1BY6R2t5e5/i6vuZAEkGZQ/M4XrqddshDV4bUg5dYWk2dxiSK6+Wxs
SZp4u2iyBHZv6l5hbmknztkmdDECdoXAFwVrggWk3lveV845c1k3lPtiu3fZ9PoBA3XSkRSFNkom
bR/mjP3zFNMy73Upp9fBGTrCaB0OR0dzBS1jhWIy1RfhhkUIPFZewHSBhH4u1AMpjREb6P0B4ntM
yzqN+sSgjQFolxVRAvBiTYGq+vWRaYPqzTtgmZmsQXyigntQfvzA8cwPrzvygk7/EjVG+yJQB4Rs
85P7TxGACJU/0D62icEXDj8mud//BHSuhmj1ojNV1XyW4q65iL5CITSFlBmGnkDEBUara4Rur/3p
BCfcKSYq8ZCVb4irb+IRHmcGtN1rLP1vRbi8MGw5Az3HoxSKKn7iebEWhQgCNq48Sy3AMEhY+pLs
Wk4lvzSM2hZaTRsmKMMpyO3Slkth0ioZaPyNjl7xA1OJrFPtojK85WmLJW24sBASqnqVr41ge5mh
L9+vYWnR0frNVJi8JP6pJApMQLp4+HlXPgCrcIrIUedF93HwiTJ2SPVJCbq/Xv1gqMMc1jh/nVZh
v4LCvZqycU+UTm17toNOzBvUxonVEawSN8GXEOsZdQijzwAPTaHVYVUudd8hbPbZS3D2UFxsXl4L
d0IGs6Xn8vBdct53IgPN7cNJx1OUk1TuYkVr3UV304ZjE+b0h0HdjoUPCxbKCzC7vhMsfTDtXnyW
xqZ1WhPixeObQp4UQsXzUfywcC74abwF+1+CmsBvX699HqJZH6+4Y1vmsNTZ+EOATvRrSvW7Cu95
jyv79ZivmN+iEt9orbcOjcJKmZlRObvxfGjkFP6Dsgod9U9WN30dO+fC4LCBZHEYb831G/fCHMy0
KDLabH1obEXI5zJpcLBEmSj2xwCjManZSCrFf+GQWNRdYExbbg44vlP2hw5ayYNW/1EB6hCy+fxG
qI6CUSVuY8oocWDqICnQOJRsSMxX+2w9mLKC+0SHURNeAGoEDHmV9hScRRjjnj19UU1FAcvPxE2w
LESOLBhJStplsvlgbQ/VKQL7Ijydi3X9qCtQZBj07IX3tjKAl8vH90BdUR73Zc33ioZy61JfRhVB
CLbjMboF1p62zevAkgWFVEhSg0lXuw0D91780WI5Mgsu/ZfffxyeIkxKklhIFAGASz1Y+mjiNqh0
KFzhrBBy0lc6dgqNacziIaFNYJudCEmRB21+101tvOEvljKbdTVsRQCHdaKZjgzWo5oOJxrdXnAR
DLPytpoSXKYoUmCHZs5RWVVkLb2BsOt7/ETYuhj+CynGhKC2MS5rPpl0szyQpR6GKaJSGaBIEdcy
0pMa41Vm4IksWxwMqn7bAHgAi+Glmuo4AQbAQzylWgNGxlfkltvkHfvelHKFe7uqqJhcuVERlghT
4Svewxg5D7/4aeJ+I//DKCUIgRBHzgu2o1g16SNRIaHuOEtkvJV4KjX9EeDqPcrJnqDVPhzKdXOU
ipPCMn6oMW2pQFe+e2s8yKJrSNaPyQF75EeZAFJ3OPWup1aW243AxeaGXyM40RMzIBDiHcxkx2Fk
CrbAAHG5hQykEQNVBH935R+/vnQ+OwA3ltkgy2hBCqKTW1WwpPc+Q9YjamZsxRoHoq4MwqtdiuoZ
664WOdmMis9gVtbMjX1yAqMgGdoL9laAbs2QoeeEcoAT9R18f0YBZsC2Ro1TtQfkF6K4ZGZ/CCJh
PnvbTof/VydLlqFtsYG6Gfq0pD/K/ROTY7edLC7ieStPeyHVaiAyfmHb623Xy8AUDGgHH/fduC8k
b7Titbnx3Q89iDjEtML6IG72M+VNYCjpDf1Za1p2juF2/qAKNmRcA2HFS+wR0J6P/kqUFPgRhtC+
5fXYj6Z96WKo/CK9wj8zz//6Qln0Ctyg9HLILtFYeKiv+KhHwm17xgdmJA6yqExm1fhilxaWbbtb
X1QYlyydGaqR+3ZRqpJpR8PAc/1nbevKT9fyZsf4/Igjz+IqU+aZEbyndDIlkOMXpgold1l5+xQC
BGDXo+pzWl5jqSbwkmEBtUDWDAfoOHHdqdBz2FJJdiq21EAiOF8pcBNQ681OR2yqnTwKEwU/ErXM
mnmLMGLTiTdJWiPLCDc5xo6p1diRWYfipTiMIDqUsBU7YHT4Zs/d7yxBBE8sNgwlbgQvKKX475xx
+6YIwk3ngZUNKDoflUcjGK8zG527BIqo8uS5aljFzZ3MG3EoP9/Z/cQ05KZia71fdIprbRpBfJgm
t/dI7Gj0nS4qniDDDFnz8X89FMyZI09B9+PQD9+D4JFwye+m83t5dhsoP5u1+S8Lawi893TOo81i
Kb02CMkrqcRvXtm02ijJUtNYaeG0aWhbd1fDF7OcNzNVej3ZJQnlIXyWpf+prsDQnL2anl3vcC09
VKYwCVXJaPtDMRHwrVfGeV9A1RVIookoPuTVkRAF0PZJyFX+ANfTTTC7t5OmeTu+Ep188N9DEAUm
P5TjHkNHLLMWD688R6o7eCwAhiYBnC6d4U2DBwRzMJ8ky4CDPHRBtviDXAG7dKe3BcPs4BlPR1iG
+ChA0Myzm5G7kJ6XZ1u5UZ4xaflEpy5I7herDKISBTPG/k+J8SeGFB0sXrjyQP+jNbl+bSASv4jh
kGomkHwsE2+RT+RNI8c9zf6BEaIrm5uQT2xOGRi1Gi4YfkoGa8+j6/h4BGB3SO9ODa0iz0chyAH5
vqeHr7eqqpJ5nSuyGOFoQ01z/ALUwh5b1Zhmg/5CT2WYK+83W3kTyS0jjSp3+UlfdQTnqCqVDVIG
khpW9imByGbXnofIuBtXkbcwnNKKK3IxgNGPQXtuI6r/e1HAKc+uG0VpGZzCl3Z/R+UiWiGQI4b7
iFcfkkp18l83OzavEN7pLgTFCTb3/+racRF7HJu/laBWI1TjltWo0wnAQmmMWkgYhLUvIeXUHqQx
vdf0W+A7zCWyTXA34C5pTzki7KxzsuTzFBBevUtn+qt1yJbB6beopJ5x2NpGIJDhlSEDMOwNfsfv
q+89sY13gO+MnWsueIHhcZy6kxY2ufevfRnB46NjdM6XpN4dwLX+mD9yc3jAz4omIpM5RZMGbY7g
z5BmgiHMXzRBl607fH1RGGvi9Idf4GbDzcbdckBco5805Q+gl1o4TNoKlYRn3lgk8CVaf+TQGOvh
k7mK6cyl5+ADrs2ps1Mdzo7j+vKWFlkcaqj+bIB4Tcp9PKjCKoWXcwjg1LKO3zKW0Mau2BM68KZu
rb+jULkhrP+uWprpTs6iJ1l/FRxdZ7MqPbjpEplNxr6kbH+788shKjVU4RgmVb0FyG3UHs1G+ksP
JeKyKumLcc2B2oZFt/bkrGIF13eTxj6PsJSMdyAwrT8yX589hYRcJNeepgZlSiSp/7m0lKGabcuv
bdlnCpu2jUB0U/noYyX69VMHY7d5IiMBzhJfRHolYwJ2Q0YJnecFriv1a25sNzvFbu7x/Z7tVVVV
IqYl0nONaDOwQTXgTGWhp0FT1i8qUdX8pY5kN+at4EIaYMzrxXRU1uAl3StOXXDPB4QheIGAukmw
WeCJua0Xsi1faSur97ZlH38/FHInS3wU9iUzzkagpUHq8q8WR81bkrUAiEP7upUZLRuMvZmI67zK
xlUDUvInmpwzFgtKxH0ovv6JMxNkeBB7zQkN3FbvKfOpnLHwQyuPUxOs87Ppkz3jPWGzWFn59cnJ
FXvhhW3eHvOAU5uKhX8Eh8voHVS0KEXFA6F1O7k7WvyS4YwJ9oRSie3UTh/EkBFuZV/CHYmouhPI
kxBIARCN0eWJ0o5HakJTM/QzCvmgbqXR34fTJwGQUp6DRURy1Ci8I7k6RUGqLV8xkDJIpafToPoK
44kz02Xcy/gshai/YWzfS+l6diBjI4TKN6odGtIrJFMD9dpMrDVqYZmT5CxlkM2zdE3s9fChKnkc
eH8Von8ia939WoRKTF8Er+KJS+skow1k7Rr/ERQ4FAKS0TBqTHhysidqTAWy9RYHgiQb7bCkbTyF
N+ah6yUK7D6WtMBxNkPufwTDMorZaShcRL/KxmVGyf8orTsMKwgKH2tbbxz5KySHmqM61jJc4st2
9hY8MVhaBgoy+WPMahErvcUg5FwmeQIVXRnFvJcMhNqfx1Wwgq656egfOrvMNMXAwYJlInjJKcdb
LvKPTmcf2gtgOZgEqKI38XqksegPWCroAg0iwTVkFgyjyu7/laPef3jeiHQwAZ2EN16vk+yiAuqB
gRnpB86FEfxrPSYfjvHHOj2//cCUDGnfX7XqfJJeOFrjTtYVcuosJfX01XMxafCqZPgZ4HAOH5Op
HCxUg9Eho/SW+IqAOhiKXLgJCYfMhLVZ+FsagYa9NcZUq4ltYYhr6TYGADzpHsL1MMZ4lp2pdHs2
82CR7oUlej5TNDbAyZEPrdQkcPW4lzFfwb0zAh19asbhrXrjasb47JUA4TF25cwUBKXYv4Z9v00N
hWO0B1pjVOi3YIX35Hbg7l3Uto4XM4r6urxxubgFz3L6LR//0YanT83yz+jGp05A+Q4V+8zbyP4Z
B2B7/7GGfnQEDXJf6XC0y3LSVw7n6EpKN12PekJtAYY9adKfcEISeHpsFpGQwP5lADGlHf9Gm7gK
7Ge9wad4QU8McO2enM9I68fNIKLCKm5V3Qa1QGEUMgwhXJypdgSwlTwuuw9Tr4ui6RdHGyJqFhRt
E316CWly6+jFf0BAFt0tf0kBb+muarj7VRGoWZlN0cyBI6WecRW0Qp/MYGiUvdfgrq51tU/DQC2X
QE8W+ksdOLA/Jc40UUZHR7wbPgW3ri9r2qdZ4YvhFUCdG5Nr8ABLp6GDhU/f8EGSmgm376992fG+
qB8AqlaPR2eEEvHCO2CsE+2IvKRWM+66nLAbyz8PO4zfeZ2S1qBTTASDUs23xuVcR5lgHitDkUKl
5hEKH+cJqMh3EigJW0bxwAGQqW6gxKMjzitivvH6MKA26yNUcAFXO7+pMo4B2MelQepO8VHKQgqD
BrrDWpmnHEPKjGKBbyxB42s1g0QSYPi5Wt7wAQCYR7feb2Tf3LnIcOs9HCBcMvN1etY58wObBQuK
h0/X7j3tjAqBpysFwOPs6SGkOpzG6msV760L6VqOXj/lvdVUEJdDI7hjYxW6UOka6hjXwfUkcxkN
prmitj2SgaACMLjkreFzYN1qmFGBefP6LqvNbIsymKXkQZLQLneQm+EEO2KccqdnTZfei2s38Qhv
ma5p4WFD7D7l58qEyPV8Z3nwT7rPYO6kJBpaN+i6s/WqK5Dsrrv9Dm62tz79Llqwc54RNjkZRJ6Y
GvbEt7O5g7nT4xhwuWcNQejJu7HBa4dXlaf5T9/BrwCVETcNWhj/mO1pK8a0M8Uo1kyHFvyjw2ZI
vNWWLbZBQEIcqvNVcx+t2+/uvL8Dau1aRS2CQAChXs6qeiYU+bbDQeg6P8m8EEpKBG74oVESlOra
dP603C+E02tajv6ui8/HexOrFypoWSGvd2OmD39nx2E5vl6YCTtecirSLTrvYCsAyrNl6yPoTSjb
5ysbbpU2cQe1mpsVGkmpmGlKZ+j1h3dgoVl1t6g7IJFg2LLrCtpTiVsJyhhPW8fsJNoRGmBrwCZO
XDknQTgrola4aEh70t3+zYscZIuqhyXxqEs6p8mGzYvnUE8DE/3Mk7dR205+l9BMunwEReahvJTC
E/UCYCQFLjTIV0HHT5+mz1TJUJvyV4x3ARe9fxckAEhkw8b9mccvTmqEHOd53wNnxMRhcXJgSs2n
oHHgfD36sR17ZWm9/3DDwAlm5f9puQJflwTOrZ782eA7TxFkGnI/Q/pCY68KKVazzLZhCLiGG0pI
vqC+4EFCSNcEzH4OqhdbRLj1izl7UxRq9XADKngWbuC6LLhUmcxuDHmmz1ZMV3nl7a3jJqzxLv3g
fj4kXQdr/Ldd/4Mv/nOYFG63G7OKt/qiYNbwhpj9CAL8mADXw7lYNoPYBo4zvTcxQbwokItIVx0h
hp27ua/abl8S0NoBiHlosfz/ampMwpq0Y92+LDArRnN2PoEAAUjsYje3C2lei25Z0ik05OCYWM/q
HQfpqoUr13tIBC8esZ0zdrEXuPAcKNGBtiH4rNa9QIvP2v2WnGnzkGY72EjjE/xWDB72ou5/Kk6d
uSFgg0RkN32PbbnnuJPJlouzj07P/dX+h3trw3OqU3L9agapLDPTMxtQ6Qmkk4Vt/m9vMHSJ/sCc
S2NwBImoHOK0ADuC+/IDwN4IijvgNSrAOrTJp8hamjhu0cgIrTp7V5JO9HdodVjBP81WMU+zVlQh
ZCyJJ430t4qfQAgJ92UUyk9GMXkii6irm/O+FD4jhDT/a0DnFgY8auMmVDk70oQjnPaLMicfNOVE
R503LKxNRm93fEL3lWU05+o3Z3jnUR+RzZc+pMoustfiUIBFXWFKjhPMr9bB2TepF1BFvSiijVqj
5UrRdrVyZu3gjetledNeNWsOyMOuba/m+hOsMXIJq/zSvA7PxOlzEVugEpsDnIZ4w5/48AxxfIlA
xuGa8KS+VJV+Qq5ml2GRhcftM+yOdzc7+ea+IbazF5SBp4s4Bnj4jS8uLPl7hLqm3lzsbfhT7myw
DUeHAU0wyl7OXOuauBHQQq4YvNVWjdDlujabEE38AJpRLS8Sw7HNwEt1+cf4mNEb4AD3oRQAdRtV
43yJxF3ts41pN8Nvxaa0FuVkb8kezmGvDG6IVyQQdGZt3bPrJtX2VWpgKW5stKpBi8ErXrj21Kwc
nC9/lhiNKk98ZdgMdTQaXO53mH8na/yDqdyu00Ne+NcFw2/mMnx1lB7uvIqp3HoksJnoGTYgjG+/
LfbXFjJbh5R6wUpdjUW037J1lDo21UfRVkDX+V6vQWR/dx2UrGsbBrluwEC+/kSZxvvZ5Opq31/A
a+/FHcW+BI7wLsqkPL/nj+R+N3tWQYRCO06+J1eMct6oAgbRHng1ypKvkWf7z9ea171lCGsi0eN4
d683OQxyCQXltr0cIICbC9wEurh9ixZdhNyjNy6rIiiKbBC0x/oR8OAGLeu23uEb7h6m/BLGFzmI
Em8nLhPt8JEbe6XkPD0RWz7h/NPJnXhjzyJf9tz1D3/a65iPqX5N+K7b5kiJ5xszDFd/SvIxAV85
IXez//zL72C62XoEKQhtu9T/Lv4rZ+yCWPllPjhJgtA7eXwytJZPQqOcAthzCmZilKcy1fkJVqmS
HNLsRn5e2KhGeCueeBB98vrUZTCJNv6ssHPv7m1goryhbMkdHCZw66NbSurG1ZlZt5KDU+AVyxIo
wcADrFhGEMIPNG6gNmYlTeJ04jRflmKGyC2Z2sYnTibj0+J4h7Yy5nAGlaiocWZjFO82g1roNS92
okSNgE0zY3ioVpsiO5SxJpXxuGml4SRdyNF/vtV6DjwXzcjdgZTK04QtWo2A/ujWYBJbpt8MpUGr
+aypM7yIdxB4oZPamsMox2bT1/nXdYbNGvPtWJjsv2rOfcjFY+ia9t8Z7wQrGxLyVsUX/tGAS22c
E1awF1qSKekh+RFdjYHsKK8/RCeknPjrwgajcFaPJNYRz81CEMnBKzhtzdeGo72CDuCkWu7s0jM+
vio4MIYCBA1qWrbJmjSZPsFzSqZMGoMoYMdnNCTcZ9iGr1uX27n6Nydm8uqHc5BE5K4NMDzF93Im
6pmYLeBpv3JOz7q4lnpf4FEu9uCeqf/rIkIa7C4VhGkoEg8c+u6KUlt+nIqQOx90785ysn3fBNQw
8cFJaaVD2q2QlydpitazFRkLJXjNW7/nfoaSnFU7/P3ZpU9NsC9LFoZ7rsEGydd8DDdA1rzLfmbF
eFVxvi3HdIGeMTD7FNEsKI0bPkOrcFhlWIp1X8OtL6X8P+8yyDr0ETwvEXAdekgizM4vt4TaOPdI
lIwirdvy/Ga+27TmKy+6X+DxIou6SMxwRdYVzOV+fVQG1njAVDdIvJH831j0lJ4JGxOK+V1UUdii
jKQJaFvOjdYdAmaCt7QgmnQXo5JxGaZ4z9RFcz9jxMAq0D3qYmqIsLqrzjD+6bk9faMhNdsUnGn6
PDE1IgXcv6O9qvYwxN/TO60ooHxzOO6qwn7Q/J8aiBN1pVX9b/Z/uY2KdoFZzWjA5N0jnUUtuLB7
UkaaeDJlGdfxeyEBORQ/U5kvX+zwrFxdGngNhJghktBRB6FLIZ+V2LmQzdcb7qT2N8IC6u1hoZyr
LlHDwpQUJjV9CCYqDOnUVnCTjRRFvZ6u1hWAkgHyA/N5JN1wlp0YDD3HpZmtBJVAh4q8NVvsT9rz
BwrpVAlgAVeMUUarrVBofE41QCU1dZZTMIEgJSesDDdwVRaz6u5/hGiJC+NM8q8PvqBtI+tAztXm
9d/9Rjtqfra8uCkcC0VXbMervqvrcX0M1zUdLXFYo15K4Xs23JWaXHClyHuxTz+4CJKd0fcrtVhg
USuNgDRXulzEwU0KM262aWpfioAMg9iH62G1KOp2UPnfxIeIs7FwS8V40umw4GhS9Nl2uNgdADV0
01iERXFF0by4IQ5DtAWP2m3lMtLfvV3l6z7atkQdeqS7jBvWWbb5d7xqZfVFm0SDcAwSbI6S3Wge
lrMx6J6Q+vYysYjTpdQYbNG50MA2RpdOgWcatw0bMB+YqCMlULFR54VxgI5e6zRoGAGbkZMOGANN
PGw2hgcpBmZJEo/iOTvoA2ILEdulmtg3zSG9/JcP820H+9tSwSwAQuld0b2lvwh1te+IYSeJ8hgc
1VSVd0eIwzCOhknEybzA5gFNPXR0vGGX710NmjI0s5ieiQZKVpoq/i9WsjNp0J3ue9wfkkQJ7Kqi
ZZxrn1Hd9VnvoKkN9IINRkKOxZtzWcbAiJm/q+itR9EAO3pV0LZFJzMC0IsMFC/dxTJoba03SKLy
au6jbvLS1nSw7Ivmwb1x1L+W4dAn/MNR1Pkv6Sg/cW6jK1DohKk3CdVPYPFuMFYZt0Ran//OS1Uo
ZsGegU9mA2PpP2veCqA4BcPWjtM5hsYCflgm53+Fq5+vr2iaabnp9XPSMX/5wgyhMqlSE4bOzqS5
QTVOWzDLP0PuS3XXYYLsyifzQFtqWVSzNl1l6G2TIcGhzOecidSrU/th6Zp1BlwTgJZaIX/HasHC
LRfk3eRHfyYPqWdJocCuWzYj/Cro21z9fJ3XXEoQYJaOrSD8J8Nd9mUg2EDPusofrSKfd0MvvflG
8bIRsKSfBerpaji0fU+QQ0GII4tSrIRroOEQm5tUEA/iX3ukq0Rt8OaRAfhTv+QLi/g+N/bTEzSu
EIxWa26Jpc2L+BZMOiwPrPen1yutIfWQizB3F6C77NbxRirm0E5LdHo5Jdb3DmKLKNq2/lxlxo3o
/IC2Ce0ab2cfSR/tNCnhpWXGldiuV0jWNpsBZs369wrrjf7R595GtxASCdEEZ3VLt6ruLXS2zUU8
RJVIXEK8tsLaNFZyJUQ8jKxLeLOtE6qAYYLMaiGZc19BudWJAWqLHnku2eVBPQPoE37899P793Jd
9SLOo9Gym1VAXp5YXNkkiOF6f0KHvJFIwdmdsiEE4EKIcpBXWXcig1dgj7YVf3SS98QWasGgSoF3
Yumh0A1B1fdyIRt6QOk/BMaiMe9hNwGQh7KMKOghPY4hCLRmZjNWLVXpk+TqHrUUqkB8JYkaPNpf
XMu0HFF41WSBVmMpIO7LroreARiZbXiFj3LK/Pz9sozarlyawELwIsotnEbnUbnbwdNa+oH6AiIT
pyKyqCifBvkVMzXYRf5W8vMsycaPZybxxvFig5x1l76TNAziiUR40oiQ9a4hgbNhRqBMeSpz4Q4R
LBEk3uERRIdogyl2tiwNAnsY4a00w7a6PclDYPjJ/rKwi++xt33aje9HD+7rU4fFxWO6vl0QXzTG
CrBpHGreqmZgUYxpqYPMSUXYVDIYCNybH6uzy32lL/3vWeWVHjLL/FcPKLomUg8GnXmTsuHl65jE
MwaVNHJuJvigfzMeuMPV81ooJfbrp2Gybl18NfgZRFIkR7AS6acCbNNhIhGkHZoDYJsYDCYkhI4t
WwZMi0Ws1uphkN6GWmCeKi58Q8yHZcQOQLNpoyRoRBtcEargi+VTqzaTFZzsR36s/o37hAfrr/BY
9DQnN3cSxRTiQdBZlBchpo+iHfOEMbSPCRNgGBOaLh3+iJa1rInmgyhY16yrm+c/3nKjOf5mVCzR
Br0xh8VlP0tC+0wOLGLUM/pv5OIvvEsNggBSA8h84ffLEKMeGW0SMGrZH0LtDRKgsdphEKcpiez+
IKjlVSR/d4JiNxskr45EyGNdMiJK9W5kbgdaogyxOWj426TSLYjaZ6UAnJ38x+GqsQrEsOgplCkk
XzRZZbAXwidSC+YavVOVt1Tq3pQhM7lNusyroaTNeSEWfsFqjAGAgRRPdLO3d1O6gxpCmhNkMpEU
7oSu60UlX8uD0Ocvy5G55YaRbSsP0Fl4aGOAl67okULK4t4IHfV8ljVHepMerUrckFvU03rsDxkL
LntGOM/tCunuXuL1OSEna3Ifd1g1hRkTCFKv63xRtLzQFk34rectvKzet0SI2P7BJmARXx/ll+hs
zzQV1PDCNY7d9p6+tu1yQeLpwFptCXI1gMGKTpu4JzvGxM+EaVrfhOjjv4hEmmRp44zFplMBmWsG
L5PiBeIHdBy2tIMqmZ5HQRgkw7/g+fJyy2ZX3eYfaGLMIYc2N/O0IX3CURpp6P1ZqVovFxIbsCWu
F13V8p5vph9gF7sq/QnCQ9apTACAnm/cWTZ2mLCDOcp/S9N4TZcyFrSM8ozX6/X7rXVl66B2zyMs
wrIzXe6FsTgifIqEketztPba/En8y5UgfUCYWVjGCu1m8ofbJj8TimeZjW5LaRJxscaTg7ZNVeSY
xmY4hLOLrYxyh3HgtjIQabcUzokCDgkaB4RrvtSBLsjnUE6x+dkgZ87AXEkOH+Ca/X2yvpxl0ybq
tK0hOXbGujjM+SGeG1YgQmqy3hqy37DIb73oggVP0ijVPfpRXIYHH46FlrEU0tPeM/Qi6m40Z3+z
6HbrQ2DAOaAlhwNhTKGzhbbvJb8isPod7aEFcgnXzVFT6L9zoBjha1QJBtVqSMUe10BjENFoAz2d
B5Xime+g3zoPoF05WGFexj4AokJHQx3sdDZUFhSYiSD3we0RX06seLL0Z7ZiqNWjEwBV8y08Ysif
CTBfU5RktrSeDyyec7qiUayTK+XIeoWXZKtSaQrlBFPxijyxk3wlAKamwtaRcgN6Hj5z9e9ULt5y
CHfLA43jLKXHjuL8O+AgPAE6F2vljP9FsnTqVN8qWfz4BI6icSqycAHYv9y1sl2g8S1XaLOvCNE6
dhbd5b6ogBxIl2LkvBklIhd6CWDcBVQYU9IXgugQO6rFVnTN77AgZCewVllFzkBoFnR7Axy02huJ
LXecSjXKYbjbcbQOzh/caevcc5yx1wek0eubWboHOs3sAcTvZFuIqTjdzwjZZHo3NkJkwUnVQjdL
s3vXFiJApOAHL6PTzpit62cdCzJFHgTVwbS4z0cI4mNz5AXn79di9cksqbadGK8rbX8Mk5NV+/f9
Z6V1LrI76G+KpaIk+GP43Tp4qQ+ssVQSheYvr//YKh3ho2SH49EPuZ9HClJ9aS0wZ/c3gvNhikl4
WqXHicbWAv6C3XBwykcYFuu4IEHp2/lcjyiuqrroWVBE9w6ADk8Keo+L9fAttWIvp7DEwi4bZ79K
xITvZveKSUujIGXi06X2e6X9AeUjiCXTU+RMPnwj+vzoxROgOlgkcN6nsEKP7yokfzhejdJaAIMc
ndO1p4/cQM/NrqDcm8cDkD6pZywLoIjcSuMeA7z9gucxV7O7Jt6SZp7qhIvkxhrPvY6HLHN2KP+9
UBY9Bwitpw17bTz3EgDGhWTiBID3WTmZXQ6ZpLeoISiRtUYvn7bstA/td0SrwQABnufds+DHoOr1
2v/nkCj6gW856o3ZKDj8HvnM2ZQ9gq7NgdPcny2q2t8X9OVP7aXDvFMiJZuM3hGQ8vc6YPVur6tu
XZQ7w29Yz4YCdnrVN1ifNVsae4qwuohvXvdOocuSehiDow7Dnu422YUpmXU283vNdQ/DGMrLM+HV
YBcjsVGxiZ4rQYVv8tMryxO2Ar40ayEHP6q1wikHqIqy1t4LlPVVMN8PLG9TPaNxBmaRlTDuyEMv
vvPK10HoOXCcYYA2QrQPwRzGFOjRk7BNy0apAwJgGccQiNQHyi9OK1bRsvrwwUBomXOszsKgfoLD
3veCws+3FFsM5H7dj9+Wj+DFGFuRkIiVHwIm+ZU9veA20cebZIAm+KljquQIjbJGynTLbvVDR8R6
rz2SOI4KaczV65rY264tSNEc30+64IBwuDZyHRWCyeSrN7jocHjhmqdoS4+grjH5A5IaOiIQCXKX
ed51nTIW4J96tv9EbOJ6HEFr3NL01fEaqgXKoPgqTRKTtRNGBxT9Ni+g/hOChcrc0eSKLCPyssO9
baGWqaYf4g3to/tFPJ1389ezaJviqped/xtZd/w77mJqGbBYA+EUBKOt0F19B2pRy0o31g/7ptWP
b8i4ushJkOzOZu+V3lT6oApgkcNFZlbDKU3NhXlZiGvnsQC5Cnxsr21qbqjW8w+RVUtfpXfsP2Um
6Vo2AlWJ4Z4JlyXxE2jTZvsw2TXBLUbAQMDnYD9aJ1b6xHuMmi+t8Be/SAJ9NBfulst41KZ67/Cd
jhr9f1hubeEZYHPxvCDXIPaeDD/vUqyEXYaNudvMGVZhQoTUiBzxNSs35QidO5t9j6aY7Hkzug/f
EsSoZLZrcgzK+RbuY5qrEzwr7oPZ+jcXq/E/ToyGTxlANo/u9/873dSMZAM9iFY584CjSWalxSK+
DNwZkPMUQZ7ivPP3CX0YTcUDi6MMR24rPG/FIdXtaHbrjCx/GtwXrmaJYsOcQs8HacugEmK/f3Pk
ELDtcyjvfuWsdbjp+kzp/czjJIMtvHnoPRo6k7rULi5QNOAnttBNdlVt52C35KTHEzIksxLdrbva
2psrfNH2hNx35+euqlEJUI0HA5Hi48XTVl6/j4+Z5DizBjGAwHz0Et2Aw7GoP6+TmOA9U4k/79xy
FNWYB7uRE9GSnV1O7pmCbnczX7HKDc/GR0k5pSs9uGA7LN4fJy2dhH0a957E7YStnsU0dTu8dxV9
TldfvN+73xj0un0YFgEVe6llwqOzjgBsEu2uMm2VS6KIUTEX3PdWNTJDRUqLuHyD+2dCDqE8Hssz
1wGtmiZWpguIFxDiM0XnHqqXIX7SEhi/JSQU0yu6+Ne3p5/6Saq6jBzZieRlVnZL1xg7+UdM+r/I
3YvcYWBbaIeA6crWKXFytwpjqSGCcE/rAr6ORzibQvh7yzo+jTlz9OP+Tvrg3nXlBfQWelHOWQ/u
XKxHDMbyGlVKNdZU9UsQYNDjnZmI2NmLgzzi/jS0We8xZsq31bPvpZ5nfvcAgZU84FkJLHwsLi2S
/HAKalXDcPudkPyS/2Bt/2oKdAuC1Y5xhbiYj500UZ/zcWuhWZWy6c5dofxKJ6XUlZii0hs8opNA
pC4B9BPzQQgagTZjgqORei6gsYRGzqdsDuD+TEEkHwSmf4z0cWkmZX0eZ6fiu+WYNImM3m2irY3U
kSGM+sRjJvn31AmVBbBpcbS8RjuM5+W2b2ox/yQLqeAIqZdjJY8Aj9OS0HCviLBVGpnBBF6AxAFE
3ArZdo5J+LKadArDMqk6/rfFuwNOSc3fB6urv027Asf0VC90ZxjjCVRmSsB0FhVb5A1aAxn6G6xC
YLVEsy/K33QBLYmHNe/EY/H4Ewj++L5LcdAViZD5VdBWfBMVHiTsJjs3F5XQKL9UzjVdQaFguJyf
6GlCbuFr5kfx0SHCDhSxVJwp1+MmgObwzKfsW58bhNurGaYtSUzRkhGegKtCZn0wbbb6Xz/YEJ09
D10UtEV+KofJyhUAqKa27kiQOmUj4WrxuGY51F89lv8HSnLDO7rJhRaOOE1kuPlOe0O58vY9fqjr
GqjEQMQqnN9BR9EinXqh5vmTOD3B5DlvF5Cufu6nD1HGdslNghU6Wvmc3vKEt3e4VjfRXmR4XbNz
JN/kJK6XAGo12irtwUCUAo26mgxz68tWHifUK6kv32sH/z+NIP/N8HGV/VLmzSgqyzg5Nqx39guW
LRA228M/NnlGJXpQQr+Q9gAoGDXSjqdqCFSnpmasLgdZBI1GvNyjkofMBaW5Rho+5ZJ3XlmWdFYu
nHm74Cv8jLAL/VydhupUhpuyTY3PYSjrwyHpgRwOCcm4iqgJxE6Xy6yW5CU0eLYEc4cPl5KhnPPp
GrFvtNe3oHpHle0a5vcQdnecfXv7KT38gWTeJaxpivqJP58Aow74spj0I0kOvoTP25ClOcPIFsaH
nqIIPbivu4K4lir4Amq7ibT6/RXME6FjibMBLWhx0jCXaQYVNUs0RAEv07qjfn91YglioWRJpCAe
BoZIQsoAlPI6vQL9gsg3Sk8AzVoQEc6NJ+YEs3+DuwcvPgtoLvh0/nLFxFM4OfcoNFPlK0U5vAK8
2esF37Hb3aoL0CK7kCzLtk5Z2fFcaOTmJQvFBXRwdetguee809oUyPxHr2MfrbiXLh5/rXr0t7nY
+GKDlviGzuyd4pLzbyu4Tih4Ks9eKAU/sbAXIoZBODXYCA0KDQzRo2o1ttToJuhBQGO8GkpI5Oqh
z4dm8nYDCDodg09DxClELGFo9Mw1xQX+q72nNnCXZKQ32Sxls1ZIoVWnSav4pr+m6qYb8S59dmAm
f/ptfPEmRLMQd4zwG9RXGsy6FVXtHLPql3TOY+3DyMXzt0ky3FLcUVj579N8VWYcPngSJYrEX1xD
JrxxgmS65fsY3o/UXe76dwOcaWnwLf5S9K+qnGem5fx4UfpDksWAhcg429lyG3P8IO3YUEbN86yX
n1bpho2GkPOS5SUXhCyCqDLBL1tkyqhO1rr3vd1puLPpSMiu+YkAkIuHQxRJWIG5Y4gM4i9b+hPs
c3XClO7zys12dEp9UufHeReIBfaVHaNp79kSR14OofMpZlHYyeyVhk9uZPcYj05oGNJq0q4RIDgJ
xpy0IUzv1qFRpeQysdMImAzJR7ZemL6H5l9aNAGpoahCkP4TvvznM1c2f0f6BK30mcNxIP2FYDXb
hFgg3yOjtDWYZR9/XpBeqnjphQHbrQzFV1ulOj12iCc6g0xFokKHbsSEBlP9A6HxlvnlWwIVe7Pb
pM5jmos0OL3SQ6nNnIj0Tf5H2S7jLT4YA1YO7z/Dqamebf4SZIICLCB4cgt0yKzaxYMwf4fTME+6
lc4LLIJYcD6ncPvz6rRW5lSp1dOOvPotumdDHyx6DYFuenJWii3fIopmiaU65bHMVmkPLwzboCqA
LXmijoXOKKSxrbkh8SNV2+LrUv9BNja7qEXknhR6yh4I/9fadFeBaD1J/GowknU8iVUe7qG0BQp9
tLZv+B90sXt/Twsj7TGM8rwJg1ZZvJhiHM4Zub/8S99nIeawyMNtqJRyE2Z+4Hc4baJhEVNScUS7
vBL7/nAcW+praw/mVUbSSjgJqk2nKaPGAiuOnUtJOLQWxXHbkzfQqqLIELzVQFnXFWksJ/nzQzM4
jFrPJO299f4YbroMiP5XaLDD/n4Jy9XmtABir+AFho7/j83bCI6BXxPneukPMcFoXJkuIkwDlCqG
gV38VxYlksU5GlAb71XmqxJ3Y0cFMl+uyVeSbI4F4HkPwzdbj/rlUg0mM+f5OX3g3Nh2Bwwynmto
fvRQrxjXTM3qjNdYUoL/q7Q5Ihimp7SUBNuH/2lR/WiUM+FLtsGUUiMYmFBKLWML9O5RZ+3kproF
qD0Vu4laAeYmEOIpzZrY2bW69jIGSHSYAaGmghPgyRa4iG8XH12PhOY7bEs6E4L1KwmhF/zELzhd
FNomNUHfx10ZDC5ZYkSstIbuL+YeLml7syM3XEUvQfXL/MDEWIPWFpp0BNNN44hiLjJpPXdov7fP
/1C7uWPd6RxasI61oR8Gq1wOLEWfSkUCuwDEwgxO7rfBySK+Jg3RA3fhagjpOsXz/FuGgawn+1R7
/iIoG0sTMjNGcey7AEcu7eSB+99Z8SbB4URc04MG/aRVkPwUiyiJhmmRF5qfRBJeDhvw9/CEhwM2
nPA9FZIz55T5VO5vmHoeWTCW7OwopO8wFO8U98iZgXXnqvhTzadDsRtEd3bo2wVJ+msJpqn7NAqg
bKuMaOItnI/4Mq48FLpUUU+clW3sVlaFhHbZ8gy5fDfwt0U8ZEJFtVbgT/yOtzoYjy2VTg2XAuiz
PbVrPRv20yqOaYWdADPokTP7TJ7JmK4DxvC9HIjy4VLdf5ZRmS9I86oVR+pfisU+BCwh1oJ/SktD
c+cLddVmKs2/JWx06Ll6TXzmz9u1C/SfX5h5rPCQV/7uSoz5fnY7uyUO0B7BL9bDAw8atEIWBqfM
pX2oon7BYa6Jq4iCGtG81dR/7/vcccyAipCqQ+E0J8HHUwu+jBlNVncmHAlX0v5n/d3GhG49kJLX
3lo5JDpbx85AG9DfZCVRACB9K/qf5tCSctliUe+cmF0NFAYLb7U+b/urJkkZtzk9rjr923TpGIV/
S/RNvqMsLyHP2CSQ99eeot/78BFi46zvCUfDHRSMWrHtnZv08mcI3XFD0Fq1cTVa+/MzRKbn69VU
nt0pvTcwSSvy4esVch1Yz167NgWqpwa5tDGOGNP3lo8/gDOkkvd6WjmrTvEurYS9wsV9SX8aN/rC
6fExqyr3pbQAkisJvEEBpzJ7b1sd2zeQKpQm5fHKnQleJc7hDC9Fq1c0Zcw52bC64SL2bgFT5SbR
AiApL8hcEgnirJm1UUePzI7Y8q3HeeLIXfAwUQiomhpJ/RL3AjBk842iU+MZhs0wXIentKD7aa9t
NW1iYd+9ER68H4aRe4DKBZpawhdK+no4lKhSI/piRNx9rCeOmDhAVCut4CEkSEnajm8TR9q5O/c0
nIvOWlNu2nKEx75mn7hpdSalWXOfEXo7irFFuVURybKqo2SKIFaGMR6iJJBeUohYjcrx5on0z0cU
mtojpNdjc2QpnesAgZTD8uTNgU+ex50vkPcuJ3v0azB6dFGryxedhF+VzSGV4+p+rHEQw6iJqbY7
8sOWl0tTUGscuQ6kQKVxxYPOl9e+dhwQ/nzAP3jTxVKOWQwIW90BRi9hRkVJcpvCZLJDZXep+bZL
rYrdYrbdLgZhNBax5uO32vgRECkL5h9LSjMYhOFjRIQZZjsCR7C8STN9qHONQDfgVRvDPydXcsmd
tzwJRfIuIk2PBf2Tjk1/1k6knfl7ZpRWOLOgj6UjWuObY6zEIPdxZcx5OY9z7sQNjyV/D6cW6GjV
mCEOek4ERKnnZD5zwG2EMYookhLYuplaPsY+9UkRhe4De/bpu4KCu0ffNXPfP3DWwGUvbz+sTTi6
O1UJdnph+HGOeouwuHt+yAoGMAVmZYUoHB0NHy5Y6ElyP8RTLvSmvpo5gv+WTUOgwqy4VhVvnBMP
Wq4UkqIMbdjWjKcF+EWwednCcAcBSHJAumOcRLwT9GdSDJ1CtMImx32sH2H/zDW3qM/FdB6xWH1M
sVcHz93mOGWYa1Ua/MyETISMf3suShVsbB3NRWjk7rWWvYSCFmEV4otRmjnNcAGIKTV33W33W2jn
bVUCzplM6LQrmMG/FRjrJIAijkhAYttU41JZGk9mcbn50AK2/GubGDznHvothm66B6wl/9rLtbnX
Ohli7FI5A9FTbn+nu8NhHbiwONT9XcouHxxP56dg6uKj5y1MTg0FXoKIX7jmmujULuwryikXQor0
o+J5c6schcjb6K7IlC/NgsprIbFYKPi5qO5c8ncEbEjgmcX9Si/D9JABG92L8Wm7xUc7tmIhH7xM
6MBq5tq/dBHlsTsbBDRJ9r7mT9Gscloclx3KL1Aj7yrO9RMouvRsF+RZ6qPHYaMud2mo/AalOwpn
o0Pz2uLG3cIf4C5BMGGb/NfUHOv1MW9i6bx3PB4j+ta8o9eHzyejnjiRGfoM7HiaUQ2OmDXkRVKB
jvNGlobIvmne9DxygQ8qeyXiZMi02/UducpQG7Ha09i7z4UB67bXh5y9awuAmM2aCYwixfhTLPAo
RqjfKzAWNo4yUdqzCQAqTgCs64vhCk9NyACYbkZXs25mAkSPyq+HMUJAHFX0X21e0tz2pEESBRKD
yZstCtSww9/4/dZTKvMdRDIjVSN3wVXVUJil/m2JrwVvZQhTODl4SLJWWJeazWrncqWQso96Dwzq
f4aRDaFihKTBdiXDiTqu7L4RJSbd2nqoqU4jP2ykGjIWkT76JIeDKTGF5G/Wja/hYd0IY0izyorz
xkzwGQKomX0BB/Vkpel+HQqHGKEtE5JR6rN+jMVHNsD366BTeifosW3A4HDJZrvF1nJ2GFSHRz37
VbPMtWaFz9WYIK2/0Xp7OH642gi9Ke558W8h7WB9rT9/Mmu7/KHQKE0+WZQYCEN9qTqJbbXqCpvG
J1MLesEuIKbwspeFIrEYjja3R/OOeutMvoc2N7zaa8uSoc+zDrpklwyaJiPDYq9oBURoC+3gFD88
LiUgk0sfDHvKKOdpgN2o2POfFIZXmQcUgxiVZCyspIg7FNMwRAFWg5UNv0TBpYrGLKR/iP7hzwlb
kOwlfLHoE5baYUB50eS269GUMiqTfTIVWBZqmtXUfWW+GRLw86CkDSoeE+BJTIVhfIR0Qh2nu1RK
nJyt6dOnYFZrzvAZhZ79vOlxHb5QNqj98Oo7Q2qvM2xbHaek2NCfWf9J+uXkSLFGNb50VeAymUN1
81lw6zp0kAj+Xgiq6cmUeXjX9V9UXOtvHVit6PAU4fRDYfJv6YKGs55KFYOQE7cKBcEKBGECm22L
mZpXzj6wulGSMKCr0X2Auut7+x0hp/GaxnkliPzByCnnWvBePdcIswilEKC6+JhMIeKCKKxquG3V
flwQWvi5x0OV4ClJJZw9nfLt7zwe1FI3P63lFZZD9OMkJ+lJoJk1zro/CKKtGf2IRD5bqncwr8B4
uF9H8mqXhXLrZtMkHWBQI9fii1cIPFM9S3yQZWJWSzRIvVN2NyK9zRZU8oWgMPtTSzNz8NZyDsLp
w+A/N7Qw5QU//mofpGrvxPrP7c666UyJlK7XnzyqhWETNgTfHa//GdQNRouNbFFe3WApUkY9dZoC
zWeCKX+bOFY8L/2rqcjmE9IQbafiqPp9nFOer57tbeRJ3yrgLwXThtBKtiVE53j1ArsWvaG7+zT8
bFXH+aswU9jxVIKUEhWOvQq1ep7q1QydYqwZ9/cupAbyPagjlsqNws2GcedyaOxz+9wfCog671zY
3gFtFQ/sU0hxfqS239/TqHclX8cZEpu5QRuUBHT1hNvwwyLhQTdKVYpEEkh29AnXE1HvkH4nmpy0
FlKVmkhYn6SZd+0rsfMaHnwarZItteXfTCGNnZ1Oo8QkhTd+afy5RfSa7gFTEYvJcw/dGCKW2kcO
pKA3cvMIqmEnf983bxbjH7+F535zvd+y7Dr+HbnvoEHjRo+I6zP+srKFXDl13KfycdpipobEOyaE
A8uLe88n+cQqxlCBf+J5bs6snU2+GKsk30BycMyc7QNpuJAP1PVsNqBj6ZNw0Omd13dqDJ2zvmYL
PVt1+bqGwR4a9FoKlIy/NNWgCGSDi7VXICSliVORlnBGn7Z9uMhZFgM9UvB1dc0qhk1dlWafI357
I1KZjblimXVF2pBY+d3wj7Y+P7RCQtg3owzFCBiZwZ8bsrdyf9jzV6XfPDmHS0/lDeQq3FnyfaOz
JgfuJPdrloPmvRaKrttvcDquoK0zbNkbIaJ+PA7kt540iMRMZJ2uoUu2HKFWjwobr/OfWpiI2lya
UlhcSKY72AucPsXO3utep6HbHtBR1fXx1agOzPq8dLV0QDjwRaMSP2O4+f71CFGf8IskK2MluoSy
wmPUUbPmXGb2XFukBh5Mvi7qoHW1A6blLBWxFqvp3/BbLCLEyGxmTVGRPI/C0r50UjN71z/G0wxm
YwVKfpRoE7QjqeeYlF86OQsNjIk9PRnpLzdyUnKjndZOLxkTh+iQculXJ7/YlqZNjbNs1bTsUgRO
S6lWBu836/Yq7Iknx4kDJ61hQVZ34IbgN0qA6MeANp1lU0I3il5l+jA5qeLPEU0jmYxl2HLXcf+z
qWH84kDsekDqv/NG0ZetHpslXFsOn1uPgcJ18SYYMGVB18+IuP61C4DexnwDfBxwCPna1p4IBOBE
pM/q+XlXeijocrsue8CXXX5U4dQISyrN+wCIp0zr/EmkU9e3lcroTAm/rhjg+v1+RhAn3lcj2Fui
C3uEle0RyVoB3y9Vj8YC6NFiSARVkfWn856fA2ZwXtJ18oay9kZhXrZgiubZ0b3dt7hDlkGRMZTo
p7OWNVLUZBDstvxKyEnB4scqAk3x/Tnua3s0pWx3kIbMzySDK6W9lW8aUXo660F39ouqL8Y987tw
EqZEtmUEsI7zzFFPRpGWnPrEYs1ud4gi2EJm+GbcbNLGE0DZS8oikgrxqgbs14HRJmLGfqrFQ2+A
PuUQjWRTAmwnwouCfpxiY5BEj94F5u01jdlRgaufjDqL7g7rRsEA7VWRjed+S6YnIlfezY9UKgC4
ng1p2Un1uqn7iAPEmnMsvBV0QTTlG+PSVSPWwH+YtmZtMBzGYlWfJvf7y5VTShzjQw0jLmR8PJ7V
v3Yammkn1JCnj4APFCknsmGSG9A74CafInrzmj5Uc2QE0CIPYg9QL7jFCArnIxv8v2X0F9ClGag6
7iFF0dci1YFMKIBBLr7o9jsD9A75W61QKdsO3Ne0fGrsuB8v2zaAM5ase5xtFL+y7n4O1N4ftG9D
znNUEF+gMXylKokCZy2aa4fB4qwEUx0ycqUTuj6cPlMBZFQKqw4+TtZcVOd9Yh3TIllywCUtHwpB
IqNL531RxIdS5qB6KKIWbHLYYBZMBae4hqivEPQ7yEiPAxKwuih2HjgA0x9SyotZH5tVudHtja6x
DKEYlSL0jCOlKwIBOVOqn5M7pM9wWVpUhwauuOoMymsqBmFd7a1mtA5zUgRwq33R2l8hJ2zm9VjD
WiyjUnocvEpab7KB+VhtfhoFPx6sLvohp6FQi4rmBuHWHSNO+qP/azrXkitG+dfA/UwPkK18UX89
Odzxtp+yXmhBRyv9boLzDBK/csNdNpU+AEx4GaCzqJWnnClyd2kOewg/J3HOe1LislbXrhtEYg+8
CytWaTs7VPb5V9o2Aiw2DZiG3ye8mmGab4rp5glfaY3TP3IaqXXmiZ9ojVs1UEOC+o1bjPsH14X2
nI/pSSyLvftESzlIH/v4DOc7pCP69UkjJ0VS6HRgjAneE/aQLum903z8U0sY0p2As+3/9xSmROs/
IuiRNKL4ZN92VYFRTnWCG9rP7Zow9YhxsxUmMRDuzjEFhsEN30oP8YZDWskeA9cm38tT1XCG1fag
QeRAbw3Dss1cANTuPkVMySepPjFBG+eB5UhKH57YXhHfj+WnumnsVwyjOrzI/pbwPKUMk4Drav7M
LR71JBdU6RQSOx98YRfIauoSHp/DqVxRcSX2gCyXuW+LLFdibiOrgawK7UMBbkeueNWsgm4TP4Ea
XXysh/WorvzCvAlvXvN2R4R3R0gKYsLhy//Y0sYgSXGbkPk7g3RLy6sOybfA8yIRnUR7c61enWua
4/TMrCECZBwuFiQfjVAYY2LUx0w77mBIlmlEwnX1v2XW0+AlVScrW0LpqOt5NbDcs3aw5isiIxOG
QGgQYg1720gs+YDG2pVr6N5iq2D6PBELgdC2/yNsx75V9Yk3BU2jd76IPw1aXx1b9xVD6miXEPW+
unH968ZrixSUU2bGJPy341CDyXCZrYy1GljNpJ5pRHLsvoN0y3PNoMtaKEzS3Z4rf5zj2Eg0UxGd
arjeyUIzhFljLwMcKCHTk0F+bvrOyhDzHe1oUsD7c3ih8slL0tQAMLM1vmXiVozY8IV6BEVbfDZW
Xee/ae1JWj8WjxS1NP1ToolQ7On0k2EAJdFuCwIxAlRWaVhsf20w2JwS07yzSOtEVWqxjtVeQC87
GSgYrVYowQ0up2bbvTs2T63WydlmSEeRASXMf4/kGtulFoEqiSauJwMhNhtVP+CJMY/cya6+QaVh
4mXO6nikyjZRclrJzqep8J6SIY0ZJ0lLU7y0go+hSI19SOTqyQ9Ezylx54POrtbNpwOq/X4JjH0C
BRbu6RyHiniC6t7qPYlQNgZ1WoErqvUYa+wGyEkVOtV2RW9FUx0ErSGPySJa18AL+D15eRBxJ8IC
TzD1coVjP57mJYQ7CYll6uRzuVRqGY8R/pH41lOctyAxVJdHJGfOwdyI9t1rZoDL9i4vn7GcOwef
qxb1slEdp7bWTgB5ZJhQ6ygTaUOZRAQ7CI0h6fOTRwqdPr8BcKL+/J8/3mOaYPMHdLoKYyHDMsbG
H5npL2D6Q/2vQrsC6EiOkujRNDcfqTW1P8J9buDykauOUf4CgB6uIixWGFIz+86cyaHwu2Xcd3YD
WpWdXhYLQmvmohG19bMdkPMyZCUujIfxdgKhjCcTaul41KYTIUWNrXGbuNqva0iiT/Pr7ILS0iA2
VzBoYljqCHwZ1bHCdAQwiDz6UBoKlzkGQzGlifgOLslRfF+nrL+SwKVoMGn/nD69qoFhuEyDH9Bv
EQ4YUd1dxGnOCWNispZYP1pS3clQX1g13rYbjo4iyHVUBoCa5vY3Q+bXMrAEAkDc1/h43KtDNlek
L/GMgiShO4Ah3uQNrALZYYiztcri0pcJFgLhC1khwMIBM0PEKEmTxu0njRqb5P3mEIaz/TTbA7G1
dzObo8w5TzbSatSYgmTV9eDUmuRkURkaer2m4OrR5euW6s3K3H1mxDWkbKnO2YdTqlvRnc8L2Hx1
bp22cC1NAtNxjNZTlgjT7HSQ182ncGYYw32zFP2gH1FaW24D3bsiVUzgOhABBGj/Rbokwm64YqZy
2LsLBR2sqOHqSiKrOffLj6LoZd7xncwvWjoPdd5epEr/AZczn22dgTuE7vUR3NqSaiCl67qmO/Pu
3LFTMOQ9qXhz5jD1DIKtHGeUwue+E5hYjW/gMPv8GBx4Ha8/Xpv5UdIj8Y7jgrGmHdhNJS0oL3O1
VtcCpKx1GdmJ0zm74X/BqPgCe6Cp0SPiqVWXIje7jeivqfc33E0B8r7vfEgNmVhrm6CMurkx6syt
XsWIPTqBO512q9bu76DoTQetLEVz/aAmSB4jAzhmlfYFR8bRV8S9crADaJhLR9/rp2bAOgoenDKM
zVgK+sHm1C5ABR+IKxzcnP9A4M3qhrO2qif65AtEW/sbFjf2Xa6nfjwCAVO/pmbaoeA6SJhLgkfw
/pHMXYN41MqfjyHVoZjvRItdfOC9hbZnD1uXumh2uv1ZIH23X1Q75UvgvYKo+VaSittw6GC8t8jQ
XqmvsYEUzaegV1cQD2kZ5jpJfmDwII4UQzosqnYdenBFAXVby1cn9Jq+L2At0escePNrjSwBmLrY
sBUS6SkhBFnIA/v7uXfC2L36M3RRegVHgePDkhL4Hbg3oq0sWvu6/hhVbJAFIbY/LSJYsCLgOkHo
mXpN1hCmJSiLL8sLV5uaJIgqXaC+yxdbphmfTGK8hsTyvjY0x6VAmkFVJDWmv0LthmqpERAmWXRa
YqxBRbhkmclRQaooU1QFVcPDxudiHWK7v3w1YwCTcwVgaCtUymRu8YAJ0VR+ywQmRzZyPx5UchWw
TUHDiWzpIhttDLxRPq/imToWrhirx4edZyH1Vga4iqKMnOlTLef/A4rz6ds+RSV1AFsBRjliNkmZ
OLqjLCWozQ6CTxIZqZ9F7qe/t21cD8ynTXLF00ymBGQLA5hWid06aldjVfEFlxTl7Eb+pRNKM+Hv
j80vs4gqZm/0xoNNZJTOD+mMUwes59ACMxCpV9x0T6ocJBvfNWwvHeG1lBaGbBFVYQla5Y8f7Q7i
wLP3vcbNCi72o3Icbo3YVXaHmGAWUZpD6hBKl4KrxIqJyJfHosxgw6wMpiC29/k5ciPhWxMZ2m3i
HaBX85YNq03KiTZD5OsVMsGZocJKgdObHwfUug3OtVvkL8BEqMvH+xnntofYGUeo5jgTl5VQoqU3
3YXJzc/0rT864e57RgQcZEiwE2QOOJq8nvva1fxLdsYuee3HePBHhHxBAKqzfFC7kOTn258S54Re
1hDR7mTW+BfJCHnFxhCyeBn70+ZtaI8LajxbO8FA0uV4SMfOp0Y9ANUgYtcSM3hW+EbJtPO+c59t
l3uQPoKwQR9LWaDIHhp1B0Z2hwot+H92brt+d/CKRzCqC5TfZ2wk/bwsxSXC20LK2JSvCxmBvX7i
88EqHhjyw8vVlnL1ZHLfyWedlRAh5kTtx0L99Uvm/zEfBE9RsfAPrL+5kWTOI3v71J1DovyE1d1K
SsAKIzAF3viQfRBKknmmOCctMsFGCI4kKsx1aTlUnpUMAe5xQKl65ZpVPJsqOREIrNBYKPmyLh8Z
W1KAz1JQra+49/mpbGgrvmIZ7juaDN1LgGQD5R6W0oMR1exJre743OUE1aByh7WM9EYZ80za0xL8
pBL4NQmsREobkmW45f7sU/XarZBMGpEownmknOq96m7zMWdgL40B+HtXj4KIxZXIQKbwN+9vdwvx
VEr+bVBQhB6u99qRAG5QyzoffrY+LcsvGS1ytEJd3CG4xVIrbxtlc+IjG1NfwzvabLsWWG4cbZoa
a9lGf5J6xkRoAcKya5aAIqkzehN4uYyvdDcIcLl4LMxsJGQTFqqH4Wyu+J+9iElL/2puyr7WWqYe
JqwsEbaoypAAYCVLXcCa8PfICx0GWgqB0FuXT5kuImM3a2JOYveRfzCxtIg8eUjm5E5d5TnhRLlX
WVp33RlbmGSvygbGDvIhE1FkgfmUR2d6Av6uOLZkHbDLqqcQ4j6xg6z/NORxbIXwO8FAEs0u0ZGZ
pc04tJZySFQSMKxRpjouNpQua9jXDpZlUZbDA/U4HO8KYGi6tNJmZzqd94zuLRASwp2MwwJcfzMl
rZ6ksHMVwr+hInGo1StNz89sAnKKdm7IQrvHeYfrUwvnlHBKZYpwlT1ZHHXQ0RbWhMDVXs3hWZm0
N5DFQze5sAHUjBDibwBz0ulKK9vNP8C0qJgzYZAx7jgJul9p6OUSFIRajydPXddOkcUqgwEHF46m
O9lyWL2/U/YfvvDOuSmNF6/NgaLUoJD0Samh1bAjqoY8VLVXL4RhmmtFyYj8o/LXZFpiF2J0EsfD
2lWOtoYAO4s4PkMEpQ2GBoN8+7KmIwL767D0tejGUeBH+Wmn5ojBh75GlU8OiHtClWqkyrbb58ci
DM4zJBRYFEtubD+YpcVl8GS6jm7vveM40m/qZp3mbgcagtmPX5Pmqtiybu1CYlzY8GGV9Z9EapMm
SOdaOi6Gk4HnguDUv3YFGIDnyaqZzWbvlJ2cRqq9ZPe4T4+thvZt7yl2XWFG9bu0q0AJVCRO0bpv
Mth5OkqXsf5ryH6Tzq340lTPCO9n6Ew9pCaNMGe5mrFQBriYxakHyFFOcQ4TR/kXMxS096p8putt
e4haCDjHLhF+/JWvc5E72RucmMOECw05yoRkSCH6FIh3uSuTilX3rnzEJcKT+sq7TzI4xu2uqwXi
hfMXuzpQUkw9rFnm8yt7dDxFUO6CBTVmliO9eI+HuzR/cxaqulpg6++DN6NhL1Sa9Gb/8xE7wLXX
5DOVCmCJvo1bHLn+MZTXI07gkb7ICfohDowLEta5HKxbTPZDcf5f8s9mYMUkFVSzZESe+R853cIS
yW+sIwFEOyETmojX1EoF7qOQTFIN8lqWJs+SzDoLGB2UBBuM0g5A5I7qGdImVCuh0llyNrpNCa8i
AYa1UnBQPoLVPjRtj2trkLZXFDGAzXiA4KVuRoSehwnJbmFcM+b+LnkKPhPmibTgw1qlyqWrrRCw
4ChQUKfSn+rw9LHCOUxOMwwAoXPBF3pdqrmwcB2iUmNGmCkiWVbh4zwsAtGEvWuNnZu45vbrc+W4
PbRRCk0lEPALW7yX0ZflcP8W1pdr4tn54prIAY0zOiHyasE8LQ7lGdxM784N76P3fiMQKByKih8h
TZhKVo6AfoCC5/9dvdZOu7CNhL7kyPi9atUi1Ee0A+itYDrLuzj4W+9V8aw+Bs+U06KXIzbenWNS
ZfZD+ORRp0qS3hP+RM3paONLgZ4dW0Oj2JtNSQQ0OHqHWTX+eCAgqDz9M/gDVPgd9xdHjC89Lboa
iS6vCu0JJn9RYWpuEsiKaaLeQJ81z+rt3ZTjd6Ap+FrHtrCWCz8yLHWzZspfSnN39U245o4FWGUs
ZEuJAv8gYzfVZuQm2lf7b3sRNJJ6YrMpbIJGQCc6CrhrN4MSLUvHIm5ZaF7FYcePl4Bc07Oe5YAP
snbT62eSPtGPQg1IQ6GaUyZh9/+UUZ9ouKdtJrNLF7MMnAptj57gDTFSFI1eHgLYjWEFLMQ24Oep
L2/LBcLwoF00o9C1v5KnM7QvM6tl7NVr2DYz4Bl93QfqWdMZAfp4+whwln+q1LMz3zRWBmxyAomf
d76nYOwkI6Ihl7YNRN+kc3JtLmADi9gD9+nbvHNMMFQlilZKCe6M2r0xfj79gzOAVOnwi4/+3A6Z
vtDa2CF6difW2mUOwzJFMPxLk5vokk7HhH2y0rdTmocoP9SrVAEYnpurrTsQsXkpvA5yjQCm2PCg
MLHyEDU29ScrZihD1mo0A1h9/mgvl1xweVT5saiLbodNbBcrr+QfNfmniq0GZhcKVdnbImyzOP2I
TP41OLpkKcJdbiPRFqpM36MVizly8yR1vJNT4BgkINCnhdbYxrOlcLD6ub0+nh+fuW/aNId9YmdH
tuiUZ6ZKNEnBxlqrbMPll2Mg/f805qrM3VV0Gs9hwBzds58qDQD2aGjpz8gE4scbmBVsyAcUeHBh
tOiIWOv/wQ1pOBZElipvAGgQXtDJI8zCunC5qlNS/VNhlk121hCU/utB3KJL18vxlDbvb7PBAfqJ
dCkb9P6/eccHx6iUHDfAfibt9rdEBaEN3L5MQCsPE1kTXtE4/yYHOwLb8Xxdco7Cybb2FF3Y+psh
AhinoMLjyGYCDKiEnu3p/Mz6EonVVQG/Y7c9o1GLwph2fFp4jdckWglgqrw7+ZXb0cBLc6Ds3nFM
thFZRVJS6b6D1h8KqNlFgVkEPr0VByx3PXoD0OPbg7uixewjJrKNHTMTYn7AUqDg4Y/tNOVH0WoN
TKn9Tt5akfeF5gqEUZ3MRyDW2r2cr34nmjwn4lOLn08CYjwCKBQ6KKIA7rpXrhG84v8goRPHrtgq
R+4/EIi6J7P3Us+BoSpwKNMhVYs2YJGP55hDX0SnmmBKuInOjPwoGqGj+0qZSz8VVAxIultBaxyO
a7Sb1i++WSZSortIcwQUBY3p0PNj6s0I/FKbyGwD9/pN2eyQphLJZl3Qw+QHMIC8v7HdKe/+iKVr
n2I11zG4xLDF2XG/LGN5v56Cutv4C6taoTGi4glohjV/kKqCJtdjCeYqPrs9/vpGEz3OAG6pKk7y
VIe6PTs6GbOFZwagKcWspRluE0fassUXwegAusl8qhI6NN9kvKIZ+ncMvs19nzKzg/DhfE0wRQzC
l/3iDVziIdTXb6cLbXyryAff7INzqFrvmO62F25rbGuficnQqvUks08Rg+mpdxt4Q3seWonUUaEs
eSh+Kv1g4n5sT+lhlK+B1WvPnmzhCZjTx5L9iBnl/ymkGcTiF6JbqvCiIYsihy/dfV7HFZhlo80o
0GdHp06xQRhnJJykIS2nJmb5788xXiTQUesLhtmg4w870LLDZMSmzb1jMVj6pHcOKpaaZhc3GWmJ
e7UxHuT3KP96TZ7CtwEJkU6hpG0r1us3yo5F1v4L2R0zq6n4RPFwKrOgtTblo8Ucfz6Z8vuq/Glc
5kdZjOvPjuE/6hVbkf0pYN5/sI9QKXxFSyymlpKSC4NvcvYArqmqhAALVbJsdnMuA/KdVy93FGAB
wcrHtzdjY50L6TUOHpvGJR4kufZcHwgnv7O0O8PM23Gr8J5XtFEe0C51EXsw6eWetkfgsdawlbBG
JNOjVYuvVKEDADoNLVpeh5YKPNXL6FzmPWbad3DgTOlmLtivXDYM+RJA5bqah3FeAZ2f+B1OyaUW
0lnDO0tPeFtBdPSPu5wyZT7P3WkYo4Sf1XWA4N9iyEj+GoBw+OAqpdRmxfukksJVcmIcHDhpF9TN
gZb2VnNA5w239Rg8wlmX44IgT8mnK3OkWQVNDRke02o8rrWSa1dkNbBYM5kPkW3tt3KK1APYEJJx
ULVBFyAUJMpraqQcNOkwa5nqXQRrbiKbosCEirQ6+rPNaTwA/NMtFWGze3iOVlbwB7BNIvV9SsGF
ihKBggPRM3QH0IzXyjbHKo2Zx8FvgKFuPYBd6jeznw0OTUnDEAHD6B+Ju43QbCDtevGPBP107suj
nvJ+C8bwnT9fWY7cxdUEpDpqVpGN9raimLdWgmXVnpxzzS430HNkbLYrAwuQd0a/ROfIVyctyqA/
F7XbOgEIhMn2p6Ky9zNDbbUOUnzKv9FZKGCnbmQmz5QBb/ePO49gxvbO6wzJsXLVARfnYIqmTrDS
513wO8tBatpZhmQ68IAd19k11TmBIVClMEr8MBTxN863sW3rXHNt0QQ0lQYL8GZeg9hSpMRFCvEL
KPsRSzR7uUc9S8wevWR1bw0OV+OmApW0Tn7HfBnTfYPkGezQEn76vgPkupYPap+JKaJSGQcP66+s
4qTPACpK5JllfP7xT8eUBr9qMgA/pfn+0E/e8cMG4R22a98KIUh3mzAnRBqKqIggfYJz7OuY6bxT
b5R2n6X6SQ7ei89n5NlihiwgShrjYZuOd6N74G+iLBSJJSUK6YMtL8XLQlvAznWowivi2KuKCCKe
QB3EWhKFIpeemfqeVI/N/pL+EckPXqEb1mgrOOVGmTDboZ0u0h+ogTd6ePH//+s39JSXXDrFiMvz
AHB8XnRygt8G7OeT6/0+sN0L3Q+SbcRRAGn2MaFkCXH2DySWJlw00+vwzMvzVoDfO++tzOaUnAwk
K8MIHjVlJ7pIkqAXvx2OZtMuCZLqXFMWLPANXV9Bbs6ypFELiIh03AHc78rQh/u+Qr6xVuKlsMC9
xyeI2mVRWnahN9YoHC8qr6IyenzubDTVAblP8JrDlqslD3k1ap8seieCJJaobIx2Rre1QBoJt/cH
HQJ3f8rAvQwWcnY86voIZrmtt1EY1vMz8aE+QeRunwVlFJTtW7LsFrVbZNHPLOe2n5726SKDjmJ9
7E75PR01odzMw/i7ojtCrPnTBYWaK/66WYbxG6DRSul/p3gNd8QzGJNFNxEgfDpmYwO7P/bAn+bi
J/Qr7I4fWl8YqKUxz7qDwj/sUGxX2i7YhsLK2uCi6HIIrWS0b7Y+tr85D0PqqZBrb+g5Qj4+TUH9
IgGCTvM4I3yCWwqaGK5SLHtkO7ozcTSmtCa3bGniDdy2BGHG5IXgrDT6/Ia1FS2M97n4sKaXRSuB
gFYwrU90RJpYs+5NFal8bIf6zpmaGxkPK1GjYgUEZms5fcgF3cFGY423IPTW6ICVgFoQh8IIlXzO
iLWfwR3VmbzwlkCqDNgytkeRXq88y0WMR6kIJOX8l0TQKgnRG66U0jR4YLz6IXShRhfztWnWLkMr
7F34ZAaK1HwVr6fAhdUApeqsUFJ99RlTvdBleUDAwBQIzbylOPxsad7SKPOmUFwCUIiYLK8JVk0z
wg9VUWzrEOpdkCkChwGV50J6ZWXer8IFkVve6bM9f5yE/k5oagkIP8Ckf8qx2eG1UI2QlJ7Vmy95
+yhXX67qkXzVyGAl/PfOB8zhm/nxOxahaQ7KZ9J39PzLx/nO9Qn9QifyAkypePYeoWDmPEOWMcfW
knszFnEoe9afip8DGaQo2cxU3Is6e9sMIqYD0BhdB8qlcpR2nunctSmvRWNkxFPyHMrQ27C1QFSg
F8OdOAKt78rOn7BZdSrzsMvpBFr0hadqwk9rK8xbiIyWHy984PLri5fHWUe4HpJVwB3c7xG3VpPL
w/KM3rxJw7fiMGJ0iZls37hpgnTeyCBaKIUmZ1gFmpfZzRosHsrEhl4k6QJtp1xv4tpVtAfKgm9i
CBAdsyzSCkBxu+loTROHbTqI5SuDWslSsriWlvC/TRYM6WuG8xAmwrY67HIqEJJvnxYueaG9GZvF
+MUngtvbrPL8t70J2S1UqzB120wuiA4dqsp4Ls4OBSRWIC4tkwU9+EBSbVSquudWtT6iodMvd+wW
wv+4zKUOqro1B66C+/0Teib+UVElsqdsN+48venDCQk0OvbG0HGIllkfM8/NcQyrAuYDex0xjtMp
JRJDqMM1OHpA5rMmpImHFMjM0DBHK3LOiO4Ihatldw4QYTR0HAvC5pZBGuRx1HgregugYj+oTq4w
/JTrj56JLbz34ZDjEki/1pPRX1towEP3tKE0S5D/V3D7VPv0QjrI2sjsYJGBXEdnYZePDbiIgXHv
eTlY/ih2GNFZyZh4gTuML5PD0X/Mi8m6EfdDegaEHfSlrUVlrXS5YdLIBcyKgabyMFrSh1IXJsBs
cRyO+aCVmevrceYEa25NBvuBkyrA5ktiF8ghC+PyoK0rIPZTpwBi2tiMpRQum32Zs87zQoQCCRDz
TiUycHBHJZLgRxMEdtXUkf2+7QD10uu2cTU8YSRZNQjDOSxcSAwedXZqEzw5eoqkOlhIivM94+dW
Fdf/n8rNddWGAWMM0+ljqEdvadnx1uClr/2/B8egZ7hFKkuj3kOjTMfzDm9AywfAwF6GSwmz84zf
winwcbCjDeftbOzKsHMPSmRMesPR8Z3DIygCEk+cgMP5X/VsKfaOiGbyDVvXHzqnHD4Yfari/K9v
pxPzC+/PJ+Sp8fIq5VemfPzFmzAvOGoA84dPFOrzfd4z08nETUjKiarnSyJSxuxcurNcX65UlaZz
qqTc1mDhVee8nGbKzxNF2COi1Me8UI6ENQg0UL6qeoBkw5rJm4ZmXQn3RUuxfe7YUY7qnUNcVR0y
VmyolhNvXvF9IjU7MrBt1z2HL7XFE2FPF9fCWdIQkUFpesJu0U3RHSeSHfhCZeEhf8bWXqOOWxEE
e2dm3hc5lNiAUgdsAU81dnf8KQwSKDp3vgweWCrYdJcpVyhtVKznbBT1HaHE7zeMQhld6CHpAdpi
SjsCFn80hCKcxKqmKS6Pd3193ZLHTqjoGvN9QTfeT4J0clhP83mBV7wcBbqiiRAQRVPm3NvPQxb4
bKqwHR2R7ZL2mHOe8D0wmVjZ3rWavj4IdAmAffIeBXGFlK+rqosk20jh4UWKA49EfmvKza7kC9mi
giHPNBOP6XaUSiFfzF60MKWSoIMQ2fkiRzCw+WPHhiiDi2zeawF94ZflCI40tr4JOdcIY0ZODJQt
of//LVy6BlL4jAJ4/HE9tk8MQWf6TYWzJ2u4e4AMeVfH5NE4bmV97aDxee0LZ8w525FklITCFWtQ
Go4ESyFUb5RlGA4+q4oCqyJrqKCfqpDznPZvjVMsjf8IBHCTs/KMYMk/vJewVn/fNa0qPb/XSucl
QCxXQGsf1BCkPkWoj+JAGcySEQ112agp6OJRrhLMM+wz8toVxKQZj5ufzmZDAZgCFucO71YDPIJF
ZtOmD9yfB8XlDl9iJpOqoplpIExxVjIQZGerYgIHdX0JMndSlvO5fJHV6uug3VEbeDCtXk/v9/X0
IMVs/cZk1aN92tj0/8uIvfG4EqIrQae2PACz8nTn3mGn+lQ9nSI5/xkQ+sV58PhMHkP6ZlojDZ+H
mDpO3l9TTZs5/uiqTV6af5qWjE7Yvg4k6SzULEApFFRJn/UTaYUnY6KlSMehnMxKQDeI76CBLtwt
iqQT+urLfUyvpOTDuXATpRmbkS+kEoV5ogmp+zlzPAZ3/GfM+QKqG7xxSdc1RwKOAmtUh9MSqthP
uWZb+czBfASOU6KDKRAj7UidJ722AJo9gkN/uXyZd3dJLlWRZxintndN5tKVIP2hcC7890iE0xJ2
AlD4cbF5Sv37FlV4r1kK5QSc7vvS6L5fc8ufWZqpGsSR9TDab+k3OQomaFd6df10geRhL3NLB5gX
mAD7IJdHlebH02ItJ/pCD68coJv3PDh4Xyqgs3xhHsnxhQm9rTrxpsTlLb081rUyKXItwJ0ZLruG
T3YrhhWQXmiWe6RXplW7d8uwpLTzuv5q1ouUUjb1z7PghVDe2SBoBwGnkGxf6ZmB1lFQy6sL60p3
TU4OhYL5ST54edJZp7Y+I9gwDVoFWq4e3MofAzLYSp8yweuNtogwo+zYgHmxBEgTanWwxXouS71W
pRlRFBlyB5C3r9Ubp+ZCLkOeyTPBZEHdNgjF/m1P4hBdavYImlMqq5NrhWDH+L7Wa/+mx3pNZZyB
QhooCY7GXA9PtLZ6RAMrq1nm6lvbzcyqT69BQfWBSLjDGChKe6YKw+Pq1DW2/jq3j3a9WVzqa+Dj
LgDq+LGU0KM2xqvdJl1nMEbGEB5GVVRvdiCuoB+vsTn9F5RDx3Yc6Cdy5GgV+yoprujkp/gdYxN3
uizWeSzo7ds3RztmtgoXwVa9cZWMQkHxCMT3z8XQXkkocmOIi7jxQzeq4moKNItZSEFHLEYscm8f
tosKnhe333xyS/f9zocIPP7zeGYb5FiRYziounuyOQVD7nY/miz5+HFjHkmMjXUix9UMqyOsJJoR
FPpqRa0bD4JjsgcH1Ax1kFPKX4CS8kMkBcJ7+UAyB9BcqnwRL5b5D/LODjDGUnJ42Yxc1ovLJzTY
P1yPTIyrztrWd3y0o/H8GAW7i93e3khhXT8Ynm1HRDpLUeyx92fk/hCBzSjgO1Cd8ES5Q1TdG5m+
KRIWdfFk7m9pCE9QcQgt8yht5ANJ7nf7CpGuIhLtIFCB0CtlbmCvmTqLROd2R0QDUzDWAQx8Te9X
i6FAN9dUKyCsoVhHZmGOfb/dOuXBkRbyGSqKXf2K0FU+NR1xXaMhSsmyQnZujEhXL62uMhdvJVrT
K2HlzKiq5owfuLxGNuL3LNeBrz1VLd3sdQOJChO9zn/vEGFgWLyr6xW9RexaoWsoAsV7bQTsA8RO
IkrC4zvAe2v8B5NRO4qIfkMHtFow3AFY9zGD9vIoe2gc1FCsgBo7JVO/SRYlSSBLHoG+CH9KFAzc
siUA8HNnY0d65rx2SHvg71JNX3ELKWl7dcfkSCd6y/MkCtGRBkBwRSpMkFefFP8DV3dupoVgO0u6
umjK5zabgekdDXRB6EjnBYrHd3e8SF4ODSpO2IJy9P2q+wFBAGcIdbc3Z05a2yVdOJwetv7kVIPW
bxlMHf4AZdG5M9Ts2kwMjy+g710z66Y6u2qdo44tmFMyk6wKLRGW+8BhrDveYbUdFWqYa2eeeaWD
lFw/MITs8m/Gmvp/woiNgT+GIG1yU0aN0iEowr4C8GMcBJ8Z0O+lcnuQ09aCI+z39XsPvKSOTJRs
ZebB2UtEPr1KpZY9gzm0n9PnHWTi63eqevksD4uJVgZqoyYA9BNjx8kervx9ZNCrLzzh/80t6n6O
Rv9ZNpbRI/MicBfSePniW7kdLuSIwMBwrdKi6/8aTT4wGPDckhOG59ynAkE1U7B/xNEZObkVXMHo
EAZe3Ci9m6Xg+sIjoO+gPLYmrOn2bpUTBItaJZwl9QhGJ+lNOxBFoQAbBPDMyuX3w/mbCMilRTIk
+OcjCZau+gYTLnk7xBTjSb99WWApeLTAzUtnUwZYxZFQUMRvqSdLpSjJChCh+ppukxSJGtsYW2dU
tysUN47fLxw0ww8LUlV1BAI0NG74wXk+Lbii3YQp3kjomz0OoItKJRkwpiMB96EhjBITVs+De7UN
QP2N7h3XLUYw1zBHbOWf5CJIcsQjWH2ERykfPmi5dGUIAW2v09IdOFuXV2bGaSuOd6rOhHZ4CiNA
FoVteDGkUUWPIWVcnBcdGfK4Cn6remj9QivLabwJcHK4pw/s0824E56AVNIN/RtvrrAdgcL4pUYt
XnXFBeVt04a6Ef1p+Bp6FLC7WUq7kz+ujmTIq1DipC5vZorfOwKncV/+dEKf19OryC4vZH951/O/
8Oldo5h0hY8ppqTJSRGCUpNBAII7qXKex5oX/Fh+N3Z52pPVPYYgyXp22gcQAQd1UKi41iD03hs7
jkLVNmEkmBqurM7FjA3N8W/3HK1ubkccu3WUMPDdaK2Cm313EkiR4c5jGDK6+wJq03cdkr/2xnPH
E835HRlRFiJpTqAb/QHZrFNcmex629seNa2PvDSb9yo/jUAmrr9ijwxBjjyJI2UDzomzRaiAYorT
g2eeEH85kDs1PYiERlTd3wB/wB3ZFs+cLl9KHe7ZWSSolrBJawRPu0ln+7pddKsc/UACq0gSCREW
PTYDqA8klt217lIYmdZGF9j0flOI1Y+eVmONo6HYJoVu/pKLJslQegfyxP8+1EAUxkMpopHYyaru
ACYY1Kt1WAajXT5Iie9cggK2Iqx1gVLfCME52L0uin9g552Ud55G+HGX0tOgrXu873gkyOCNGLKi
qtVwCaE9W+OupeirtoP8xRzQ1CblEm0oonwDClvLfYG9Q/aNzSgn9JgvD45uARZq3P64fVNo6GyQ
369Az54GVmG6wyYFNzdLY4IbfRDXQIrbWB8NgpVjAvxd1e7wZ6quKxEvun4G/6TH6mywS3jiBDDq
IqHUrrqcyRN3pFE13rY30EKxpuW/p8gDts9AJV4jdJX2wEfco7t/vXFTaOmZMJf0giasvhx+ZpHD
h+x8WLoMMMu42fq/QAPRPwCOpGYa+xgF8OkJ/9rB9vOHR+epsQIsQHuymFQNW8IWETrLtXC0WRcW
FcQqIIJJar8T3rXOycMDJW47dIcGL82v1e9GVyFC03tFQIj1UZzV2V27HEbZp6/SrKRD3vAZZ9pm
z7cyw6QTovh6n0q7gYmOKZYx9B3B+MPZ0WekgUZzRDFJf1zRGLztX+lBqKXdZxFuSrIQ3HPaqaFe
yCvZk0+7ogCKgvVHWJQ2PgHbEask7aIaEVFsdMhyn490eW6PZ4fm7aMOntL0fQr1aXnULkhFipfX
at6phF+mBnFnulJ37D56YJteovJwZMOdbpQQM0z2hQT3utrwrhINtc+1aBvdbdocI2OgpkufBiYZ
ZxQrkY4OBzpkDPQHjB1tcXw/uVKEsdjMhCxVVTq+K22mWc7PbJifR8zdYhh9SQNlAGE0wIl98TkP
w314/Nw7LzsJKMmT2FW5rNiFsxzbUDBW2a/gYR63UNWwPMzkzLMVPUb2y2c39BP2EvB0toXjHmJ6
VcHf9ihLLpJAGay7pYk3x7OIoq+QPSNC5Bkjf2Uk/KWN7SALkO4EppvubuiPyodRQup2L0uGo7eO
vs/9QoBZsLq98SDOrNmDqHnLEnfi6JfRBYWKgbCUUeQJ8ucMGgc0SNfUqWTVd7CBO2CYanjo/uF/
9u+Sa/HJvXwTR/0OZIOfQa5zNx7F2pBzr0yO9XjsbDB6t0bwVoQe2rp8z3uBEuFvgDCVqhygLBOt
cOK08q76htwLztwHwDvd+5pi1qQISEHJSdbBoX7jwZBx6n8Elu6XgGAdkSWAzdukqzCpWjLs8C6v
np3mU141aPTVgOeQW37QyOoZeiroUM0z2Vn/NXKEKw7pV/zopHBUSYIXhHPhxOvk/DMrhTHRjN7o
gKQmmhJ0mTRVIhbKWIhRZetIHjuGXV9n+z62DDWBCFW/X6RUr9DThkiBtRAOsoRaHJ/HNW0UqZDj
in9sKlVX52yrPBiw1mgYDz85AJLWkRZNgQs29R3ByqZGXzV6L1WFxUO0T0qP/rXgxMgyTgH8ADaK
vg6y/6XtXckwG2mDlENqa7J755kolL2hcGZipRg6yVSMy4YBD/o6m1MK+s2ezQs+SYkAuIf9m2yx
XgYytWIRmd+cU8uBVA0BhrEBjTWYyFzRuO9zHFZBqtjFRNDxyGdNoz2ELV8t0uF9G0caZW9dyczY
xBdYTTVpE7tXx7yLtYksUerzkGyLx7GKdyyi3PiUNx11Le5vnQ1TOOYMZRti2zNoY3BY/UGOnPbe
ne3rS6D4VAuFVjGtLchqQARwIwWmoRAdopDPhhlLpNTKb848FEszqIKdRSGdvHOkY1OxltV7KczY
Xkj7dME2K11o9tNGV2m8em68JBIU+x554DBHveFlwHpHoHq8xftyPDTAT4DGHtwrLxXPmILRkpm2
8gnhX4n9dEHsridxEZiDHaWkpRrbNpXY/6fu2VBi4TQpQ4TW3KYSrbRF7JfRsYn5da+JMxH9ky5z
e4JhOjNmrXajouU/LSvfN7unRGCUlqLqZ4zIZxXbEuXu2/8ISSRqsecNyarLXm9VYbVlKBPjdJYp
7tplLfqshGIwOOvJV28+EK22pbMKdhSME0yrv27Xxk19ESXb9xRIHG+kSEpqBolZWTTcGe3sdw8r
nk8VP+UpBcpFKayW8XAykxcGjnX8e2OQxEXoVTN3EkzZikU9Umx1kN+ZGbijGTq7NyUK8+8ZTtmT
ASkqOa9ahpkgQtiyi7scAWqpZ0E+sUp/edZdvgNDG8gN5uNmqxCNWmyDl2Wr1YcsCr4YAEN5b2Un
smQ75/SFUCj9zraA6objEyC5m6SNULHci+UMeKBmQ3QSMP8Extb0JidHpsLI1AKyIbsqhwLzbYHL
TOV403Qt5WX5Gi+7U2wowAFkSH6QZwpIiHcx2KPbmK/e72SjBbgH8E26GNbCYKrj7nGk6N42eugW
MyLFTaBJJ8bLExBUVjRQt5UsaqLlyJh7EdmFtGN8lXmAZa+nKAxTizR+YOQc86Sg+sDwFW7Sr7sg
nNNOYan9u7hKJzZnqb9woMF6gkxx3P+DVAFHckYQnANQ76Dw6+9owQUMWX+tdehzsFDM+/FAE8eM
0iWAn/rbOFVF+XWXYfu0mA3bWpCxJ8+qNJpgMtAAfZ1qHURpZcJ9bMSRP0xy3GCwdrpzRLYdv8q8
9sm32m4U3ZOPng/dhFyD6VZe3acaLLHycDpQeplLUOIjuv3VhTL+vFuLP4aMz62y5kA+jo6yxHBt
0hFEiPp3XXzgh+cWcjFUy/TaV3uoZ3a6YRHu1p6d9aDd19TnzeCVcCNwMNfGEv4w59xlLO81SnJB
Rfle1ZJsdN49OJoQGcQDkBy0oXg6V1seYNp72O1z0uPJn7E2DWbUNvqBRknSFMotTHOXe7LhgEuH
s8jB/PXJKlGLIxjmeqRubkvcvUMfqiOUrM1OfGIsOwb5gyPyXRdVEtSNfKyOBElXphFNbQCZ8rKM
gpE0Yy2ZxgFZgenxghzA+egnWewtnlaes/+TkwZKAzG6xYWU0zKb9RPP//PfjV5p+/isGGn1nT43
7U0suGidwxnR1AQLkIZKBuE8STBmDhg5drensjd1u7N6VNP4UInF0wq4MS0FIdtP6ZQxB3fQpqTM
Sjp0SrdKnVB61Uu0eVEdpWT7tDdVzEK+nJsHP3r0aw75IVqbMJNKRCu7SawtjjvUXuatqFG27s0n
zGk8daugPNqmzqj5X3peAJwlBVpTUfDSrDUFlgfRtZQC0lB1X1Z66CYJzY23ThgcGftu2UQih1FL
bUde4PEHgy/CpLchMpmUGW1+tlX2l6zZNC22tdJyORpva58BQEBIA6WEgfDOW9r+d7WfwBNxAskG
BcIQkc9STdz86yU4dpSBcIINeCPBJE6KzWkcVqmH7LY2z9U2FWtXwJyCyb1u6r+SlL8eqkSWcWK6
1lzzOR9LrSz3E0cEilcYPG79AmxCCdZUUH3jsVvLj8HreSs7ANpX7raDXL+pfEJwkekkm8+sbD6F
AI1fEBRE0itW9Di4NXsMsTY7kQ+NSU/NFAgM/TOixeD+Yg5aYV+Z+LN7L56gh4sDO6UET2USjRu6
HK+Ama8WNZkVfHAscAMtHIcF5mSjOxE8fYO+D4harYM+YQDD0g4vm7NlQ5gLuPka2BB1Ywxr2ly7
0jyDzl2Cn1f50fHVSNgL3NMZLuyBEZkUiVEnl2hSdVgEob5Rw+WqKNkQvutgOcuXMZRRjBgXl1yi
jr/qYommebmh8OWbtw5hwaC11+QBIRPbxfpuKhka6drvwe30/HFkMdjsTvD8ldyVtOOII37YGLVn
14ppONQqzW+hMIaUe8TBhn+jO+D7Sx4axLmbZZSQDMACO2wHzdHk0jroIbDJmhycAXP39dkS3D/K
wLN7AbZSkE0Mv04jMof0Bk9Bo3sLu+ugx4Ldd9Op40RIGtGJ8Hoa5GAXfpxg2vMRa0FA5MQRFE+l
Z5ty8Ie14yvejYlP7VnAq4/WJ2FHHQLPOU6AA7Ouh7sh3rI7G5Sob7C7wD/Ypt98kJ8LXhbujse/
nGG0K4z+wXRG4ZLhtwV/0bHhXONBm/hb0dXpDQPtmfch/EcSRYr7cuQJlNuEUEMR993X04M7Wf13
a6BJ4hO9MX0915GwfqF+2h6tOyAJmxsmAwx09XCl7a3RwTkhdPs5WyIrEkgPaYddWoZAT+oGCmGc
Eo+pNR1SHLkH9WjWXpGUU1jnnnIzkbcq7x3JYT7ZHQKaON38rIkD9RFas1RJU6l52X/Dn34WT8zv
rSSQoWTh3SsUo3z3ltFaxbmrpPbZ1uLq0qQuPcEWM2DYie0K9whe9YRPYj9dalXY9Gjguw3T9sr4
uDVaN9fTGnh8U2lXv3DsJeP8Tc6RGyJwKMGFRyKVRWjGWxC6B4WbDB9tZQxqm0yD6bcS36MvsgsL
+2rMz3GvSpwEEoMzDTlpjSSXYw+aVjx8M/3tVaXBqatbF6iFz25r6/glaMvez5IeSqPmicNdJHjw
NDFsle7QeYgGpgqcOFUxkAqUPh4ypoRpTkYAuc2juRs9lldzHLivP9ltrQ1xc1/kdXk9L+2a92Sk
TFhxThXcvyTyeJHo5CWqiVqT4FMBWSjsASkc0ZIDMq+mR0wWp4M+QAOIi1pYcONEsziM2zB8/4Uz
EbOIFeRPz7yRd9MBVUYJewofkBkKh6vLMK6IXeglL1PE5fEQnrsFsgz0PFJfGMGLGlJyQuApbIfG
RhGSASfhIz2XsyyG2axBK/en6HokzA0iNs74Y+xncb2zGR5NdpAmWsJArPJWSxQWbw070DPfv/Cv
wcKIUdhThc2vAyVvAloKOmt+X8qGe1nz+d5ztP3qxZ8ECUiJ0waM6bvCdA1T6Yc+RsJCHrYzvs8d
Fa8frlEVdox1hDex2dnFxbgismTBaUlwtqwAljNVpAqZGJbbnaCOrfXyp5UI8p3W3KQIuISZ3C9t
UaR3GMC0dCVzTxEbg3VNKXQgHWGIiPOgFBx5P/e8pbDQOCKFXMIgbUXFlDjJEc9+KKerCHX2fZCO
PwjteidOoKHYZzFHjSk3GmhJspJFPXModxU4d6c0OuI1hG33qpBB3PFDjzkMGFsQLipSlUa4FKIg
ZGczSX91qNFiB9vrDPu5DamQV7vXB+UHnS0bc4YJV2q7QuCTBt+JmWfQuNyBe6SGn1ygTZEVgDoi
VS//cujfz5czbcmAI8PlWaxR0wjXjnfFgtabgovXoZITsiF/KiRdAJGR7jjhoBcwcNXsVn0WMQZm
uq5JyePM4AR8ptc3ou91vOikx9CjE6y0pfkmz2kROyUT7jH1Q1UaS0nIjPAbwpavwwKN27mZa3Q7
/K558ViIXXDCq9zVRd6ZYSEVNGMIj+LpM03hiHN++eptEifwL9mHqQdGR9w/Tz1cD0dpoERAcF30
nXwGiMxmcSrGfNN9ZFqlMslEPgN4UhPtU2mi6lAZ1bee/JDIKk1blC/EbNwZiIYplpImPsTYVyVA
RC/AM7oLj36uean/EnIa6YiPhoE0+2PcGpFtbl7kba9D+yAVPyy9ahSz7bWEJzpyGKilVzQHmayc
RuxBdlvf1DV1lvT5C0VR8bDXM0nmuFOlB+HEhi3ETOVWjmAsQvLtQpiI2k9p+WQ6qnhXZZ5kXulc
lXWf82fQvB2ak5PhPtTfTBv9/Pdu/a3oMnE62jq6HcG4r2obmt321MEpYzNvGTASH2gZJr7ITknm
fLcu/hJ58AUM3qb9C+NZ5UWrupKeuefIO0hQCF7wz2Kqxp+GmPLHoH6QOi7hNIKf5OUEc5V0UwYu
YvvofQe7E8hk9dfAuMYjBMA/q5s8uVzRIaMWsvs9P+8q/iqE9XgenP7i9f+aVp8Khy+WeVIT+j+u
k8O1XOE6yScXC9MGyHEOJJGhVt6Do5ABLeh3LxaQr3jpwLWox93h0xlqfXnkSdMFrPbAOaH04Gn3
++ZQOpIBqkKHl+V8kL7s4iUV/+8j6hoxzaRFQi1xVbOVPDfkKju9GKLY1HFzLAmOeFKzE9cfOiZN
AGnXHdhDkM5WmItVlmgZGd+nybKVaH2Vs6WHtJkHuQ1EH0KGmCC6ZjaGZ5/fCKlBcwW9GkDtVh9y
/z8ptf9OWjMrMop63dfD4dar0N8lrT7x2R/jk4oYOT4vzRU7PTyOoedKmeNTYN1e7vjLxGaXFRNu
fCevEklwUM2fCQ8uzSkHxbsJPMB9fNZ01ltMtW+8G3cd8fUJIkxsxg1FDgmCGsROTg7RI6lfw5Xe
kcvK5TxtArlOmJiYL8OvUn53GAQpwEpeLN0OLHhgeOw1rCWLlWqI+8YmUWot5L+2xCDDdOd6Ez6j
1+lA0MSvTVnWVwvrQ+vmkvYDsCz+0JDFKvCuDSh5IEjG840iCVq7v9XqTeTbdie04E6GVps5mIZn
HcTiwXilXxBhpu1Ft5ZBUZ1Z1dO/WUBcqdEgAx/n2lXRs7ebZZ5DZrbjFLIruLtYxsvhsCJTQn/x
NTBjGlee/abu9bMAUolbOqIp9ZJ5pZBpTAl5KYuqPF7SVzCseolOG5ZaCKDAZOiWvTZSZ6E1zXCC
WmSDcjR0vMXhHdJySaGqjaLlbH5ETMmPsGmyAEKU97q1XDXSc86tzxmYP5vYWfxTc+O/9n80I1ms
ivVvbv5uU4MkX1jvbSKJ17Ql8Z+JvuFFc4MIyMA0xWsF6ahzuEB+Fub7VWdAPTsQdWUllINYWraU
aer5os9ZOg4ubOeVqJ/c9eLbT6rm0WpmMTq7OqVeK8sLpaOuG/vnAr580r98oMQYUOez7eDEjCa7
okRUDlhhhMsZ9oGclXNsibTwhNBfXV9issvUconKB2jW3X6Sti+2uFbKCtR+C+fCc8tsPV48I2+5
9AoNYA2E9nLx28T9iWfhR+yfkXUunndtAeXCbv90QDdf163DRP+oY/4kBRMAIr7tXqWY/A2P2jIF
6vADp1LGuReigtyAyFWUGeZavoSPuHrGgFg+BPexDrFUubOsIkwEzPbQ+ef19yocYOHufWHpJ5a7
UoqTWroeD2ehxSRKAjNTs9gk02yBN3M7O0HQv/EuSD0iyBt388mr4Beq0Ycy8STDKU1tn8/6rOry
uCHEX44pIB+eNBvVl1dgBM1E7/UCwW9D7sJD8sCs1d7z/jAD6Z1ojK8tgTUeEpD4P3zsRVlNtjDD
nVbPuQLPnvpzYEB2/EtbgLj2QS8eWqbXT86r5G3lLLAEVk4uE6Vj2Y4wbUWjI3DSqSC6rSaq8s4n
Vg4OSd1E2bnOS45DvPAoNKVh0uAWh4dwruF6XhMOY+/v8fpIfggWPYtiGZ09cQPew+brOidKihA6
c6xDCOOAcYZU9n/Hinoe+sf9gWCzWx/N2tO3KfKROCmben9zp/jOgO5vKfjJI1jQPj/LrCUkeQMH
dYnqin803ppxpFviWBlUE89v0zUOBDCXbk15NK9vzu+rDnNN4yFI66s8ndzuyBDMgNP2kt2ym+aO
Ivzsj8ujnnqOO3BTiSZFCP8cs9r0nP6uxwTHhHGPkITxzW46ZT+ACXpl0Ww4mFbl5o/o+M3u3tpD
KOL3qI8DjlJpThANF2b0mRM5zAJ6xf4BVDRWhoVk26MS1ieupldyhpir5WNuUy02+hm5MVKVRdoe
mjuXniG1M4QNFaH+/p26iYEWhIsJhv5oKpneATT021dot71b7KjOsAG5nVoTL/wlwbFD3r0tS3NW
r2iXF+Udw6Mw9pSWQbyLDqBTARG/QXXh/uFiR/BL0NHHmjZKhzq5dy60amsn52FfyB/HDdXd1/Qp
PEsXbSwLsVutS4MZOnCT4SQkPF5ILc8DwCqx8OcJ6zz2gIoyzrkuMjji1YO+vbpxdO7YEFaH9kv9
59BEfMw/u5e8uv3LqN2WcqbDr6MWBPvIrq7oYNtzqW7R1Vm19HpURdGdST+0GPCY2i0gADsJWhit
67wHz9b8s7cSjamtvffkcppxSqV1nQF5ppUMNna5xs7/zlgVibf1lqz/6KU4qXkfoBZCwpB/flOM
T/pY7aCQJo/8CBTGlJKW2hOnijf6615pMyeQB5URE1fJeAn0QfIDhkCvIgzby0ra/gH9zqbOYUMY
hv/8DWteEeQn21l6WENmRwO8vFC75QYzS7iDwyT8IM8jpmP4AFSBVa2PRUkA/mdh7XQv3oDkntsk
cK/4lZwWDh176+ZYxeW5GdNlUkRm9iS/X77Zl5P4FpaXo85xNSOYwwqpj5XANfVqWfb5azYph8rv
QxQGGZnVhADLPz63XtPA4rkFDBEmuJehSj4OfvvltnSc95JAt238cLQqqNBsDwOlvBxjL5JMkqv5
Mlm6PtSaiWkiACFDBcJOCJGJTb5lbB4gNxCE0o2ZdsMtkYSRsmaKTFEQ2PCl8JV+LCmEERqLGGJs
reagyDrW8h0r6wp0QImXwWqKNTDcAQIB3U4YPzvMLRHITpeMMeoEMDbgChVa9O6iInCUCiPjFoCg
CkHAZyJnnQz3JMHxJlx6h3w1UGhgMs+3FTFc0GnMVsXD8dWA47g4p8c8McrJlix19nZ3DqRLNX/J
qDY8YIwIcrKwdxFV6b099Pw2J9hqVBfdAz3LUWq5DVFdDJ5eYhpwi/c6jQG1PamOfIJxORhBqXMU
YcBoBrTUKKmBXTfkXlVOTY45FQO6f37Ypmz01sygCA3XMjF4kkgZgelbM7Zzwyxsfhp5g3H02MtW
odMmfpAjyxfous7gg8C64J+3paOZYz43lxg6CFEG2VQFxAzUBCCFmYg8pW8QX0QhXHbvhXdFW6rO
4Wnfa6ewS0LFeBMwSfZd7pCghDjevEeYAZ2TneBC3yICb/Cqs578rOLd+Up38U+Z3oFhECkDuJnS
mtQtwrXg1ayahF3OuhpZLSOBWe39AhDoR23/7kkC0CDu55ztMYAolZBt4PerR0ZdN6/VWYZPrKYl
XbZPOzHk+0JVhSNoSndpDr21uvvMqPd44R60E4fUnNLavsNUqIySpeIipuJbwZg9haekOA7DSZAA
HOgosfm+lFVhfk+n8zfyfTrDxgSwH4jtGmeZPmKDCmdg04Y833wBynMo2lixCFdCi3JVuhank7ZE
3lmKPoRerb50jgDRwIVv4vDdKzA3sxwkKYvBSy7hJxcTPqGpMx/3wU3wGzD8HbRBKfCKKJX6FUao
QGeBW1rSiWqqjbR+IevKR/N0soBgcA6J3NqBcYLHF0GkrqWq9NuVY0aNMwF5foIUH3FmaRhlCvHn
KBlpnGcRYDAkLzsm0F//5fJrFup+3slxOCrvsGmxSfUAAfsSn1fyVmiWn0xv9sI4e1n9kQSeonyp
x1aWLXONxkj3kw0Yj8oQLfUhcoIJj0LsRBO1sLUv4MsPBH/2XfUViYNw/1YzHWQ9NanFYT6Y10L5
RinymRC6tkCp+Eb0j5yEyWkzDT46rCF1BOqeeUaBmnUu1wAlgAyBQc23lDTjSYS2icabnEbdzhwi
jUqDhY+dvObJveSlk5lKu6G9MEjycz1Zl6CN+Se31WT/WrkV2E6fTpjpLYNTLDg/ksfCR6tW2r4K
61j6oupicyM7EQgz/QjnUXf4Q44a42f59QSnsuvcrxV7+h061TdbLzOC2EYPfZIFrld2TZ1NI4UJ
6oLRdydQRw+Ev5hZiN3wGubn61nqXqsIT1ruxZDc+e3mFAixfx3VvU8Dd9hN0a5hKNfIPUeU+vSb
3tW8R0PVqR6g6hf9HKHzgwEGDhN28FXxs1AJ2JqDjeipFVxCRqfJ3Z/MkgoVvubdo+Vj7r4FItz/
PYPn75a/mrF0IlIN7J3rOPrvmBKhwoqr24p1TKu/RbK16zNGKKRZV3cUUnO7riMBHieGmLdHJxaO
n2BgQgghExdXQcWgNO8GbzLA3n/0NRrwIh0q77vidCI5zUsTIBLRXE9Imm3/U2CcsV5LVXj1qPs/
zZgJeCIjPEKHaTqKcMQjzB0ASTf5CaXNNS/3cqQ5rJJxJfEQmVjGp7+Mm2El6QnxQjjjbHugY9MI
JYUkyN97ElryPIJjtyX/EhufY9V2FnKjXxI4efVhpGhKdIbbyHi9tEWld9dIuYRz2ACRmFecSqZp
sLqKyPk++5zqdGbX6H5YgYfBGcsqcY0pP60Fn3G8612KwBadmuWdS7xlGfGaTp2Q7Lz+OsW77eTN
AvLntdrGXg6YbgHOop6vjITf3d/HVSKC1NYLLNgaXjEGcqfUiUhLxRFE8kEdi6m2+2MBMW7V2JWX
azKyW5To3EIIp4d3Vxn4Q3e7Yzj4YX7c28ke3HDa3q8ouoGmE7DyLFdHbyIPO+xT62bXNBrKkfPP
5ZHDkhjXMZI0G8t/zzijGhYkqZGiyTYF6AuVxD/pMEWLJj/qn6+38bLsSYefSlZKXB/HZZHQKhx8
jpJvmu3UlkPz48YTeKF+pdysz++aQaKens9dMny7V+x1wun+f3/3QbG7BhZEte1OgU8rJpUj5Vv/
spZMC6Ah8CPwjJeJwLWQqpSs9mhhNbSpSGdKXN5eJcabZZ/PHMwqDdX81jdKCV/2cDmwRH4BKO8r
03/s9cfNhXcBaxur6B8RhqXkc5GlncSZE1C6hqUFFjL8JG757757DkCz9IbJbb/7UYTcKrl+oXJy
RFHUA1bMedW+/duQI7DhyoKW/PRs1CvmeWmg5jnr4uUWizxJKOU5zsJwxP16gVn2ZYbtwLbtmSKK
+QKr5+EHy3PcxmkfUIm1w48sv42yXtv6CL9cYo2f2qJSrTOibE9Y2ZnTFpW4vGdU1A3eNE2jUgVP
yLNud5V2+PL35eIVe7FxhlOgz+CcCoPfZJAjLDDZJK6nRCRpEfwU7T8bT+Bn3XOyEkHGMYqxM3KB
jcLRkbtf/1xIPMJkF9y/4gvg1ut1TF6HB+zRhgRNSqt8m5VII81bBHS0aW6EaSYy/juZsqw6n0oe
Aih8eFAqlatYyftEROrkBXfbEokgIBdQTq2lrxKBLwa6HWRM5n9zYZJR7JSyzaBb2JPE8sQRNzSK
xOCTRgMlfA4yjTwJBU1auPXr/ssydoB4qhyP9TgtpD9NiNGT16W7tvN3nr7jTUCdXBmrNjmqy5Or
Gre0L5vx6AQWKB0+zmPDwJQ5TdD6Bb+gFuztHo9lCs/tQHCpAN8AflAAEQhBgRRM64407zxS3pU5
EnbkH2xz7gaxubXhlL1pjw1Z3yMFkZ9LJaj2oi/5Ddxwjh4Q5k4alPKeXWQ16aRuyoveWjaC7rn9
Yvzlf8pS+FGlz9sjz3vFwGxbMHfhHzJWFpZ+F8hSi3044jzYk/hBsoYNdjsRe+mpE4p2rDRWuciK
ZLqI1r+9v7X1nIXh/40Na1K8lFgyav33pKJFeIvtGCPfsQFlaQ5q7wvyfPM8XESsOd0OAzS0RX9R
PYmRu31PF+8ZeXBH8KBglw4EolqggrEUba08ZDwMQJZ0WWo60FnPVVZfVlTtxf8Wt0BfNXsD4kcl
p14dpRErKkvlszwgeX60bwIm4g99SdDZstNc4+Plbni54HGvWDT3GI8C7x4EquiZeDXc3yHRXJVH
P/ZC/eJKA1s1cOtu95ZPnjRI66IFWMTopAu5Bf37XPqbdhbE6iWbn3AmzH+YoQt95rz3EQvKTmsz
KQmlIgo7k2ZbfKYWIbHhi8rW+lGmBPkuxR8lOdr0ZxKa8fXW/xK1AarKPxlbeCp6mQvzQ0G8c9Eo
lMx0N5fOVWJ6I1cDEMBLlU29GbMtHBasWbr235EujutMVysyKFftsvweokwuCH9jiV7i82za9e6x
lAk1AwvqMbBHZuuzx0xcSVfK4fWRPyEWJM2Tzk6tvgZ/Qy2sqfMcNXaY+oWGpdJK50pW1pJe2Q8O
Ps1UbLnDPVXiARcTrtjXkHA42by1/CugJxwseQQrjCLcFEiK9GPkzmRfvvXR8rqTp5Uf0PRRB2yO
rceY4VyXsokQx/+eMfTx7jXdepXtYsSosYG7aB1TvII0sPzpr5/eCF0rQEq/q7Il6eDBsU+AF+lv
ZklE7smKQSLpuHLdr7EJSUSLNGnaGhbBiV5fu2AxDVf7q4i5FDI3lnqps3XzIiACwrx7Q+yodXZ/
OmVsn8P50lGNs7s3yaC5yOhHzWBIUHUmGbZMxhKNGjg7laJMSPhGI+lpOTVb9Ff6fA0FAhBG5CBq
RJ95lJahvDv1DCJw/a+v2bys+2FUVFhLxE+Vkehq4peyepKtbjRir+7wmojnMEz5BxEi3AfYa+/c
b+humz2ATyBKfRiDaus5R5kja1Sbl8/vH8ygCD3EK7QVcZ8zekehOCNkJz2DrBnkoJzLlp9psg0r
sFNsiUgxAEhB8nlTn4gjaI0tgx9YtQj33wM5Yps3INHuQq+ygDBPx+uozDpwwk16ejDlg5HIYnM8
+wjrtw/ZXKStF08mfoi0c1fOxonKUdlmZDsTU7R6VnrD3zcwrdPjlZWLp48NoTKe2heoJ+TX/jEi
xrvWxxzxLQn5aHSzRk/Z/gXvfiVcuylsqOzthJgpkRE5cksGHcXSwNZjzXGa3qMZv6Unp31lgHG2
SYv7y3NIYCS9bOSTeDJCQiM1TqPScef0mW0ZzeN804Bv7k6wwf2/T2VOIBInXMBdKTmW9Eyy5vne
shod0fz/OFm0qitGmC02663dNb1D0zd+P03Ugx4D1gyEvtgznlwSOJ8GYH5ZvbtbgyNd/AJcZ1sJ
De4+/GuVG+tKZq5pftFZB2Stfe08QfFLCW2wwZjQPO3+5b9QGYSDXIQzPumpr+SG4+HHOandXyhG
k3C32ZacYXOPB96Ox0U4dcVkRggaUR0hICg/ElreZz3E6O0Mluy5RlSgaxLFe+j3baHfDrizI5uH
DEBQePaJY6pALaVJkbA/q+Yz60pEuXhaeHkktySVlChTmWkmjaOHr0iQ2GuvtlE4cbzIU2NsB8/U
su7IQ5RxndWmaHknZy0OvpDsU1AEqXXKw5Ma8+xYncRZ+2JlkSOWkIWNbpvjgU7b+eYZ+qbdletu
uiTXLMqMy07/F+u4DPbS0rigzKLMgMaGXkVj6ZcCvMzfMr60dTxTUQ1AWKFNx/SVhS3VN3m0JqDm
9Wp622jpttcSBNttchsEi2nsXuNbNfv8EopWPevJKp3Hwo90kOdUr1nPxNZQ18lcPVJzFgrowsD6
8fv3csqLz/s9vQjI/Pmv5lWrq2YjlhfEJdp64KBgCntmyg9uhlOIbfD5Me99j9Hv3Nrcp0vgSrcM
apIvVS5E7GJ+kyvajcrE5JS3F6LN77vE/eNC6WcWNloggNRgQ8/gMYY7LBf2NGr/Zmu23QezjoEm
Qklr8j8MSoATF//8FrelxWANv8wlPV1oPm/jPzbbnkyKFptnHbu1g7yjqA/pUe0wdhPMAcHkdiR7
VfWsqWHqBJdNtYom8EDcr/Qh0MfNKZpHNjzdcEHFk2b+kCTIJDyKqM5UAHTmtUyBQrmpi9dKikj8
16hqjoJwPhVKrwUPvDFsyR5kVZMQomVbwrhOv32Yt002VAU1wh7psAPJ/6YAKi0avl6ODeiiHVVM
FInIllo3WpxW5x5rGY/fEq1AkzvjPHMs1JfpQTETgmI+pkA/3CUAHU+XsBHBaCvw4pXl3GEzgLlq
gXdwYITcXNTW+nyPDqFqBuqtTjTw9v1cGJF3JPKXcf3YbHq3PYC7Ky+W768N8zueolyoLQBYCVAn
VlnYMTu8+VVGyQoKgKFh/oz6e6R181B2hmfWGIf2miUbO2lVNeAPnRixXhkTQt20OEXfqrgmaRse
Qxk8ekamL0vZlRQ876NCuwj61p4SmMcfxOXhBncDxXLQ4ldTvU+0x8LDDXR31jeU+Iz/amKDKGbq
FyKI2IsAABLhgLa/mlLYnVDjUFwUGLrC4ePoXofl5l8vM23kWuM/gOy/LLv3ONYi2IRs9oJDOe61
pBKaYXGj5iElbVgNGIR9VWfcI+My4h+K47e2K9uUU4f7C1143thIH5Dd0aXtct7ciRU11fKbcWuK
sQIClyMrN6M1Vp7hBJ5TyvyESKnjPn5vZKtR3JPKBpBZvs2XEMEav7crjgUxp62ZzFDh5PKxqtSm
akLKLyosgdrYmshi+vjdeKxoFUvScLWZdRojMzJZdx2whj1cUcGWFyMwmDBS9HN9FeCdC4qGVOmA
jG1/IA8e7u4cS8rcLodS20y30NM9vIX4Sk4MIwtPLuPZcgWPUkEyJhN+YgvAQf67CwXpkqofQsmA
q2r0iQaZwJJrh5+vKH/Pn8aVG4tph2CHxUyWcIa1FQSyBtyjWtZ3jvtbgVnsTBxFI3oGsBMLPoH+
NqemuCMfN/Jr44uBO7Oq8sFHiNWoK2InfBAmAAfH2VfpO0dXL/rKnhKgcI6jntilrw46Q+yji7CF
KTNRbWbenIEuoZK/IUECiGGCDq6u1pRqfWk6S55GTp3R+ruxxV7uK7Pw+BYnaqE2uMBwuvBQJk08
ADSS7PUS57rBhy1I94uSX/UBPoBoYtdWml7LDKF8bI2CEX4jzn5yKFFM4YGpwfvfJmbRhkgXpSJs
2MG5WARqAyV6mvkO9gqgU6hs+buKRja1umJGLRBVqMu4n0mg8B05knCU3BQXuFoYa82we5+/foVA
J/EQMktNPtRoLWryEuH26AtaGBeHEVHTAqYY3cMIpZCD8yP0wwKNbTWfZpjM7mU0zbrGpAuBKLyu
yetmu0sEBB9+zOk7Ie8/Ma/VpusPdf1s+fXgeHeQ09leCVYBEgGxG20llqeZlk5oyudGo31FwkHx
Wh8beelwYcw0Y0m3WES35yPCcyPtrnounPvEKyiv3W+ALInUDPwnIfxn4eh7vhcvIEQGlfTmyR97
NVQfZeQ90702Sd7Pji86Pgf7XIBoTmoqAqiPHPnIp1OOmEGWZBDk4e55yRamJD4uc4cx8Q8M0qDQ
z0BTBphZcHs+YRjl+LATfNT2pO3Ky+JivoC+5rCuPL9rq4SVUbFA1frMIb1WmOlEXVkbNcrjGf3I
dV8sQZFsLowq5cKajdfyyEIW0r7NfVDk9xFuaDEjBYKHf4fzFbputGGD6TGy4M+y/DoEe2DU1Zrw
RIOFm+gIpKfO5DPLKTtKJQMYONaQaoDPjjLDauYOJ0HpiBflryQRUGwqbbbvoH8Z+FnCwq9JtZEU
0LrK8ZJI+/s3r2MoIQt4Cw3FgMkiusGtrnlL4WaV6PzzYmiWza5P1+x/rXfMfOyr/e3/IXpqpy8K
I/FbHDdy/JMLV0wDD8YUOjTlcI0seKY8iWA/gQVuVoAOh+k3dL9h0kJj5VGyBozEWYI3TJ2TvYLT
ZjloMO0BBOj6XOXCyso5pOVbQcVUGXXRb7upKmrNxsRIyoMLzGCeWiHrB2BYiFFFaBkP5Sgw4qvE
2piCy9nGxZz9lP7WcMZz9yPerbLe8MUwtSrRJMrueQ5/u5I7PYGWSkmmCXq0KnDHnnq58IlsQr8J
jvLuEyu9x0mo+QWGi4/g0gBo5m3T0f9F5h+gLW0ZOKYpnqoqHp+F1T/XbmfpbzW7wzTSt7icfGT5
vGu6O+i+/pR9LON8RhTguXiR9N13/LzRdyeOCK7BoasCbJOu9Z3R51H/BdR6+ZYSduUha7b85hKU
MY4xJ+hTKhfLYZtctkYCnnJaylJgprnZWicV6RAP1/I90+39erL8dLAmZia1MnR8FCsV0z5+E5WC
7GD0AjEXxvWWMdby3L5ts+k0ScfWShfqnQ+Hy64HEcoiW1/wfSxEmqgVcJPQVrydDUjFg7Hulvcg
jRih0sSywxiaZWdhgu+V4LD57f6GauWCHcyAHLpAjHNIzj2cSYo1AIX//oG9fsyhYozsUMuOtAMX
8jhiop6732Qo17vS3/CvKIqUoo9IrHhClc79nwCwEkJ4TPExoTJZ+eUk5w3Hw9mBx0VFgEXi3q+3
8Vn3dwsZWXAv4rUxVnK5kBlEIPzk1LYU2pK/hlSmTwXBrzLKn+JkAcCo1SpAx/aeFOsPOoeQu3lx
gyFeiD2ZvbJOgNiVjdbXGmn7VyR7FDRAoz6rMxgXfipFWE9zaUw6CE5nTmyCdYMx/FgoIOBD7mbw
yRaOX/wiR0hUUKDYJ36C3ZcKHMjTxOhCYs6GTt18d0akcpCtRxhFlwwnTKIs2AfbGZTuE6CgVuuh
N7Oba1kh9hDPZ2OIQteFW8Y6VOHcYZ/BisSYwAr7lDCrhgR9IBOv77qSPUwWKtsl67r/gERAAxBz
YvUqt46DoTtpXnAXsVg7iC6qjHwOsx0CwTAC1aQdkv9n2IkTJtsv0ILfgHZbdm6hMz9unB9AhVPp
bza+kwjkLdcT5j13MOnqBARI+IOIWf6MLhbgXujnRszwEYqSCB8Lb8TBrWIJ7Nn99TMfLRI/FhHX
tGIRCIZ6b5duBZUA9aUV8ktGJ7SesUK+Pe2cf8Tj/StPHPQ2gxRnvb28iyudPR9SgC5cWDs49U1U
NIJ5UGpb0sVi0ve8wBU5idVtCx8YwliiOsn7Mvv4aZwIPPdaajPL5b2mrZRjiFDXdvP3SCghX5Hg
Q7lht9f3bASPfejv3iD+WSvTAlFsQWvpgCp6dKs/FgnzSTtnnzh02WHam672sE+NuA4255Ns7Fv3
e0I/7CjeCewzPxEYU0XULkyuSLlCQQwFNFnC69pKwEXr4npYDWM+tgessNaesdTkm8acxVl1m9PG
3hz2rpqfPKBUqo2AwjepUyn8w17uJyWfprLFhhTL2FxejD2RyZM6zm3Y+ToQ5jJFlQVbyG1A3b0C
dNN9zWfBBUOrvmIXGHi6/3JF5jS7pevJ0C9RTZUQO0+H/6p18VOffn7257uixOgsJClx7yqere4e
yxXKiVbrTtYf6YtfYvAZNlTtMneu64yTBVtdCW9xT6Ty+JPVox+ijedXR85tQ14y0W6F6rjAa5Gx
diT5bORwg6odvCU1QNpMRonMpGMF2StIBTZujlH5PwCeVbNOH0Q29jCaqLe0wNdwULh/nNze6Pse
i4CRdic/lqr+X4trFBZ0H8ejkfNfFgD1EBTcLZDZv3V+YfEQqkGCvwSBf8wu7DPp8JENXtltQO7N
s+obIodEh80Mr0eiP7Nq5lVjjNYj1lhpgnnjJISUcS0/3oBPUVECWo/BOlpDuUBONvIPsWtwKy8f
xtVcRhmKX2e58XVuYuDuFWtG6HiCn0/BBkmKBW3spd2aAa3cMaml8OrHdtvJJ1LDcOH9dJ7Gl9Rt
8EN2jfKEPC87vCAgyEZMDpXw6BqMQcKxAfoGUTpraQ3K0SxkLNEpsylRvVZ7anBARavhXfuKxjdE
Ve/eP8BRRzB3IqVjeQCjR77LkKW0lCeQHv4Rihg2yAm9Pv9W2JtBNvUySBNvJhSM5BxkbWuykcPK
a65aQFhQuEgDBQf7V4nVX0j0lVXFhRI+DPqZynTw/OnH7NusLoYUcH1RXpkwPDmWKA7WesyEBsR0
r9X9xKEuxnmO5WOs/vVQ4KhzHdBHiO86r4OC+Vx8PJrE2EAaSeBHpH3gwVVO5kDXHb98GHVjmzG7
BPzNlxGS4GZlVDuUJqTEmKi5E7YHv4vUm/cLW+oO5ByYNG0FIJH78HyA02iQTTXX7NFHkEaowe9k
QZRIQy3kZtUhMPG0SOqy7ogRKOKB19cvJgmQda68Zvm0Z1allQohFpaeWuGGZxgw21WdKQT1iGSL
UO/jqFoYA/uLFIzqH9FpvsHVykeUi5r6uKRC8GSDxRox7F3Fmx0PvkyKnWnV3j1pmasRwfbHyYru
9JpZ/lBTXyZip4UUaqhfo22qsDTjWeA+wnjRTkwHmYHNeAyNzzrpsoN9X+siW0JNdIynhMDgX5sQ
EGx8iWlhCAzHD0tU4I3g+w6OY9qjOuW80v3b2iA3UxPjZZ/3LCZJWxmGdkb8JBlttliocYp3WV5y
1qNHpiQoKWZgohEFKcTQiMJmt/0JtA2eAaq6F+QtCCkkta4vQwIYRCOVUfPI8atfW4QSRFeMGTOL
MHzxXc9pxIiIIu5VXpfMvMDJ65q1hFSX+QJ9+F3n/UyAlJFM3pAly+Rk+iQR7EVoHiApRW9uxl4N
hEEgLdto58BJe3n1Pk+vMF7ot0GC1eAS7QyiIfTw4qV2BevutNS5FhmK4Yz08WmdGeS/VflRp3DX
oCEQbeIQczkQbTfUKhtgZ1kacaZp6RcDvwDD1KyL//83qcDE/GGZiJDQIkgxdRRQvwQFIBbj+6qi
IcRoqFDQ84ZQsDaPk3ujGAJPaEcT/Sptjqr53Hz7dma51l0xvZ5d2ofL4JngKQIH9PjgHBELO+wg
/Nz5GI8EVhMVkbYylqclTfXauWP0yLf3vKFOSxZtb/yvltOXAMyrUobCBlsUayCII8bQgG1QE0Af
5dly88DmWKYfmArBxvlvBRDPZP/XsIK/MD1VSzDECnmfAPy6V3rk5h/laqW6zpxOlkIT+LH02iGY
1wQLUrwWyqKenxzlgSbHCDKaJ9G6x4xr1FgxriW9N90GOhCaaZJwKMpCf+9BspxFm1WXhgiV1b3w
bCJLOC9HFWtQdotViF9cU1jPOBvr61uQzU1SyjM9aug9sX1G93PoG+hsOngt/9xMOM2au/0a1dAc
dE6Mi/2yAoPBf3CC3AD0GPoBTTRCjTA2SQT1Kj8X7qwORGn8Lc+u9PJ7mocrgPXS0I+6ntA9QvVs
8dtgMStMlVK+fI858r+6V3qZ+AkIo5ON6koCNplod97FUwdvxcoLk3U1VeRm7paQnjWf4hHKqynQ
EnJLN5Uaw7lrNiQutB33DljSN4kODI0LGJ02INVlv9itii8XHv+QXunNg2XVZZoij9+tjOF9VMnc
EM3MkuZX92DbCGA1fOXofVixwpHLsNjG1Pdgw8fBX9fmIJOVeGRknwtNO/9PIzPUfnuYPFU47K72
dEqe3+70qiUxL6b6BM1lnPlATA2W1XH4lJo4vZHyh/E0GF1wusXb8yIjx8wZwwNQYVvBylA86Jmm
qg49IQQeDtCCFm5Cb1EeWmXyvpZKISn4fJQuv0LZ1C2pkiy032m9CipSgLTKq6qNEPIBo82DNw+w
JSwjYRBfK876q8pKXFceI029k4NnJxAJwYUrtL5q/gdU0zG/mCF5VwSMxzRpC7Fff6xWVrduNH3u
L7zgFaGxZ4KXOrMuqUSj1yui3dqqXVCKqPlW3MpgNuHBGRNDVa9OGwaR+z8qW44GPeDouofMpxYD
adfQOl0Jt99US+qumsdE51VW2wclZPK7V2mB8UYBeP1Nt7eLOZCz0bIKQnueINSnneImZy1sDFQl
BRHIKxBc47rSuFQYYS9p6Zg+ptJjnRvsL4YSiNTb3UxU1EjA4VDiNpV80CEIoRQ58ifV3wZLZyX9
aTx0U+NxCIidFEi8MZJKoZOm1OThC+qqln//zue5vioIAISRXxHL0gQtLR4cgKH3cyvP69ioop3Z
9zRsI4pUE08lF/WxYsSVZ70fMeq53gq5Et+FhRMA2C2mh9b2mgj2gTUMgbEgCiDPfZo+FH/vOx7O
o/8VMWt4Ly6/sq8aKheGUYrGN05J/rTMQFGghLfbUO0L/5OCldNIjORkuP0O4B28EXreAljjHX0y
b1DH5n7SmWPwYqJdmpa020oqVOEvgW5OhyxVjiw4Vk1XNNIMcihYQ6VGn9oy8xoWEfyLlqwaBql/
5YW57PhMiNYiCR5mW7awLv9WoOpiB/dQUkMoYOumuub6cLzDuWm8DdAwS5kg6U2YnRLbP6eSxtLR
wTJyCvjT5Z8nxYWWiw/U13XwKrsSbIs/0W0f0fc1pFRr19D/rXoEzgRfXnyW2HxDPNHiM8xAJrUz
xmcUtVsYuT8eCGiopd02AIzBWWVSY0cX8CgB2Ad3BzTEW5466HmVs3yN+EP6Nq7zfq3724btI+RP
+OpEyttn3HqMON2HRDa25F1kXGuNcac+sXBR6TWNkU6DWt+1s/rycYDLCeCAtgBrhossDJgvWIH9
ZSM4iPvQqldRphQbtCD50xNCiVJpm4Iq4BYMzlu/vxUNqSCj2mjO+5Fi4tTiVI80MGjJ/dOjCmwj
xXIbsWIxm/Zx8mcrU57aJGb/4uP9irlTCjy1tDlF3P0/HkeHZAy62xpUzwRQxKTX2Al51t35inAm
Rvd62oSKTNjBoucJ/4pSt4h2nwCdXMktmRvMOB7Gsk4He/NcOizgFAfW+XN6Mumpbzdid3iLtLSl
kZEbsCCzvTikEERtzrWz+PWSG8sGMr2NR3SKHjjr70MXtycrZOeBhEbhfpEGtYAU0ofHWZ6FWSDL
Sffl/NCSS3i8QJOIntL5zImEULUY+sJvG9apXxajA2gqVdXJrJtaBqoDyXqgWGe3VTGVIIA9cljE
h7LaiUqWNunzCNTjCCj2EutdyNbkrDgy2sblQTYBvKVkanN1HGiOq+iSxffd9cACz0wL+eh10cZ9
T78C5JEnA4lHCHXZ2dh6/yKNVzDwbR9EJzchGhErwu7mFUxbZpF7hmkqEqazmECrYj9kSSMoT1U/
KrINLZ7g9fas00ye92hlGxT8IDqcn14Spm6KgUTQVAvRgFbwRT+pi04uHmJDhvfT5QquY1mQy4QU
fMKGFld06bhtC/OVGZcJydPo6ZMOB4ZFIUm84Nt72nODGmd2jREt+QsHKnhQperuTbHgkpFyvlSu
QQql25eVqg2+JwnYueW+VJ4dmZPvHQY+fOZdeJk6g8UJgz9HuChFWHTY/FleDFjTNaOBnPH62h1P
tzQGYa9YcOUOhVDnXV/0HI28f/FvFQ6WVIoVnsVq/tuolUayig0yiDubtIWQEMdkf7R5tp+wkKzv
2qxLUY8RkdrD5B23f03PuF3pUmOfTT4B2sxoo8OT7N7+eyjL+UKdoblaXLmtl62GAHs++lrKkr8V
brtxFcK/lM9Zt8HYS9713kazv/1tdDxW1e6Vd33Cw/1tztsV7y9jOzRzzsW0R4rGAjmh7+YmYmfz
FJEup/wlv2LYxeZGH0gIk90Dg5MeU4pW1VBvqUJj00lDBiFQ1+C74w7mRaO5zi0AXcOPTd4jcUHj
SgSi+kMJJExNLR8/jz+dxXMSQeEc31VuFaqdv07CAqoFNaQJIYNcxDg/yWr3DQiddrxOXmh8qgkB
gojHui1NPAZ7CVOOEsjiDJ5I6zq7bhAMSG8jeJnN/Cq/RJso9OxRqWvC+eIfaJg/LtvCNZCtMk4S
E2h5plUXdGihdUK70sUJXohZL2J7ihwFabukmANUoWkwlvV6uFeyxR3cR3wYKChAMJJzIURjHRLH
BZ4P+ZuO9fytoyaqZ5cRLrzpMxXoqeQmVCfCTkXswPVxfnVg/HqqpFei0zsAffRpK+cs6ZUZoOSL
Y4K+Zo7pNVWSF5FSe55cbPXS5T3CXrkb7fYrOkGLo3osgLkMigKaxuadCaUuCzkoKe/CvG5jn24H
me8H1SZkpXGbW48wi4KXFN0fRS3KuIkSIpKK4zn0vS8UmK+0i8nA38eB6qUEhAcNGLMCbK58R1Wf
O1QBNhtYv3/SBfAfEDPDtJV3wHpawvx9ACxWAFQEQILIoR7OFLNEa4YpF+uZe0AQFUPROeWaGZN6
v2Mu/f4h35IjBD4Z8853mH7ToouZKyTVRJkmRt1feBgk7dm/5DlQXyKh84D+l83B1esGvTy+PPJT
C5hQNIX5098LzBkSZXGxSB12C41AyoTKWYxth/fi7Sp7VxG26ETW6xHhL4jD2uBjykBtwpgNwHWt
bHT11ysHaBCm85d6MOvtaI/KnQPDoDjYAvS5Jl1dP0Kd0d1lP2+H83QBbe4p24jW029C4jeI8IUJ
1wo0eFirkigbsMQOBGcXC3T6PAGFykRZA7r//5H2fcE1vHXYM+eR1VI7KXLfgCinUnMp/fJlo09o
ZYX+LZYX4MAKq4RE9Uz/ChSAVU+TbCn1LWq9dhDvsk1eyZrw/Wsipk5micAyGM5Ti6Rvk/hKSvfI
IpCi9YdeokxOhZ1dxpr1JyWUFronzExPz7P2gRnkESdV9BO7tx+9yS+txKY/AvxfG9EnFNPAaD7F
TlbW8fip0D1K5O425nRrXW9T1u6NTLVJydIwK4u6/gqMOnnOdR3LvMtfjdVifI/TC8Ui8lPHtfjF
V+c8yHMGiISa9Jty/IdqzS06oOZXjBKVVRIVZ0xaPtqlezm6lp2Ifu5VA4yD5s4X2JS6Hi3UAYni
uiRgDZC8PKu0nP8VRk0/9WrGvRR5NXJ80QwA8MlH+4dbyouEmMtdtUbH0HobyF3E2Aw8L4DhKQVa
oz86UROLHroEDB6snMDblu0wafuv9Na8eq9Pu2NeopAEZYsxhQiAexFsSk1wCTMAGX9d21dFJNR6
X9KfP680GAaqhXzo3me3wL65o+NB6LdeXdYRLWFiob6ejP99+amLNRBrF53HS/CHyPCLdcTreGMM
buHyzCHbTuQXEqjGS0G2TEDBTUaVF0GHaMcJhVv07eE+pjd4kJpGkh7wUswxEan0lOFYlMP4IEAf
ZWEcY6jrJUBd7yRarOCNiP5/dHaP9WxJ0S7gHNhSlI+6sI7SvF5uiYftyE3khN93lIwHPdGdniNG
y4+oPrc5kyk4mUtTfscqOxboefpAW9v5W95/Apqsra6ZdDBXmNEJWueRrdqa07PnyEa4m6R9x6Kg
D2KXTp8P15LGB1IIGDiFbyGCfXJOOyECclBZ0S5Db8+SwTnTBhXErpIkPnp8Z/wBTH7v6El8ZMd6
igLM+sEYvAsqgpNQk9gSj47cLHxiuTrEqZCzRdLfaintiohr4WQ/S3HBQCC32iygDUexI9ZRSAK+
AonspzcmXwJsHyeSSL5b1CsGnku3C+8AiaeuS7YjPIylVnSC6/nwvPc7t9VZcQ/JiV+63jSEuv3G
ssezueeoG1rfc7vKk46Lgw8RhvPpdsUWcg1N+Z0CfZOvzyHK4QpmGatPep098GVGElblyyCbKt6W
Hxby6L9f2jDMUYIMM8DS+c98QVP8sQK7FH7rAYvHKhOS8ToP5J9qoZ6MZMpfRdIAOllQtcEiKJ+n
1dW4JvXPr8sQgFpMBopFjk0/2uwFEE42iW6K1UXajIB2ilMhbKRnnAz7fC3R13m3ZX7I128/sUq8
49JWssUjATdgFrVUSgBcCVbN+hJsJYnD2OhFAK7M9ydkpxQKV3sWCYBlrhghW0CDvufItPvTDple
3NQ2Y/1pSEphQ4ZQaeufhlFgfo1+PCH/NoRpigp0Cdq412RsTp9E3MvpGg8WgJwnZPoujPdc8+1V
OB+UQ6HAIHGFax/D7wvER4EzumXEpoxNSfVMnAI0cT9SlElD9cA8dHcCRSAxcfslOf/UQQ9hNnc7
ahTS/BTz+jkkxV0Yfxu6/M6iAc6xwl9K317gyg8Dx2cMx2U02dL8aJrvJ7C/Q5LA7lo9Grf8zot+
lJr9O7R+6eNXZHqiJVXl4Oc4xQqK1OSXzBg5q3Ura8Kzs3M8TthZhO+W0+AQVq0d0l1Eql2ShP27
tM3mFzrZaIImDlEMA5jEo/DZDVNY9OJ1solo2YtAKmdQPHP4CuXgBArpQw4360S0Sf4V/eHjzbJ/
QkatWsgUDL8wOPP7mngjGYx/hRtXfErs+yLOcIzw9Wh56/rnKii7lkp9i5nTQn+EhfefzYmvWuiQ
8MeNfB/VdYtV7oRA0RNTKVmu0CNVHo8PkwLCaLcH0yjSn3ONSCLOedB1mgNyhrIdFnAE5/oiHQAD
HYuqLRXgJMUqpeFE96nDz8/9p/1FyXQh+PVacmYuUPTEBXUnZp4ipwpe5U3WRiCIM7zV+YVxeR6W
8tlCqfjevwhmTM3DYi6CGwmvxUnQ3emNmHmLIsd2v36xg6c54/1NiA24046+It41rnrdTh2WS7B/
71LsLFniY1xhPkdbolt+PDekBffhz3nqtuZB3ftLqC3Jit82Eiw46+1QWv5QJDMbExkfuSyVB0Yq
ntvxc+IFdpp3AAiPX33IYUCWIGpGoMzo7diGK4Tala3cCTYYvBghXbHyz+3Kc8FEbCuVDUsk1vz5
TNpMbwmFZBxuyOikUl4JThnsWd0eGn0Ir5jqSwuBUBwsxyZBNJhUCRd8UcP2rHEkcOtGKJRgEXX6
QauMvPW1Pzr+rsG1WEdvM1q+uo+zef3U8zAvymTeD1PiNPK3lcU3R08PCByS6H2Q1ul7vkc8v8ZU
AvDY1oZrp6H4XrComD++K8eHkUA3vhn/xkBtCqQX1YsVdj7afZA3p27w7/C8o9h1ZMoy3GFX3XeF
RQV6tzJbm+3DgLFiL9v60r7/vRu4xvp7FhHnGeBAjFfmCjQ5DE4ytZTm/0zZtcuAF+r2umIpuowM
A1iSx9WoTI+7xrLEZkbW28/IN178bsoYFRiKhB963Qe6VEFXNyq3pmN/7l0KwEwJxveC6RfW6rLT
nQFJ7e2FTDSaZetf38P/iTzv351RT8qilSGszm5K4AR8K8xIkrseVxOGrOVvqqpuDROnPSQ5490J
pV8hvegf87K10OxmvzDe4OsNezL6bdcp46e4SMEwM7gckahrBMP8UdWmJdyW8hIDAJYM55wXtIBb
Ywq/aU7ok6arsY75YJWd5axaMOrGMjbgoLpHleERm3kCbRdaiHGx4X8loRAjIjD3mjrWjDJSRwF+
mh16+8xL+aBnUP7+V7/M5wYd2g8mZm9jlXGKNCGaTvlR7K3Ot0u09xVXY+gPva5bJdbaGY5GiY+R
d8PG8VlHrZwbx99DQa+VJp+4iLd3N3f69ACfjKD8KiHNGXPbWXPi4VwZQeNNcdNYyf/Il2IofNi5
D2Gb2v+7J7ytVd5iuqq4cv4FaUxuWD0zX38Gcq19gjcGI/V9zUgjPUKFw39m5Et5u4Dwo9E12sGb
6y1PI23A5XAcJgOI3AStGTCUSDM8z46TuiWIQfFwW5VCn88/HzlYFamQTLuszstOP4SjbGycTdf4
rK/PaR1wKCskfvh3ViSJjaMr+yEQMbs7mGlNKspC+olCT4OFrFpH86GWr0ZkKyb84706i+2ixF70
oNc/XNPu6LStjRZxhSh0+Ffx44ecAM+1JFIl2f/wclrgwAToqk09iiqGPadlsjrjdt0HDYWdaZR2
ImzYA+Z10TqQ/nR6ZRp874Zk/K/fzKd7g1fa9DKe8uqm4E6BIeyXWJ/7dJPFhz8sbCLHLKNxbqmc
edhOBIfKaukLlo+AhK5AeP//9Xk8pgxf2putXXzPaTLZrkEza5XNM2V8XLWTPgMD0vf3Bik5akmV
AzvlLOkxEDU0jV8CFIEnCbrC/LJ3WAPr284JH0Jzi5xh+V72qvUItx8f24+/DSB6IXuT11ZxRCP2
zcaVuzallYpZ2iAAGvdyNnRMCPVvrSq51I56tuYZGXsnGnmdK0o0hnfY7rB5gO9ybNTecLxuYwod
ZpkPqVYXrWYpyP5kMJLxmPAzBzXvzztW27GPPCkXf/U1uKx9IcJ+c0Fnvnx9Z0tMVGm3lRg4o1hp
cErDfaS51SP5+77dZQtWYkFy6WzgZIXeLbwWHQA6AmeLm1DFJonYI89nneqXBckTeWhBYEjfqxUy
t3VO3JyUsWb2+xgPkqIz3t8xGAJbha/I8MA9Yzbd+37dvyoEij4v+gBHNYDrAiKxvKuj8AXgcEap
L4LnmomGF1ojGRpuJNce8q1Go6LJO6NQmtreECA2IKOW+YhX0u8oMgiAHTJCWUAqyEuNBeCfTmXG
wJ/8i7I7v99BraYH0o3HKGtN2maOTauktls+5FpMGY3IZdEawrv9m39/9B544vUK2iknHsiO0z1W
DlRtwpQFT+BUWBxuuwRzxuWTfUZQXoQnQao20g3ErqTqJVBBjgKAf3h5tCzDnBeoNCuoPNhZ39AF
FStpS+vhgYfZ2rC9+eVTDeSP8mEVb09/KZrbTqv+8vvqMXdvnHrfUbFFn0+21hksDLm/DOGgqeHT
vN4BbXcJv9DpJ7odvLSCHLIvO9DV0LuX/8KVIbg1RAOgV4G0DUgeG/KJ4OR4Hpys4+xt+3kRnPaY
116vZjwZjH/Z+7ie0GW8jCCm6fQ5QrhdGSYNop1WEUTe+HJfm7c0Jl2/Tww+Daf5S02byVxQqjbO
eiUesyYZ/bHoKd4Zg/MHXYr8sB1GO5E62slkNPwGfzaJLbKdkMoZe4qrB+HGPy9TQ/akWlaisE2B
4gMBk0oB4/DEFSBJCDGJVDksp2Jm9/QzcBmoSINcs36HyMTZne3rljyXJ2SCyFI8GbRMa8vkL1+3
kqTr/YlsnDMLDuJKlgmEYiT9txIr1Xede4atEQuZ6Z8E/11D4Qokz0N0DeNCSd+drbur2KYknVPu
8c/54NBmx3m5ozzWP+nil3S7gO6GJUXo1BwjtYRDO/iVt6XaNeLJ0Hm9no0jYAosXnBh6y9Ce02B
NsBGI2HDL7kNcRDEubJXpgNtgKjQ+rnyvvGjCGAyfORGU18unJhHYnlptx8byZray4OCQSiWnAqN
I73PS3JNLzA7Y2Zdr3UxGv2Nc+niSDw3G//GMIBTSQmgAgQo+sxEUXCombALn/uiVN4eDbZCEEmd
vN+mUZgkjBUzqgPpClZBsqOuAQB5qOz7uU9YieaSVWWkQuvJGw0JQJyZGY8I6JK61gYHp/13Rdsg
6gBTzCIDDOEy9pQDqzugErwZgc1Zh4VxbTxJgQ7V3I+xl2UUGXrzU0tATTSUE/GCdF6SaZdmPgfE
KC6P/EkUPrp2/rDRvG4vdt9qNPufaD2QoaDl8V+Vi29J+eHDO6y6X7H3HGCfzWvR8JCtaW7eBDRY
mIUPJVMhIB9CF6mGdwmr7p1MEdpo9uMIB2ovd/I67lp5s3y5cD/v0jpOmeBDbx3umQKv+nd8seI7
jjVqdl9Mt31tWF3BdEDyiRMHBiG4IKmm4H6eZi1f3m7+V7q7/5ICHuPAoyIoZ9dn21mF+Ry6qvSX
2iqWaqwO4ByzJ4wtL4EfPN/98BZcCIS2kCifcGKhJnh+sc45EyXeQxKDskXmdV+JRNKJAX//EQ3D
i0rY428MG2V3MBCB1zxtlAvksR9gnMu8ECGnthUAyDAq8pV0K0r1IK+tAn4G2IF/DqToLIXpZWvA
4ZI9StsT5YDX84JRZgWue9MxtkdtKV3XG2OMsofMR6OhFb1u7N6KX/WAaiWJbCL3cCmFUeAEBjBt
MDGu5lIPt9IfZb6nubwVzDnUeQUtxOuQth/fvjswhAqSs7mgDHGD8VGf9HGXOPE/yhAwmGw07bHs
vlSCjJFFcM1iEFRgKMCfDgSCteBVmj8sEsAJgBGw/c/EBk2M3VD1tRKcuPevgDOP76Rp5oW0ZVxB
3G2X8TLxIYM6p3E0LAtGuwPWnFuy6bVtOWGyriGTWgzlLoE7S7921K8c1N9lcFmqpMOrC5a939qj
5j70AAByBykXh3k1HTS3jfkK2C19x4ziv//aHoU+elyStuNgesv+wzEDeKmv4C0lOhSZ4iTJLWQe
4tgvzsU+u3uv4rV9yuuokKK+VIAbhKjV9oEJIkdT/pHpDJsTRoeKt3RCoy00kkeqBGhOsstMkxKe
yur3CA0tjOz9782dibX6lDDHVvNN6Wz23+spov1dv/fCx0r2EZ22u9EmW4hqhqdjUhJ74/2yY5Xn
o9H/QAY+OhrpR+fZlToCB0Krx+/gtdSTv8mMvnM2/vMLofGnAp/oFxD5bHUO795Wrkseqp/pfRTb
jv3NO4pyJCbANVGtoztAIRGn40GR039Rd0vV+pwZ7Fr2zkZGJWheu3d60c8o1erskKew8DtyZjRU
ZsJhOaJO+qhlzGkyW880cWnNoQZfbcV43ESlH31jB/z/PBARRjDpedJxnQwbB/m4wa9aRbmSx9h2
AXytC4npBU6qjTUd8yGMPuzkQ4ffZJVj+m3N5X5O5IOr44o+fsa4s8it2nJhNfk23YKyMHznThfv
t1JK1wHi5Zd76oXCb4P3NBO4+uEtnuMtJllDGA2gHVtyUnDlsMsen8KwgodHN9i6QAaKaYhfsmQN
SJYfurV+3LRiPMi1A6YWcAZZRHiW+kTjyougShReduGAjfDZbopLaBl7G9F/VUNVDWcwydAF0VvZ
0nfB2ZQQ9yFpTp7i6W8YvF8J+i9nZ2cwG9y7VqRoVO1oJGnI+7ymP79PXLLf8EG15wL4pi3jcwI9
QsxvgA3tkCQeTN8PmItQMQXAQzZzcYxvXTRhbmG1jeIglbpBNmjyVLYqRS6Io5ugy0psWH7mMKqc
vn1YD9KnBnDysJq7yWuqUuQrXLZEoEBxv9E6SC/e0M24CieRRnSg1Hay2NL6j8m30yJVQBiDOjJu
2UgIz/ZsIRKjq7AVxh6qjS0k984tPjG1cbe0juCOBvF+a+LUJhkMC9jHtVdEYyt0JuBV87n173cW
yFrCcRnXuaN9Jv+37wTTspqNdH0AZjqHq7FuToOCHRzWFTELLgwGsfga2CgEIqA0ckFqCLkugOQn
d/nCOKgo/i+7//JrvK5n47wju4THBDZ8lT1EHV4iKWM/PxUPj2cNqnZ7NH23FjjqsbiryTdFlFoO
9KcQFEt4iJvEq9SkyupedUq3dM3yw2DBaXwntPQINBS3ycgerZqAxj8O/f3UEhqx1zUL5P/PUKsq
TEd0huj0Yf8BDasxMW4qeH9dlTvRZgoVl63nsCkZ3Ww8cdeiYAM2IBxgLfEaXCVGGWXvKjP/wzoe
sV4fMZBcKVU70eUizdn4Hu9K6MHBjxHnfprY0HDADjDGyOQldkVVtUSwThqkY02L9AnFzatKMkJ5
NuXjXFAmyMKaS1PZ0pnDtbsMuusW3GCmw8xCo7nbnW5El4SzDApGFcDXULOA96ebqhxSX/Zp2JMv
7rP3i+0RkXwKWBTVw/7RxV/UFcvw4SIi0EaW/i3hI1uQdmupvaXa+z/0soGLmdgg8uTUqHwR26QT
KxvixgWaSBMywnrjM4YPtJ8SefUB0hTTJvYRCgb6ixqAZ6ylxmJTLfrO0cAjxVlOSmIXfj1Zgu6N
Mm/uevHZZ/c6StzzEkF+V/WI9EaceqBPrPaAZKWAGxG5OOdygpCk6R9gkgoJg0oUf04ggb656FMV
qpiE7JeKy2UIiUyGi1+S+vwL+TzGq0+/YW5yB47kc/3aJHCd/eWdKJp0fBQneBZ1y3BqTPp3PZ4k
UE8o15YnpqR9w5gx5aX7fSckKZalZGaqpRmCpD7ql0u83UfyYcMNuk+XRQWZlNLsQnxp0p9M2id3
lKGKMKZNOpyqglnV9HtC9dcJtnmVDDAe9kbT8DJjY0dXF2PjysF8fTUav2uFitrHWvUMTuoYLe7G
jOwH7iNGnBMXW9yTnRj6QEbfZK/dtdGkl6yBdCurSTXKyw7riUoZqWs900rjh7uCXgVXfrjAbz3a
vMYSgWbq0DprgmRcbNh6MD+6idFRo0gIfc3FJAFFBMswKrtGj0ombWcV5o5BONgNuAE+sYtkryEx
FLF5h2VN/E3q1QYTtyqhC2IAp2PRQCAJPUPaK1smPDz1LKVT5QlQDDs9otH/6yCh0uqgA86h857F
6O1ux16XL+46l5QQsAUHTLsoH3f2CjseuLts+hA0nyEjmAQJVO9I4aBMQWlpp7kQ5dezo/jYCbAY
1t4yYL4GLETELlxahXK1WaXNh9E7so1TbOi5bkIs0kCA9i00EWlwgWUHjANofSvaCUkF9M0BBMzR
BBCbJVJYbgG+O8q590hhVP1UTtU28egGmt2iFFh6VUReIRGrvcX2rA03OsGaO3LAOAz0T5paJqnG
bfGG+aSKNBh4YAoEYwyaxJcvgIVsXciLrmavTKIdwu7uRqY+azor5uFq4vyjZC8jr4Sl4mGf9XDW
FuD9XQka2hDig26OJhgXh4k8w4z7/d/Q3WcT5yFzkKk98rpOemQjSSGibcZK81HzfbhyHT/f1oFN
86Y+5tcDlcJQvVduRBBNLp6Km/lMT2f9IJmJyeFnfrtDnDvMKnCNN1kfMUIF28QVcdRa+UAPYjFC
RtI1LehgqTNRtVgyNa0eEx1FW9obEAJR9L2UNk5J+PmweaL9rN2QaFmA122a87fw1VvFf4SJqHFv
sHznosJbbdxm9sagClgl+Ri/aJPuJ0cs7gIRzuGBc3GcnycpwnO/4uS3Xz4Z9Tv8Z4Pl5OVvAorH
qv/qLvPFIzJf5PCNXz2gYoqck+4PXqJCEFAFqghVUSA8/LWKB8y+0ihpp2eL0Pwpjzz1n8XvRkuu
tBwkpcnnmh1j8vAS9hT20lPU+eT1au7vH42XCjCXljOk7GaCaSyjJrre2RqWAnIr2AGINFjuOaxq
nRAKogNgQphA9X2UldvrL5blrX+iMZccd0WJTozxRcEZFS2ycS9efREjmZzk3Y2dZ9zUqaJBkJz4
8PHgaZqGzZoQqeEnZWYtVmG0ZBtiFeXMaEZlCDR41SVeHzltbCtXo5FxwcNLEtEmHNWdRm8aOkoT
aoTY/xhm/FERPPqKRZr4iuxJcKkm2gH46Lvf5JiAm4aSO2G3qY7t52sclxXgC+yjgh1Be8AQazts
1e9b8qQRo3koTl2GJTIlk8HMz/WUmZ/x1coVKn4tWKVDAfgOhoHvhV2AGMnjH+Ovafyre3fUmvvK
iBPQw50GHPYNx11knbYqqyjGHU1bjM7k90k6oEfeo9kY6D7VzcrMHHU55bq7LDypA5xFmR3zmzXq
ykM8O4IAj2PbGJZadZFv5k5ouzb5+uB5Bsj2Le9mcjTvoqvsbFVt4sUyAnrXHwYtyGYf/gbsUXn9
FKkj6IgpG0YMVZA+De93KJ9N6j2zXVkzWSjbjgPNsMZAQlGhfpXONyqM2cIQWlHYOb13ptKQyUtQ
GwAs66huv7LOHgIfqd69E+xXo8TqnCN/zzet5Aah0QlHZe4WEk+Fqh20rjcVwRercWMXqfxtBTCG
b6DfQRSJIMpcaraxfAclX9KsG+8S3oawshFFFGD6knhZgRGUpqU1slnd8HhuWb8Wv1G9CtRINMJ8
INe9T/6E+KkD+W66ZXq2oEFa2Al/tXY6q96yEtIOwpB6JbjeTfdyQZEz3pyZsaEk1Mu+WySOUQz5
9xeZFhDjvT28piMD0nOWhwLGKy0AcHGIWNMkvTI+JDKddmTBL0RnEug06voQHJizELm782QryhPu
GSWxytYyaPOn4MTYf+NptxgwplNGE+wR6wCIRF9lB0x9PD5+68s3fgZEK67wWu+AfcZd1br/3N9c
HN95BdSR/eLATHiLRsA+y2r3tYNYGq4J+O9IS+3ka/S8dMG6Y9fHkahXphpdblt7Vbr1HZX3HF4Y
mRj3eiEC+mfhmpyj7j5uRmjPaERco02h5agU6kj2ltoGIsPEPFkIm+rXJu+6M2A2zroJaAS73E6R
RrOJjSIs9iqKOdmZGKvE8ZLeFXTVnmBoPdW0nOOUVCu8wCmpVpIEdSVJP/LvfLZBiNx89OHr+JMA
IeX7lvayaDSC+ibSRZKvSjhFo6qV1iZh8lbBau/0BeVaJ0CS323lTaGGb+7aj7AJ1EdCSyStS5Rd
qCb/fHgVJsUh0ZKNdHlyYPxD3vX+OFbjL2KkN1/oZH1ckvnn9tUUX1vZgVDY+IDP5rwp2xX+D0rA
KOZcRHjrSQPBcgC7rqBtR4TK+ccuwnn0Z0HiHFv0sIklV9FNGEvrGyNlKgd5ljKgVC+sJzQm6QhA
grzIcr1foDc8Fxp28r1I2jK0hBtlNElLmOWgEv0Smq95MujDMd5JFtinckdj1Fs/FlgFvSJ2Gc6C
0+GOLejIb1kU4dxkzo/61Mrqq8Rs07JRR0Eyl1IzSCWLIzKyFOPHJNLn1eySXQS3SzLuRFPkqDbt
/p8eSiN1TmJfDUm0EMTfQZi+32UsNv2REUPqQ7NsmSTpl2XOb4GqMQp2s1zHomXkzxQUtk/OSa0a
O+X2j5M6/PzcP8QXhl6jAZLhnKODOMn1qSw5CMQg9tAbhN6jGB6SxRUviq7JPtxwOxt8jLgszH+8
LFlsyITR7d/6JGIZuIRu1kGAkAGeKdyCn3v04wxWxkMHWEfEMZa2woeT1aqWuUcN0i6r4yEvg0Kk
DKsevnPw9dG/7HZHujpZw5Q6tkeS9LkEd168LIECe6JWl/GVbdvGuoBbONqOwb5vY2gdVoFsnwVY
Nrcjphf2rOtmYyQYLUZT0Ijr3VCI8o4JD82TC9n/KlLwGI+6mPwCV8IIkNZLi7XPaZv9T93LLPhK
KqJ4UUQnCPCZhSp1PcENIfe8qzEO2n9gqB5Uz/Pxej444gxoeakSgcOSutvNOwNWwVSLwszuipCJ
vU5pOotPgl0wHvHDE9aAFDc0xURvE7Ve83udwDbY1m5mQ18Hf4Iquk/sC6v9cTVpMFRN7LcEIka4
/tXH4k7zGyIyTRDZGDZ3kUHk827nqSlK6GbzLHwwbjIlqF2cRjuaKVE/6zIGszdF0FSe8KBabz4E
R2xe4MwcPfH6yUm054TuEmFgMTOvBDPSp971Yusp5aIrSxCyDCR1G5oJ6cSMHAiJDkERjqyqI6Zv
vOssfUjouc3gs5hwOeVL2i9AW+jIj3R2l4k92N7JKU0OIPJSbts5Ot+xziPL44T0+/3k6UA+67OZ
eDNl/gMZad0nPZRbTy9p9r5ouewG9EXGtt5GSd+Pmd8qTaS9gy9oG6aE4P2bwxr265n+83mPqS8A
2aKOuLDGX+/y9DSN46jN2pckgQLOGd2eenowLs7vAPgkOzkApTP+L2DU6arnocEgOpSaj0uTi5yh
VhsusCFpJP0l4Blw5ab3teCusWYEkXUrjfg42L5dM9CBxdGtUCXyvZjshHWZ5Y0i8s8uycLiCeKV
VLsp/eQ8opHH+svfyEMRjJOCtGUvp05/4R/E2KchOokHpAG9CjWCMR8CuxedS/ch6J1V4kIAHsVs
x8AfWjW7ZNvFVwuzXWLjc7bkwn1vzxhCCaCA6ExKzWn1ZS2sqtcSPyZj+P/taGXczCQfxzv9uKy8
MsbKGuaPNldH3s607ev4rKb0hhlgp0zmR5bC0YcrCZ50o0w/63r8N2PMI7/OyWvNP8pZPW/64GJQ
KOvrhV1mmF1MVtnr00IzQ4j9EGyHwZXFE+I0uMl8t4Jsp55246g40F+/sxjuiedIM6vds6OsBhfN
MVZ/8bHRIX//JkE1yQMUr0D/uUxBy3rbCuME3l7RsVfgw6dFauIM/OH8YqFfe/V83YjvyYDeu6gb
IN6pP+pUQXRev14DF7x1Ca8dAzTohGf6YwbScfkfF/Na/dCrTKiC+W4wUYiwejyosGR+5klTmKzp
Y4O4YudB9IQPNQ071ENmroZjvGld7/UP1XWJNUJv/CSWyN8ridTpaWShvbE4fqzUse4kHizs9EW1
KmcDDMbWPYOTpDM/uig2S8JAaShztksM+jcscN4bQhfn+oT01gjWrd9gW6+4ysTxc5UX1A9MC/SQ
uFtIdiKnKR+mtjYxWZyIjwOxNVUWDXSZrpjB9CxNdES9Ut9tiGffBbYgI/b/k03pZ38GuTR3+7f5
WEkjbHAJCSMzcI+nwWi6T5MmL0EdM3AL5GLcJQsaZKwabaSzUKTc9Uuf1vI665P2JSQcXD4GeoCd
XVUmudHHPKEneyPDaJSDakJpHMp2gLpb+zZnKZnr3rOsagETIyhjDSSlkJItk/YTZsqbLI8gI5fC
IYJNjQgWBVuR60muRXljmTkZvbrBttNr3WOEwCjlEMXTt+HL/bSxWup1dYNm1uvyWslyl/AhsfLU
zkLfOF8pAv2jThKMeaCR7r7dVs/KTZpe7YlyTLegATGhL8kCfLztwR6l+FDRrqPBx3BLqhRTxfVC
WiO3p1StXNYD+S6Heh2/gft7vIRToKUwzFB7x+EK7Du7H4hVjlqOum3ytNK6GI3bwLspqnx0fMih
P5BaMuNFHnOgom6ojpWEFLGeeo3Kftm0v6lvLdeB3VshW3bDPItUtoa0s6m2teIQ1Sh3wN2uA7oi
D7Y7S1s5nFjf3JnqvZPRhRlyENK5DQ1kEdx3d3AXMgxmguCWghrghcD9lrzqxGQW2fClXHC3hter
ozM7IkKa4l7FKSkIuCPo28J3EWYUZIzxE8M9ESWejjZoVLSDpvvUxdorNpMQI5pdUq/NphXoPJgl
941lnNcF5TQ0h9x6tmuFu66MqQpCyHCNjZIOnzzeOkOza4ZVL7EC/V4h0Zh7VbmwVu/W9x2MBGvD
PH82gRwNwZpXAPmvhjaAgyu2LmnkJpk/5crjAI8PlvcxU1k76a4o9SA1yTKtiggRTrd8OUZz/Heb
RKBjT9tbxsqoS/UUtV2xhPu3aPe17/KLGMSHnfvcHJcQgJ0wxvAebI2bH5nkTb+NtPRIVmlKYVXB
ESni0wpeqmI/WAQLGF7bIq4G0J0jQYTWxyWPX9hScLyflaCnZDmDkB5PyKuuhaFpk6u1IaGv2aIi
tm206yyW9HyKal7sJUNw4rMMxF0yuoICt0kDEJdcjHC+ueoAlx16W00Eb+tabhaerx+bhMIvKRA5
F874ESFBQJtwN3sOQNrmIAtE/9YfWuuMbFhYzryrGwNEyhXP6W1sucVYWcT61rfPUvqyqhsAbj1d
n7KFV5peO7IPIQLp/fR0Vw6xPgmnKI+GRhc3vFbZDL/jiP71FquLZO45unTXz5/GtxtlHTCUz6hb
+PZHSNuI0VFYN5GwvoJWaq//amh8R1w+3+HzExmpMdF69pKFgaMKabFZKq/HTyDLzrvNhg/Lb5yL
k1lGbrvzuE7r1Hq8aMEQCzYuQ7ERo5rfYJd8lE9UIZOxVJ8KbT0d6L2T/x84AM03JE1L+LntaBWk
V7XX44VM7/962r2DPcLR1/LoCq6B7LcsSJi4LIJ6iRHT8j8O7W4gfwjglQoBHoSeiFi60Umg+7dt
tyG1HcXosTcMLhNEWEvgIfqAHxCoeG3qO/NzPHNgQJBgJb8M8o8wN34QbfQSphdec4LSS0tG6S5l
i5TAOVb+ytsHRmPhaSpLk6N64dsK3j3MPFAHPGacF71AMltjNmwqTOB+GDKnQC6xKX295jVpo8iH
gtOD0aqLiiXgmRnr8UFpu61yH6JNwrVW70o+IPeGCbacg/T9ztuz+/bJKnu8gxYi1bD+ox7EWw97
eL/pWsDbnEolzwIT1IeWZufcATuDiz7lb71JrfSiHKhj/zQ9F/qPvIG/JCUoI6ZFYvlVhB5Wfql8
kykr2JpZjzsY2d8c4Netul6g4kreZAFZib4uptvWEhjcbhxwWCWmFziOlTtIQT9fsLuoHyYARyoF
Gu6gJLw+VqvPziUDSQbrUSEhDQkrxJ8XoYJnuBMsD3hkXHdFD82igEXKCGCvXYYMSvKKoymYA0Ze
n6FggmpuWJY+el+qJPh7hSE5V3D89rpRE0ZRfzTejD2YRHgQAQ0pWioWaB5eaT7k7C63nDRxfQ87
wf/nLsZKioqJM5AwTU7BVgVCxg9LfWJeYX9O/YirkOi52Oozf9PmaL/uAV9W2ibzwrHFGuz05dk4
DLLm6Wl6yJL8EsnGEFltNAe7yCcqq3UKDjDCD369UMRBzneQ0I7kwh/VAzNjjyZAu9MiVi88Vc9j
s5tiLpcy5vkuCBFlTKdhVG+9XmDJz1x5A8Fa5htTquuSKL1XAmIOEsilGXs1jTGDhXHc0ZISQuT4
Dqvez1uAuSmkYAa519Q0q4HCLhFCKxQNocwk2hlvfSLZNyc8qzhQLjzs70SgyxARZweogl5ZIqLj
PyzL2jBywvgKnioNpKR1xxw54phSGRoBmaPs/Zn+W2bVXLykwWDl/3gt8agcDulU4wvUXlSO4ViT
Ckp9fHcuOSgpK8h5Uhq0aI3OSXp8sQVxLd77/b7Oq7AbdS/mmLVD25UbWdC8nBNbzQTJAigPLjUd
vlwSM4IF8kKH5lVGjjJF03RJ/vGbmAb13j4sZFPSbHKfU/tF/SwqdRy4FrslR6CGW0iK7kz5LWw9
NpUWuvRtC8+lZbLIMIZ11SpPLRyy+UUsof7k7U1GbRp5j6GCAeOFM5XG8yvk0f1jFrMSsBp6VZbl
XBRcz5icS9BdyRptDvlZN3nXRrQLjgMa6ZUNWYN+hupQLFvNPkkOh/1z+epbSlfzNHhh9dokK+OI
MrwwWOKPumtIFLE6oSH2bUc7vLopQyDsZyAHSD3HsVc8MaFoS2xXWU5rnDMlovkyr0IrlnLQojfk
2PAsc1teXyBSbhND+onOsCPT9oSusXwylqv/zlxpiM28Pq3rJWzUvrf04VCEnF+Kl3g5utGX4SrQ
g/cwUuEzKnp/XDTZB/6AmRo54YPt+WpoLSXtuQ8feowLGgndoRxumjSpenMonM9tSvRSDEWYamCQ
MOEMYpX6Ke/2tQrTRyVBezY1HXh3lzv3l3i3P8Vgk0EGyF6TSDn/7QX6rX8YR6ELTniOQJkZtdj/
KTLdu9Ny+lRoYo0zwjNsLZidi01NpPCVzvIflPwbK01E0vU1KqNe58GFuaTlvIuFNMIoRrXm7L40
88m8qEDirJlF0dDZL/6x++ABw67cI/c0xpn5UOXrVg7aUR2BJe+eN4tmXU6VOhVYXE3Q5wEjsIrK
Xq5hcV/3ygooktlSWs6Ysjl5LSui6eKAaGbSnFK2K77NL9bCOeHfTScbxB+tzfKhRAtwX9FEgQ9g
hAeqEAkNkk1S6y8zxiYPA9KZ0FoU6jzw8UMXqvggZWgMHTwgxLUGmUZ+BkLbQFLmmuVivuMLRvpv
TTs3aNedKjCgu4fiwDquvpg61aNDjEl7JmImYUwH9NgbeSRec3XXzFVpLvfdw6eJ0cxR2/Wg3rbM
oqLfY4QAID7Hcow5kvKMABjUhCUbgtTSmcospwizU+kvTJ0Tgf1WLODlkt/iSvJm/kAMhUH8v6Jj
21+MMeIvCSUoim9+cFJyDw1AStjRyo+1+JZ/cnMsJrwS5uPlNHTE+aIhGwDLeKv9O2d+NGF4D32E
7ROvm8y/xkeDf2n3FwmYpBfYcGJMJ6zx6MALV3K9YkJ/FarVT57SQRZViHUaQlV8Pp0II+28fisW
D28PrWn/3qUlMODlgvXE+9R+QIJ9AkcnGrCamSU4epmOKakQtT1+2JnnlPi1XbPq7qEAz+JN/uuh
zIpzjJnhE4mtNstbz0gFMwcK4H95RLg9Nd2spB+fLN2O6C8u6aikMu52XdtWoEcN4jJoxIrjEnTO
6R/9c+6oqip82miHND8rILS9xL8vwWT1wPucX38ubWkk/r/wbUg0QxTvMClxB4tKRIxKE/SZwQx7
fUxVHGG/Nan+mqh0e81NVPlcR2iFSGCnI3da6R9/r/epdydm216xXgr1ENGCT1iTuQoOsh8JWSRo
MmhFHVOZwGKhxur3aIlvdn+n/zV62WVfnv5BBNGBuNTrmYrzSCgWGhcxOx0pZR1O73/72mYJxR3o
3pbU7BArAwfgcUDVC/bs3a6M6H4Dsft3estaLbfRbIVAUQAzxz4icmImakmow89JyiuUsUaSd2kE
wG/XuznGfJdFiv2Fk1LV7IDkEMU58Cu0Prpr7Uqm50bg+x883pmSYsYUEKzCrB/aJnuM+HenIOg+
RgV4Cny6R9XYi8fdzumz6sPtL2p130pnnqEUmoaxP0BbWwgkBbSfg6QqaYWwcs5RPfWAYGOtiUh8
yOFcI8NdSu8nLDjvrucQLI2o1ZG2CccEsAMD3roZ9dkoBy4zS7NvOfdBSCkwUL60898jgYn3/SNJ
MP46jBhuvDOQeL1uTih4JQUA1blp8q2GbyaL2aXPlgfSdan/WKz3yEb2TvSKBs9PqAuhhKkPso3Z
16CfJgpTiXjZIsVxBuHVkqp+CMLdyVYNVypJ3EhWK9xOrdlBGmt9RhnKxTqunUqC4mljIdnffmPL
9RY71nxmbWH/zBlhhOA7/cgJjkuzLL4h5an8WTy0mVNiOS9OY8g0g9aqzwCuV+2Tp29Sxaldukzs
AgSj/+g6z5t71L1UxHiq34rU5EDFc8X4PbcWwIuz/WZRy34PQ3HEcoV1wDFslG/4INxmihO8WHHf
fJIWMxFx/xvtbD52gAnMWIU5Id/gNPBAKyAFeciCRgdbv89Oh3ugCm+gfUj+ncY5nadxoFAfE1NY
3pier2aRJoyWFHiodduDP4p4de8uIM/B9qWEb9vvH6JQcul3tWujJ6wMmr6P9aAWlxOj4Ehe8tS2
eoJ0OP18dXYo+ruuYrXn5XUQsbrCfb4IicpojcvsgFaWnAPdXLH123uTxRetJb90Nxgwpx2LMY72
cYyrBL8NCQJVkbnEBNaNyY10mj9jjJBpjzvGTeIObiHAPqIVLZrJYTEqVEYCo4qIiPWsZPo4hsUU
4qejIC7G9/RA2h4UPR3Hkda0lfqh2bYv6fv3Bhznb9YPMAslHzUOP11a3Mty/67m7FzSwJT7BJhX
rttQCVKT9YeeBA7TUSlFBAlnBRQaWM1ZIAEFcq+3SWNITPFtCp/XlhDzmS620r8Mwx5K4qX78XAw
35rQGMkyJsvKurTdlIMOJCNcXDZ7AFsORbC/FKY/FMUGXruC37Dj9jAsthnN091FukqsL4ql0xNR
Uzm89nEEBEcpbl1nfIMhdAQsKd0SkZxiWzLyw4t1PjDMQBQqy5frY1rmMG3AFbk96H9xhSuhGqKP
usFcV5a+cYuRD7vcgsoAuI6ygFefhKnyHOrwGb1rJDlMQa9ktD+Tr8qRiDvu5cphD0iL8P3Vf5qi
nUkP6jaVFUgM24NBajqUNQSQFNFfMBNeG51Eat5uKZj4N+HIUHenPnY+ZFSYlumPLukh6fv0EQoX
K39ajSaNmd8dOMBozBUvk5fqan5g7qL5IV9bPN5dMLJ/76mZL+X9n4wELDThoPNzVPJ7DTce5tRt
Wvce3s3XUhMI8GRo3LqveCEpEHAmo9JcaBCizhlbMRqhCzmwgfBDmtiBHE4CkQZNjfrsPudXahMJ
G2eA22+GLGaRRGukz1MpGA5dZRIsqK0Ub4WgEbTifgUK+fXxSfbzgN10NPiD/qYDmBGxa0LS6lrz
tl40hEnoyy+10/Mw8dFK3DtOL21PVuuos19AY4MDp1TWc4om1oOEirI2s7kqH1v6/9gVr6zU05uC
yR40yAmDgp+pjahAwkXXrXv80XavrmeStjhzrldcrG7IhMRmV0vjy6jJnplH+La4879UEsJBdGB6
DfEg+e2GdWGn8dqARsvl7+bjW/mNHbNPClkziEKLqSHy0I4c4dHq0NZRSM3SnOmqYgWyX0xbcUB1
A01ZCwldJY9aKD4glFh8t+PU/cH5r8A0bP2gCPCEOzsws8hErCwbz+Eo9NqrrEPq211puaz9+tEk
00xziMznoJqCaFMDuADes0GOR9pqOKDz+hdrpHYx4rXzjOXk3F767Ag1XDf8zLitw3Yzv/TPM2op
psL7WRFGPnBKUbc3jKKuRSiXgFKoSSOKcV7aHmOaOYyh8xLBjBlQDrHRrIujvVR0Zs5c6clB1WEL
HTWYFfozFdem3SGQhDER8S9u/cx7kNYxGAEPgUYOy9p4tkm6FXC/QRThirO2v4EW43YNZLlBillX
ID0nYER2vvJOdh1c/6MH01p0qyV1DyNBhv4vC8hycEIoBd1yHjhaGcmhUWJzyO6rnKENcHg2WWFg
zH5rXJq/QDXKDsUMt//Whu9zu1pIudUeZoNqMsA4ct7EwzCze7vLpgh/+DmEyQH0rY8A/nm7IERl
tbu5DadAb6Wc+M5WVrBI2z2cTxKuwDJdG63vetKKFcY/Ppqn7g1jSNA1hCVuq2Q1PwrNNtYZ71CY
m4s7E5lS5DfXYkJaYdsdS6+2YI/P90Q+6zfMTxGVLdVJwoium3+5LXdBHTnqFxuNw9XnLIn/tOrE
t1GBEGYciodDde3Qw3nu6OCVz0uj5RChWRpXT1PO/NyRPP0fqTwpUGaggFvZm4QZ2p0DUOOlyvs3
L05rkyfISElRsbbucZdP0XKQAzj7M51RgBdL7jOcnjysJBOdRhGT98myd0ivQYYEaUxBk9wXKN+M
/ShJ4wp0GFQrZDz2+2ln98cG9O0uC6v0VcQSLf0X60Peknz1hTe6ncXFAqcK5N6e7ac0OTNbpKAB
aM6w02cc/OYcC9kmR0fr6XV2e620anEeNkfB637mGm2KcjUcWI200HxColE62gsgqPqWCz4Dnbgp
zhTJNmcHaekpAt/affiI6oF6mbi3v7cSTKSaUvAM800ytkb/ejN6Q3u6MAtA5Gd47eHEjRM+U6f0
tJxJXtEiWrACnftY2r09QZ6snL17jNdFhvPwggZXJvS01hV0amSbLvywTWflWBASM9FntyOuvYef
6W2QQbdLHNvOJfoznVzQ1xpOhFxbH+u2mmcIFkBckrP3kUxvdGgAwmLtu7a4QyMEt06sAaqZHeHi
2ByqC2/NnMpzreF16Amk4yeNb+mdKE40FGphrzxOysB2ylOZ5AiOjVv4ntEqZ8xGhZCr0UhUzuby
mFQ3at1b1IPjhim+nT6wxjn5ZjeyDwPqT4mspc53fGf12ztckdmq/SqXPFPIVg8Iu6fpt7uw4yCt
AkHNIr/3Q9n3FlOBI2DYvkhcu8wU6+Dj6Fgyfv2+JC+ZA+LYPke8+Jh+MY9+iaDQDqrMyLONX7BI
FR1nWhpr+6hJj1q4l6iAVvviOWuEUrzP0kYgJeOCXqQocojXyEz/mKiRGgvkKvLeRZRT1NQX1IMe
x+u7r90GCnfBFV63+LyIw/L50AyS56vawzWnI/quPwV3Rztx6R/5Bsc2v06hnIJ8z9IXxNSy2a81
QjmMxSbsOpMJMASIKL9ZD1tDzPb/VhvpifnOEDfywjY1GqwTFxTeOT9k7hUOtAlxaKQCIOkGb0rf
L4J6JecREHrmvO+TA5c3MqTqEkgOLv2dOPw50Uj0IZ1vYFhWzdk5v4ZXDlgXMrjPHkN7d3cmOl+n
QVtgYq6AJv0VpjVCczA3tkXTD5eCMak5ZfQT9IW8KusvB+yr32EJhXuuqUPpJpBCXmbeQEMXa9Xr
dOItlPxw8PFjk3O48N/ccu9+DXKTch4peHnFfwlcu7W+Uo3a0dhHQauf1/UthBuWv+2HXopXFdrN
kpp8Xri1vN/hUxIV4kA+np8nH3cU958h3Rvlztp4fFaQmpnXmL9qi+LJ4Y/Z4F/wx5bbWNByb4+9
qGCkGs6KW6/4CCw/hEiBjPgI3muzkUzhDJsH9BEdbwaJWstVDAnDoFDJbrqwDII3vAZQP19WaVs5
qci8zaj/kZL6ZmspcD7TzHJd5PheFny5rFC/Qx7D+c8sHfEcYI8kFD2QN0I5LQneInbJasV0vKJ1
eKTivUJJEYcW+yeny6HXTz+ObWLtHtlDBUqAUoAnfZ/Gj9gEpQKfUdBrHIJigxdwJEN+Qwlh6Isj
dnoYXM5QPLbzzt15/LOUVFBQ1VrTA7VP7+eAD4rQ4oXWj6zCfWNQfHEoTg/06KcQqqlm5mviD12x
3e2MJStfEeORdj6QqQMPPgaXwK/RW0LAuJPwpPinL8VnvzAHpy4XnX1E73xTMt3dbsyzzIiNuTsE
Esixa14WqxWIRlTgZv1CIIAGKWmn/sSPDkUBu874SazvRuBc4/CXqddR0WFsYvRv8DIdWhnlnv55
rI43EM10BCJPaMj1sd3gloVCqNEtwkeBAqtx/AXn+mcvvzKpE94Gl7YDlJ2YKlcPkc6W3pEn7hVa
iPCwL09uNJjRHoTuym8YMZYAemEa6a6tqQ42m9XzSjk8cSVbzkOvLn6jw395pYEY3LUPanPNyvRn
EYtuRTBHQ21IvOqd9GGWGhk+wM3lwpABJPZrN3G72s353jYErhLeXjKjSMB9MAiaaF1Kw/2DXTZk
ggGew7djvTFDULC/ZyYOX6oVLdehPWlKV/EO3ovntVFx1e9OTy8tVw/rg/IjC93zGWUVUDUgw6L9
xt+u1rFeZTNIdxBHIrnoj64BdKCZWsmNf8F7HO/Zhixr5BJEHKN2jNnXlqC3+gDLHOZtDS9Bpy6q
HHCC5ZpLL19MvY4r/LakmmyB4n2O1dtMWFLW6btqg/sVujiNkfKRgBscKgBJas8zfkfZjEfLLAed
PTAdmVf8AcW3RUdiUNaGymyi0LpDxUEKA453r16vWOkm64rC5gZ9JxdW/NzegFfaopbIi3xDpQUl
tI4mHNtWn6SXbDjB4Im50v0jKkA/EgaJFboeMLCwhtCIrhwfpLw94dS3NObyIeTh7rX5aGQsNZA3
ps0qKEoQuI7y1ZyZ28gKfGfdksRnh3Tm6pfgikwOKLgEfGnTEzFWEGaZ24cj6mA7+vcBRCAwv+Rv
UNL15cbyMHBAi21J/IiNew4166v2DuOMmw2B/FH7KNAczH7729AxCtpsgRn7CN4svm10NRbuCruP
YPP38Hp8YXys9y0+Ro+AVZ5yKinGzMuG/8y2KCuGdgSio/1G2rkNCr7hHhNOQEEe8lyivfRUZIMH
kcvkl8KEEkTfiSWTpR12Nngm/T+PEekcXPSXA6OEgNvGKdzHEOU/jIeAUDmh1PqnDsGN8qq4/AEi
GENWjNbIcqM7AkaffjDqomhROkIDnN05T6DGSKE+z7FNY7PJ8ouAU3GchffXHTvmqVlRq7En6nzl
FF9ZBw422KSL2CWdxET2ms3s2R9SS8claoa7hCx1ICdcs1zaSTmj/0jqfV1m06LfNUQwabwjcbMl
6r/sn6PTIz1rCTErotaAG60VTJMuC5xDS8wNftsDxPnv95AIZ3ESYo4dGbCfL4BnAkjUkzXf2zsR
JeZcCVZerOaIBUcinM7G1aIkNBeEDDr6AWq9qmP82ZkoydLhKtpCRa6yRHc4RUeg/TbGjznaxYI/
pOB6N65T8vlPp3/Soni+mJ7NihcfcxvH+2C9JT92BxxE2Te8ztKM4zHasPGIc4d29znTHnVXCWGB
0VZ1iJ+Wc8FI01E2JxUKyrM3EXI7JZzl+4KPLR5ENw+EU3pSow3uZVtMIoXeYC8Y/4G79ovt4SsB
mgXSRdQ0E99Meo0KkCyPz1ck87Vn9+0pVDQhI6JF5tY6cMRAbcOluBy7QxwdekVPyb0CHLtBKQqy
61X05yQh6Bi9eEQdPFAWoe8UgQxfRB9RxqIMGid2k4louz+RuqArTTRAWAtsoNnmgkvc+iJUK0DW
TbwZeTjNPrik01OhNVixIsKDDkyGyYDUrZousEyNQgVRoTOAcm94M1vj1WagRheI9ntGqTR4Rlj/
F2DCunQIIDQ1Bas55KPjdeF6bzqWSOb+GLX/51rI5Rf8+lS/L2V0VbA8Bh5EuC6jjbJb3waHszid
MxMU8y6U9uHP74D4uLWU1niHnxag9IfVb3hobBveeATMX17+3QphXRaIlwU8v+3V0K3/76pvk8xN
WplMpuQBg1/DScL5zR17g6EqPypIk0ztEcpitIUddDZpATk1/AY4TMdsEDyJNqO7r1oHaE49icMK
1++4E3PtD3cH2g/DvKmoaqSBzjwwo6rquL5ue7oX18O/wCQTWVw5gplpB4Ne0Xr+kWq7uhmfmR6e
qaLMpOX8jOUXW1N11VfFMVnexVl6pElEKk+RJ3IhrbXtDeLC2gr4PhuYoSB+2LFUladOrtr3uPGK
BetMCTXlgNpwSGLdgMRaca2EOy0qRBsW+gRFQ1u276JF3RDNrqes1okpCJmv7jOx8TJW4USIjqzu
VIuGo1gmP5yprKsL9PzjUYYbNeFtCBB8mA4DZjHY2/3TtXMZtRuRwSaKPMNcj58g2tL723l3cN43
aIt7PaNLIybiAJjO3Nf00Iid3kdA1yeDnpknSfFn+N4cf26NzXZ298ldYj2VrTrZIpAnXxwu+Zby
NJS+FEEYNhrD7H4BkU+ZR0AkUCgupDUUsDCmB27hPvnXmDHTN5rUidiEA8+U8+8fFnSgd6+41/Am
iZjOcFL/0kNBWcJreGCSaW+8Xcg83IbEYIFwN2OABJ5tavraGom8M3BG8kl2jNkm1Kfp/WHmfsdZ
d46NANjI6bYkQSw/4E/VRgvjjn/Az3FZPBJKKXF3N2e5qvK4jTL+Wi/GF26IQbtsq6t1ZdQqd7i7
i/SHbRtunvrqlKgxtvWwnhEFQtm1W327EjuNJFoNp1yQ6Ee3L9SKYQwzVrXvyTde77MOwisMrLiU
7ZJt1/HgKcHAPYgvbewIslqvHhES/RfzJbG298ld+UfcUAoKE14Y49bQ0KDNoC3t5764EztAwhOz
NbOGMOQTmrWmYVmLcyzSEIYLmI2zJSE7eOjzNh8o7eqZT2kFNZfurtRCqwwInro3Pz8bfuwW0Mdx
aG1koWl9JvLs4oUJhCLJea89H7vNSfSRTJqPTwmfSuhpwfWy9OYFo2n6Dqr7gFLfXRuQxd6WnNZG
kbX9YhVGGH0GQn0ug3or8AOS0f5EJjSsnDG0EmxcsUAGGO0nok4KE53zTGobDfe7c8SFF2n1TElF
jDqc06WbzpLEbHQcjRdOKJTY6dHU9BR4kNs64M+G66sJ+4rtq2xwXtHh5RvAYcxkOjlVglH1FoKj
uT4uUYMUYLmTZb8Bo68M9VMVH33WXghOoisd49dMngT6/KRcP3WLpoR1G43GMtlPQK2ZOAWWVGCX
TGC0c9FwWgw77VlyMUxqHQGsiPnvq6hs6u/kTIuI7CA+C1vbaNFdKHgggtvtGGx9vGbefEfwVfpA
K4qQQcftxGgU/CVBFN+kENUk2cpDxvU3A8mRGrymmnBLeXHVMqgCFTBR2dsYsj2POJmUNhkzyVuN
kPwpoVrah1Rzl6rPSB+s1MevZEwonygbWoUe9QHU9xlpr+ySCZdOydAsfu8YtpEKyDOztSvC+Exh
aSTCpbpcZhLJjAZDnYJkpHNj2X0GOJ9zcOozwWl2BU9D5NpRxFIkmlyxJGFZ1wu0Fec8oyd2UzkW
ZOhnCula99y/E6v6VHTphdd6pb9Y1/KP94Ts5vvjC5uH6gQjLVHiDpcHz/56krgDK7pdBpRjzcD5
We/BDfmwUqmwzwNH4iJ+1cxwom0TBfk6JZkcqYr0LZMd1SB/6SzUe9g/DmDFokFgODWj4Cy9AKRL
V7NR7VLczaYUmazMit5SWyTITsa5jQxDDWxLYIzJSy1QXoKokR+H+pjeMKMjXYP+KhloqWXOAnQ4
c80uwbrTUtDJfYsNjDhPFJpwFJMYrGCrgBmoJaPpFXZb4V0iDnpTrQY7Nqis+IL+HE+UcZ2Tc4lH
BWRure0/rsBsn6jJsODhIE/bSOHNV5k3VVSgL2HgylYWnoBx7jEkO36HKLYlJYvQK+Kiv8U/J9Vf
JFzxSXiWyuvcrrG053DP4W1HywdPdbhZrLn3IlFpN3r52KMp8e3RKX6nL8EEPHeWBXr149MpPTNM
BBjN190bhu4+DjyZMda3Cxu5F6W5jFvbUgwha8H6+7xbas8XeNf/4WWYCvj6NcexgUHruZIJ8jMb
zI2mrZWwlsQDy6Pt0J7RDiR1CJnReNmosPqoIHJcglMCZsSvURWp4m/iadrZtxpcDqeWQKq6KYJm
MZuqRdcxPhTrUKsnH3YqHwwNmDCCKjF4kNsL5X8sjCGMtHpUt2nH7RxAbrfxzxE6HhfMGCdPxzKK
92E6e3uBXPVuypCghxv/9bc1u6EDr7hxlqvbVd2XZXSY9qwkCneRlVlwPGg78Kdq33bg/pUXL4bK
FmsXWTMEgYcj3Uj+LutJjtlx/bD1VepxBPiKL4zy1emOdrMq1+ly7OHXnL+SW9HvHm6v8Sij0iqX
uZIU0rtwVCJ5KlI2Jr+AgMeH1BAgdSOUZq2x+dYJv0J0ck+nWtNF788ZehoSFE5kxLXS9sTjzYPH
SoBwXil8sDVs69+KNszELcp+Shw1teYeVpP938bP18xntVabLYq2nrLj8P6QnqYL9UmMgESY3EJg
+8jigjSDlEfidiBSwXKciLDHyQUGstm40XDbQVKxd/dJC9XNZndM39v/LwAwVrpOlM5JjnZLWFif
+6OvONMBx2Crt3FG7G04vZjQN+GNFt/+oso9XC9b2qMexl2kpE+39biZ2UdD+LL6Yalf1DWoxU0X
+FVles73wxsdMiTyQOjXoTcDFWWKU2tYLuYm9ySa5mm+uA4QYlhDqjBtLskd8VtMArM1nQ1eBK0b
7xK090UMsVcAyt0woBZNhW5y71AQ7BQWpflRPFp6gfGMRVZqVXPkfdZ/IaqWS3gypFN7q5prSx+9
Kcdl6hSybtd9SyRxt9d9BHo3o7eNu1GFEthqgVc5Qp7N+hfuNSiVqz5LUZ8vytkrhtnKooVrpqns
kEc+Rg8Jd4Wm2hBZQNqBlewiX5eOHSxr9zwr8ZySu4VZgQmOpaOoIbjA/PX2Ko0CRf0IC79BdrfE
wW1ia3BLvJuLoif7d3LnKH1LyqwYDvpkl/A2vpf+h9N6YO+3fj/zzKaiNVtsUoh2EbtkRmY0GHiU
9CEaZdnNL7Ao5fAZBKGWnafS/0DE8WXWZZDLB1Yv+ULhmKmpVi6xIW60GGza7OPsBXpjJcQOS3Eh
uORpmTdvuyLSu5d2w6J/BXRWGimiViF3Fi17mMP8tni2xhQ5a3del5Rm6A7EP9TPB/o4nTK2UJYN
aq5C45cxZkdgDEQfn0mh0yOWZm3k0i63iSz0DZW7AZjfkW46D2UNBHSJzObjY9ecWRLuN29IFQch
iYfzQgGmvAL+M8lPMuTXwYmnbtY8Ye+h+yh8ROdQSc6OokMpAyEUcudgvHjQfAIxHh4DQS5SerlT
Ay8E2d0PyVSoxfJafpSSwXAY9jnxfzcrUMe+U8h3yPXwRdp3lENkrglzqKhQ5WrS2BD9nPva4GiS
9J2rjGmpinPIthbYwnxiqfn+X0MsFL2ayXrBxrmnD0n4HaLNtzP8gbOjV+vuVqOkk9soC+rTFnTy
65L+QBPw/oeyRneMhV/MjqXi/eej8r18igfzV9NTejoAt3F4qL/mDq5jLPdulaljanekcNqLCukL
c1yqkQP1wZPHl2B1oB3QT4DhhFLRob+5C0Or3MLFMYwtncNHx4n6ZSJSlwBVtcwisfLVNBd5YSZg
PQFsmhXVeUW7BwgK9Fc/r4wmQMVkaburP0z3RCtkg2fbWHZQNKng3B/EEyYs73ilRIE2ftzNPG2A
H4ujjjPAIrv8GjHnaVajwbg4YUlIpARW950oKGGcySORf6q95RB58H+8k9Q8Cijc3QP66JlblyHB
RAJiqF5kRnNSS37rP3SWzcctpFcScbl77vgPaibodBriXzqSxCMn2vGsoJTTmf0xkKPHMN4nTz2N
O2tJCtzi1sEH/ehXTpyMxyMGQp3W3tG5rPFwvg6ArjR7WxGyGboUzBlH248zfwBMMR+Rl+4sve3v
5vYXMb1/Kmg/Kiet4dtjLsVZrvCOcDfQVsElKgjjeyRI4C4Ehrp8RtnyNxQw+kzZzZBDXqdrVWUE
J3Xf8tTsOeu3yI8m9SCYxxbXo6qdUUM1Fg7GdjfIfRcwVX21CYKPkBmfEQFwjLoiDb/hY0gzK6Vu
345szIaiSqSBTMab2cqi+1by2zOuB63GRJLAPcQ3vmDTjXzEBuZyHXlLFO8IuWZsDvqZzFWNrK4u
ptNZmhw/DbzU57I3xpqRknDFRpXKp77YjauiLeMgBrrfhSJa7DQfN/OjPrkGoI479zCAD5sLhv3N
QG8vOrZVqJtWwuGS4/ZD45PJoDqDD6dlpfikdBUyMZ/6rQNH1kN+HR5zvkv65n0eQ1N5MoG3oq6C
Hc1TnAaX4wXr6ARKDrcEOVMbCfT3gmyVczljYxdjxKtVNpyw2YJ7C3U2hXKBQJDpqq9ve1Kjc8T6
HDygd0RpJEq7By7aHszG/3qMY1lrk6VGYb+jHH40078i89kaiqa07nhNWw7JuLN5TPXMoHlFSr2i
WbbpiqdSAXYdXqz0crSvZh9AiEuTkq+eLeWpqeQULbjG0Rc0vUcAXiZZsyxjRNZDvMGWgZbFAijH
zM6oNWeyfK74fEdqmDy6dsoZzU8M0UtZZmOsetrCh3rVqxd/DZ9xdZkL6/2e1d5ExXWbeLr0xs6P
q5vLnhWinXCS4FhPi4X6oyUCdpKMZVXNqaX4n/ajK9guG0Rx3rqP8gF5paf0TKZgMGkRrYcEd8iP
VMMwdscap2/YJPlPpIdYsEwKNHC+4jFAFocHhqHc/kbq4neuFjRbSnpODSOY6AiDhHqZVfuE05ot
IwI8RW4nidTeVplzvTQWAWJ1vMdK4T2OZi7U0NIxx7QB54GgX2PwAas16rIwNsYoa8jI9jVh4M01
AbxASaxOldVMdTYl7UBeCfFMtgE0mwkqoNWGy7tRNyyk6BdRczLNv9+RMqBzaZPjv/elSlFjSY6x
NUN4+QLBRclj+PS/GnNr9gunyq+7BPk0A8f9fXXpiGGXfH2qoP3/HfjRTaUCVEBH14peUJ59E7t/
nl3na/wC/YCZnu3zW4k0vQt+zwI6vZZEGJcNPueRh5cNgRLcmmb0mjX9WEtsFsQM80Zs6ozcMztY
8TkH3Z/7b2Q3MLKYZ+qiXryaiFzyIRzDXdyMNug3nS34soyCwzsBDviQz0znFOlgGNaOn+l5bWat
ERVHe/1wDa0zWQuq5poVoP9EMuxCTZAcpa75WtUkt2T3f0To+p73uyfTfLCfjL6lA61PGwvnioCT
i3xOF1MK6YSNU7TGDMQAeQLNWb7jWI/pbyKoVC/UlVMDhJWpZixtHT+d9DXTF2/1IdvzpBGLtOcf
muHgIdgELRfWgyWQahieqiIA1jHINQuYTj7YsCd5w/qD1Zxr5KMfo1rL/ZjrygkMBuH/Pszhr8ee
z73NZuA12A6IiPc4eSAyw3xlBUcECFAL47V1Ks0dMOAdicRBwPn9k5p1jBzBw0KeElnPv/LkddwJ
Pv6xumISPQJFDgf7wET1s8w0lT0DKoa2cnjFGldAiqGAvV8SGcbspUtFna+V4cp1lgheacE2aizF
OAIy/oDqmVwdO5HXJrWTAa8jiZ0W6XZguLK0x/CSmzZapcnHt2QhH0tHLXPwOHmwVFetlaa8n0pO
nruS2wQMJJQIuHCDtgipFJPoDepkde1jwTZ1/IgOxSGrEyao8U1ze0FO4OGe5FD+s7LhvXMS44f7
7MvqhmXRxVVuahvn65qqRoTMFKW0rV+CkcwLIrKoZDPahEVrMBY/z4drNURZOu8Fbf9I/pYtjtaK
lg5BbAo8RSoy1CDzlQb8KBNXE/It4M2WwXntuqyZER1URa6BOhoR703cVHEWtEyoaSktLvGBA4rx
nWf4OcKCYPqhCIK0O5jDwiVF0ha1G0M+15eNFFxXk9qlra42fJ34FHGDsHcXaBzpu0nUlmFyXz40
LQIU5vg5XqNFh+Hr/Ha7Xi0/LTHVoQxnzxtrBpp16Vkw7oM0l/r276roNno/mH4bCHFQ1/dPKaF5
snGNid7uK+7jXiUHeuaTajiK2SD+eBjAZmkjvdh6CHK8p0Wyr3pYmRPXtxf0i0jWJgJK3PjZevoO
J7vY6iB5xtR8z5WRqrU7glAis2yBZcPoftnuFQZXuakViLeSFmHqVzTFQkZzfLOfGqzrYR7n2O2d
2L0Egv3pnmRd2920FYwBs5uy+pgEETWMbPxivF0d6dIcdmjRBkzUbPRRe1wLI/DdtNWYur3dRMwx
bpgYxbB/MAnZcsd84qsObcVHznLhF2RKpN1r6tfUTAvAdEfHvTfB7NQ+0/IM5gM4oQvIAKr0I+xf
ZIAcQKqSTZOqj3YY+04/VPs6raiD36vHWLgbOTSl9d9Ql5jMTtrt9hTCCtqBTc977IkOlmp5gmvw
EMoAjGJaZzccEpWXXAmZ7iBcSl5Em0tXNZetU2a9dgk++LWL/n8kbXos6dLZt4H6gtRUejlGWlRA
eFJXQGzf7gLQ4uDCydGnufVPxdvz9YK7bY6tIzueHAmBmDvgbEc+1HRCoKlnPDT1/RwrIG865/QX
lHbPvWqqbdqtd9ciIZwL34b30ipMguVQFrd+gRPZmdLcdTDOVwZYVtwDYUZjPdvm0zE8FUdqY2PO
Mr0rqT69VkMkWEr2kJdTf9xwjbHwLNV2OIFqcG+qpTkilmMGq9SMtyYmvQoiSrrB7VW5evZWPaiu
ovPZsMqqo2fIKeF066yLNec7V8IG01QkGLr+WlCugTBpUbLJCLlyWP4abFlVkyzKy+Mas/h4cHzN
eBhqWsJGRPkYmSBog23qwu53LiLP2n6Ay306IqsZaRNJxcNyFEYRlWQipw2A1tiS5yH3gx3vO9aW
g7ogd4uC687gB7rHDf43RFjDw2HO1z0hx9/pXcVIJ+YxcaE0iyE/rNjZp9EVjoozqZ0DeHpqqjPg
Q3agsTvTcaZOV1Byn0c4VI+xTWRBNi9Lvkv/GjRuv9LGg3VlJtzyDnw+O/Grrp1kR0D4z64Jxt8t
71ct0ZJK4OEDLs0fLxRehkp9PiOSAxwKHWn9fYtB1SEd6J+St6JUAfI9KKyRDCvZnxak6mFAAk+K
DhkgSCwqf4PB2h4R1ppUPh57bnNpAvncDI7U77/hmqm1eQbdf96uL6/dSdeyujdo/U0ZoF+yITLI
SssE2A1m971sg3QvKUO4jX//wobtsFo/9avlFUvIhhR8EgyGo8IgA2YoYkQXcM64VJ1Ph8xn8J8O
vWHzJf0Tldfj0PsxUWQi+EjIB8IoIzerqRKkCAbCtEeM/3vMummcODFatQDq873qMDCI6aoBXSZ4
y3I2sr01jca0hQrQ/ObRk5H3ZjoRm/zw59zAyGEr7+r2jvoomCTgSremXbBcQjP6x/CtYrpI2VOj
klYLI4p7qCdzrq1P9WEcGw6uvIbRBUzl8Gk8sTJTw/9KySEPv88sVz8M0ihOhHSLC+mmsvsH/FQ7
fixJuOxNuFDeGJXtJOqwbH1zn7VyhfzzTzCs0fTphEVD1AyZfdnw7S7ykoXD+3Q3kD/+0h9DT4LJ
8lKB/J5Lb9YRx/781FEBeI7AjEdpDeFLiFVHyEzPAS5Zk8z1zbH2bjIZj5jKYL+x+dqGtfTJGhBA
zdsnHgkPkhgP+x+T5FFOwjcD8AJQyj+GVPGaX8Na4if4sDHuzPLsqbohtAEOQEE+koE0zNd/vutM
E+K/luHcEcbz1wuc1O6uCRvr08i3StudDKgA5d4I0B0D1/tXAKqDTIA9JzeaSVb3GXR39sk+Bvhw
ZkanfVdnWNFoHP7iJbkaLiwsbZXGvhDlgdeaOQDL9xjdSWZMPdhy5qpFijqJ4q09+oE/Rgj+lWUX
AJCklR0/j+KBlk8d0D93GiVHO9YJ+yKhTt8KZc6nl23r14Wns0NBTW+MBVzPt053OeoGI+qMJs4X
9J6DK4pSvbjv0f/5PJ166pxPHqVyK1GtFKOI35xHx2P46KgzdD2F+TC/gKTKYfYcMZRIEcm6pnWY
EkKEeVzPk3i2u7/+o5N+yVhcbzZD0kIx+94ncS7GgZZzfd2RaX9+qM3vuHJkbBsDBHvUM/WvEorB
a3nteT+0uaDXdx1R92yZG87idQ0mu8t4s+BhawrwjbTvuCHDdGpvPiahNPxFcgwaUsWc44qiibSX
pRljsIJQC1JycERsLjTTe6gP7D3r1jzr5sKL/eXhm6TlVvv0Qad6OKBBY+g897ogdJXAgXCcDuYG
L+8tZaHQ/BncRC4SLBWoS/BKT87q0JaxRQcNeq9/HF1h3kCNGMksDk8jnzpq3ZovSE8hQUHUWK1d
ugQ1hCiJdDcLCKJh8y1oq0eWTWNreCB0geCM+R2bKCcT2uvkBg+pIzOb0wuwhFj/0kYaRLoMl2tX
KU2pZ8x96wkfz4CDV7G6h0mDgBPmuG+hJ7stn9ZVtHue1mYXxPQTIt+U0+bZ2XY3OWYZs15Nnoj6
9R6gqf8HAn+I7DmXUUvT43pZvfsngJZdETeRAz1IMDsA1K8+V4WtuTXZUsxXk708HnxxRzZxhUkA
IjA+w9yKeD26OZyCMzoKEJqrCe91M/fN450zLPCFB+n/Wdxm2PFIr36DQ7TjQEFbhxY8z6Qwy7Rw
tzEBRpWMRx1coCksr75FWe7y+BJBe6XMeqQ/60avScyPYLk2b1+yML25uLZtBbs79J9B8+U8FE28
WCPqaZo4ZfuqSaYIxLt/9OW21qfjTwvxIX+LIJWzIA5NE9WDKRuoYzEkQp/rxHuFRRqEf5y52MvH
wGXwmWm1xaZB2jyvGiQgpouOEpRx61iYghHGhXkgAZn+3jMy4KL8qE9Ehg08ia5mLMrn7kuvpJjz
avd24ntFGspZT3LwFDw7/gjTxVZttU/+nLbzN91qLvjH8+vOQNLE/Xh8rADKAWPnJf7an1N3IXDk
WYGkfpmdlT8paOAOS4E//EoRIK4pnPq0eYhl/PGxGBWN0244lQGFMKFfK+lm0j0hgxkbU63xaCCv
X9w64oYhBirpzufbOHv90b3mJm5J66LYJxf3ClR93lUElzHAADtidwUePuu57RtVXfNz24l1MwE5
UKgWD1FnhCCopR8wxCzY/DIUS7mpm6G+Vtqk8jMRK9obp09G+Fk2vsIK4dA84LnJZbt6ZwkqCjGU
ISdWnan4Hl1mm2kqCus+pY8pfB+p7Iog73GYh3SDwoX5AXsl0X3xy1r/cpckzfBvJV3ZqQdcRV3s
LSFYPE8I6wbp++ebPVzsINKxmvwqxIWOOrqPdjgFlYiexoMaeszRXebeofFZM8Y3kCKlSEgN+30K
qwqOSSF6UN97Dt6IsODEQbx8ZjxmyD9kIO87FwmqhgPiahs5GDbCVfQ2aZ5MtzLk6j6wT2+lIwif
Dqu+/CJ/ayub+hoWVzPUwdy/5vXHn58Z4Sy7QxgbtqJhZvOblFZpgnn5xLAz5pjq2YWsS+WgWdWD
wG+nWjnJQVLkDOHURAuCYvBsBkXXykIk5u+kfOqYq9xKa5dAXll0JFcBDC0EzuXw5lowGrdrLR89
N9sUvYFYqWuqggK7ZPWj31TvLnUMwftJam/ST8tXhcl3aE2DaI7SLbR0poEtrVb2h4jRNzSSoc6D
rOZztJg3bSDlxZiF9noT6Wt3lGZ5ZqorV9CB1WYPIXSmY34nAZ7KhQsrN/BLc1/iX9RoO/UUlvRa
/YZHW0mcO2F2glFuH9pBi4IuRXe44mvMaV1Qc0RCvVZUsRI1JwJ9rRw3M5/zKAmKxs2Mx5AEkcF9
WsQ/HItdOvNQyNRkUs0n1e982XO/BCFT8kihc25Jb5yyG3anV1WqA8ywHS+hT/uO7hqUemSUBfqq
CYMjOR9DetPAefObmtXR0ObSCkhbNTRKAh+Mf+swE0fnBoJZK33ZlDiENBWwZdw1viGkcDbFUKBs
ftlDBHljU/viNCEt2H4oi6gb5P4ebNtaPrYZAHva5h7ZnFztfXJsesa3EaA3EJ9r9fFIhutCPDDm
mvNi1SzPBly3JSPglxq0DNwrGzrUYnJPsN1DPMX1IkH4dIGxaMCWpkrWehyhG8UoVEabg8Gys9RO
FNgphTXJEjK6WJZSs3ZtEXoDvzS78KcYlrCKzGquUTMnpCqyeMccHw6Fn0VMerE3vkclmDx0YswM
sDcy944jfXWDwYvwLZuBpmb6ycUQwyZX8mkjSopO1AvJqxdD9das4SHh4d63jPgHFXSYKJVUDeAy
f5nNdMPfaZMIpwSeLufqaxXsCwMfI+YMXYByoEurzoPcCeQPpL1NhAAYM+lYtqUT8fyW5vsGLYUA
Uqa5FfXqfypouU9GbKQGLs2yte+6eZ/SNFDL0nHLQS2rQmHSGhQwglrkq6QsLYPSmTdzjL4sMxSi
CHqlEXx8Y2y05me+gwO8RihNRD3gSl1zsWTLkWGUfzG+w6rGoQowrRHT/Aa1GqJiEM41kBARlP1t
w1isHI630bVPImIT1pmZhraPBHWGih2NeUJY3n9dYeVyq3yfsImLYUs42Il7BE2k2WG3A8Z5flxj
7G/NLk/bkpIGo6cbHQnIngOzRVa54ODUAopMtv+s3HPdEFjXIKQwA8tgGBNuR199t7VZ7tmxAbJr
VdWrpbwVApA5lmzuQv1kwu/LSBIObqtmICWKPhK0M4CZmyqqjXurDD2/lYcJTqGD28qYTTDldgMg
zPjiN/paL3s06B+BhUNSqwlkiWH+wOSDKR90lrvD/MTIlnurYt+gLTfNOdO8xh4Rivqy03vYaiN5
pFguByyqCD0xjG7I/2dFWOcHatZa994KYABIPivq1fTwEyMPtz2fbPcSL6WpZGTWisk7GM602D8A
dCQST+8yleiEfiFi7MmWlbWM3SbFFbUWakuooBI/ZlGpLCrg9OyxX5FJ8bWxrVZTDkM2lxr8R3dD
LWdrkp+scFNqPMEY5Twu8/E/BE4IeqA8cG/Od+vboN/DpgH3oE/UV1vkubeMeKH+UGkjMeMHqrRc
LwnhcD8JYQmJW4UU1CMwf2Fq5TM60CWZa3EJNZW+Z4O2ifq3+1PCY5GkbAAdyAR36Vjc5fI7t/h/
34hSY3guqnTNlWVdmWDMii1JSsluESctZIE5XJeoEM9PdoVTgaPwDC1gRORHslkJX95KYaEb1/k3
phI7Zr8NzDv1So4pyzJsPcso7izwnf9XS3Z0ivFL7l+WNtKbJ5lMhAzPGG6oF7P5KBjG+wKDbn9t
bEds0fWKJ19hPLoBtYLywY99HY9cmb67V0u790XnXg5pRaqwJ2HDeT5Sgd7RB2p/NrlXTDkabQcJ
sGnuipXYbIjOkvBxI46dbY5eVJkRAlelC3duGkjAZ720KSUeDav2FBsLasuZGVz9C38Tydh2dPEU
x381KC3fTmH/76qrh4JM52/iucBzIegA2z6Rhym5/EsZqgkvzND7MwubI/oVrzFp7t/mYGdekigM
oQYLOV1z5Y2j3vD0GYNmR1cfEfMYs5I0JT0z+fPd4i74TmopFJKVIvuJr+nWEzN0oNAtpKWRkGUM
58N6Tx2my19BKus/YXIL89JUu5SP+XnTmf4OA1h2+zKpuFlyVvqgSauSgY4ikw7vdHea3iN6bzx7
W9aMK88kAUo8zTgyuqt38mynP5JCPRI4V/DHENdWhvG22bXm6Fo4Ax6+jzRpN3BcTG63v6QqJaIf
fvZCtrCo2N6CWmqjovCQp4Om7lLitqwA+0KvN/b6c+kKQambnSDQB0NvO7YD/JwMVyon2MBko24Z
eCFiUaghGkYlJzyvWAVNA8/CJP5PVKNPxc1TxZnCOcV7U1wtYGWDnII/JWUutacpqvSu+Zzcz9HA
hQymlV42tXPb49jBtM/v4C4TwiHXgFar1fTdMIPf1/BnOTI2+umZd3/ecHOB2/rGyZhzxOHpPKt5
XPn1sLLDsqhQRzk4iYZsN7zCiJxkjN8NPGEXh1dBY+ihhywwuTDDbSx4jfmdcbmQHCXyrGLZ28u8
JtdEIYEtCG9ezK91p8Sn8ghYnsQn6JHxcWvgrzPZtq1PFUiaiQG9h+oW3c9W1SXILvirL4ydQ8hI
wDhdDsTggAxolCnWR2ePCryT3zaMqxCznfe8HEBY0zbyhGf3Ex1CwWVs2X0sxcPdCmFdqunoza5D
0hu3Y37T9XxpdJswbQmeFcOLvkys9HedXViCreIgJCWPGbgGhI2S8qoSh6kLA47UL1v/jtqGS/c6
X/kCmwuAktkwYvoK25CgG7YuXcbZBbI/rPt0LL5UHl9ZU9vi+fYH5Yv3uKoVJoG5B0qOTkBX7zeA
GUGb1/b8J5hdarQ7sDGpikvBk5Z1ug2EgSJg6+PcDQQJJckAu91x76kVLCZvA99ov8xJ9HpVJmmH
mUGXw0Z98OVyK387ToB7avRry12D7eD2a3TL8fr9UCXV7eDN2CIQFK+SfGoDnu+CFRUlexPWEjMp
mhU96W5tt3hzYT7mdhvjPrLQ0gaG5jR9kC8L2chj6TDTJoaHdHtUoxujXL1ymwoAsevp40MfL9YU
6d1xEtiIPZ7S2VrncwGpo637Dc32xuMukS24EgOIMKAxz4LBtInOFE2VHqaB71LXHjVtFVJjpKSp
7V+9oS4A+E+UxSejPsLWbinhvDG9zG8c+K5K5CwIz+MJJzbwK3HPXgjd6b4ICTggLxfkmwTvBDRm
LQHaBmCGHO/MXb22Nv9IUH5BBZmVXYGcP8aSJ/jugD6pTzrUR10Rml1JrQaNs0eh1Qs5Nv/ixb+K
OHJumUlDfyJ/+aZS8kYoCp1pm34As/jvlTD9pjY0pWxT7cjuhP0rSMFaA6OwnUDL69vT/anhR0uy
LVMDb4ak2zR/N+1hp3mz3Qsa50aNv3l4T1aLMA5N0slhpzzEY9lEvktJwj3RZ5ceCG4GGDhxWvLQ
kU+61Cwo26ROABXOufajl3G7N74bSQMGyQfZlf606aSd6tni0DxHNAbU4na+nET0rupC4NZkfZt3
sp3erwQJ2hBcA1gSB63V04hMig+teAhayzAAImBC+qr7TD7BbsbhzZ0UgzAs9/VgjwsMc4MDEePZ
+ZLP86Q99nZm7Zqv6Bektp3AO2vjNvRLtfuUBzpxziDsHPYowyd+x6IUTZs8l0DAzsxrS8QJQNDu
RlJTGTxKxELt/WmExsa3vZZV9PjQzqUQCbcs9FQfepS8y9+9aeBteDtklz1HkRbTu03yUNN0DYoa
WiIFhJozrCVPsFUQqzN7jsFGMocONDk1/HBSVhGDPnCUiuhDivD4YP49Tpt9pYHcXyHjxM5OhAk/
hKogusXC9Xz6xmY2Sw5NvdquF+J5LQQJAov8n+IDXXXDJrsAm5TQQhbZC/LNtONdd4Fr5ve1DS50
DEdRGtT/nUGS3Wsq7X632gyhzMg0huNhgvv095fhiXhmPV6f9s5xGuqMdbheDQufh93EQz2n75Mr
X2JWl5cJMHGRIMCmYwOSa5OcpF4wMzhitu40Vw9b/KGFBvGwNKlBSN2rSbzzcIJabLr5kE/NbJW+
QNk/0NUhwO69zdA+/DGQcuo4no2fYaoYNWBBNLRaqh+yI7anO5qu/v2KrHNCPdKULv+4ZP6PGStm
7z3cIDLG2pCJYVTADOSRUR8mY7S+yUiizHUXzvf03q/p4M8NbJdE2pM+GhV5zIiCRRs62MrXBAyD
lhK2uRRajtnccy3aUvWWEAWDBscEb3jmHe/V5pw8ZjePon1cf867K0ACCcPqslS6VCl8IK7uj0OS
qNvK0Y94qWaQuNbec/g6+jAr/4cLCrHf5TeOUWCjgPHkvQjiBIBd1HtqSmibBDCuWt/oKXPKqbk7
bf5vBwHrPrWojbDqZkKYz8bM4RTFDdEdEGMqwtebTI6TD1AanmL+b8g48l/OGIATIOPVTmUF4oRl
O/H1OW+HlEUL+JsWvS+TodACxfjUkPCj+8r9clZuSrX8TKIeGFqFsbeKRUxCc5JJaqq8k15/3rGw
B2bikz7+9fq4NTGeYectSFq8el4tbAzb4NlkxgV2U5QvKY2er21/w7S2wUnr2CvtAtTfjKRMxgUz
r7ql4RTYlU8ajkLVoGlSWKJKyjTx0sfOenEra9vZFHCJSLE/62xj8Gip6veDim5aC9SI6fmyUutp
KkSmIRJyEv8wt7tdoNMGsVHZv00yGsHUs0mlG5whDmRFsD1JwcrP+GCj0bE8PIen7584KFVbvoBn
/uwAKqGNSKyP0MlgWj2/KrucP/gibZUj9c8Rj6DhXtjjuyDHzFCSrhWU36Dc9wgdUJCBEVkapJGN
8Nf8teBqf9UQcDPss5GoTHEzTkSSKHEyJ+bPThiwJKDosFpgRpCw7vPceXJnNOv28x26VOiEguFo
rv6qO2qAz3Ut6ExXNcmq4SIW5RodRg38yg7ALsgvvZAATkNrGYC5mHyPDWAkSUQSYWGpXwsxtT6q
jFKAQCqbQmIAn6bcHsfxfUxaFk0LfltyOFIdD5mRDxAbyLPzs5JDVDb3SqWJCt7pHeFEuDIRL3FU
/m76QraLurc06OFyEJI3cbFKvVMFOv/ScNALk2D6w4duv3Jb1EJNu9mL2KWOhi23JT48rmHtAR4e
smWFghlXntlV4iiS6vA9Bhm1JwQm4P2Yq1OTiquwQq/qrszR0/vj2XtCJG7k6MBOqBk8mZCHsVO6
IW27G9Y2A/cPEtnhDB+y/VlIqn2v9uz8VO9ECC5fJTIBt207u1eu3g7pXNaSzkfejzReVHyotZnY
tTvxhetbpB6emvENsQocWYCjTSnSSgKBFAfsLpJ6AwldqYwi79JUGakOxnRL5KeGpltbmG/Z5UNX
samsyJZLWcOiSIaGOT/GmK1uEq0fh7CWROBiQX5/B1oTdbJ5wJoJ5Dhv6smtB2amKGOVqTNr0QQs
RjCI9BlJSza3kVjh3fx9Wo7GIA3RaT6a5Fz/L9h4wFLZye5PgtM/tVZrkawoIvOkwYYHKx1VKve9
TDAg4LjwoXF/lG4AMLPg22rIikQueXdpeD5YfcgBbButTd5I2lmJUxYwqbW3A6nr61+TNcxQ7pCs
wfOxI6Q/rgFoiyfnsKQXAo75HX/PVqojam6WguhU7CGoOI5D6SDjcDMd8ny52qERgB+RaN6Ie/s9
NwV5Bh4HC/6ZkI6DWCzZ++ELhYLxymPQSIszE1nl9kZ65K6+uclIQvWZNk4nUN8eVQdsEUd4KuDI
LUAmCoMXKbkJc1WKzfI/Xlt2IVBO08sR30//fjh0gCkxN5rSHtBYrJA2pxYgA8DJTD4YhXJaU2sW
RUzL92f59GJg/HMpM21dBo4dgtIHOhw8AMToIS7gON9Rxswkd8NA0V3QT3+8Eu8FafoNF8jx2v31
IJbM5cNa320wDjZT6DsUbMqLYHgYC3H1C52Wh3vnsNGFmKU0dZMEegyugne7RxWx6M4h9UXPVFtS
+gf/kUhFCkKsgPchMeUTV5Gdt/OusAbe5EQ8nJmbeC6uYxEV+JCBQ0pA8fp8ApEz71fODgMIh1zT
z0oESI7Jtl3Z6r8l+zGlCq+XZJNLUEfQc/qS0/Ga9kSRq694DZfHSn4QGNu9QUQe3sfj/QgdSV3L
LYKXUpVb9tZwXrCYGlqNczGzAiuQp949qE1oCBDt3JqFYiocSBb95pI91FIpXlNVgMR8sIBbF5i4
4fQuqVmQKEsDLUQRYX3P1Z5Y/kyBjEMbl91vkHnWDKeFNWSzCB/JitUNpWmixTRoK9no6qxE+Ntm
5tzaXINh7d43DVKQz2vwfmkk8QlC8BP1XT/Pit5fl9DijZ16drUp24QmnGorHQJrRqsT0vN12oIz
5q78o2ozPtIWooI65ni3k+nDky51jgiyqyMoY52mJonjdK/sAvi/T25IbFZ5/vYEgu+uMqMqwDK2
UOQTpyAaRyAqFNN4pd427/3k9GjEkl6bztsjP+g9TM5kSDLL87GNaeaUkcGbE9Wz9I3BLEMzNhgH
0h7i24XLfruD1GuiZ5WCp3BWgCYZVLw48Ri7v/c/hlmploDx35U91FBWPt/lT3tZVv/2e/hY+xF1
xXHAqLhy3zf5P/pLKK1gepzRNezxCd6kZTLYn0+p4HNOywoNIAT55Ti+IX01GbCnIyMjoD+F8P72
Ol7Siu2CiI5tfUPZXT5wem2jpfcXTr2FViIulSpV9BLrLsTq/eD7vCnDXulsyPr2HsDv2gmPMMnk
0RfYGWdSKQrFUnKbePjHETVm1ZWF4HMmOFF1PYLPHaH5Llb9fnAfFEfPeqrPDzYfDv7bWE0Q/niV
Hi810XMyaAFRDDknVnGYFYe7Cy/OwF4BSom0ZxfIj3EnKNw3MP+6OXdj+0TfyJt+AEQgnVUUiSOU
8v8O1WFD+rVUiDBMB4Aevx0mizpmFpWhMJ5aYjUNB+2pZ4ZXI9Fc37c0lhHZ8+a/zY3oNFkZb+3L
0a7waArK+7p4g2ODdQqSGtow9e8kMaKCNS3NIweag3lcPudRSblaFpXXpHwKEAWl+H2LZBq4BmoZ
kSzxV77CfxgHai9wMhjcEt7sF08rIOvONDyygOkxUGSaDpb1mJLxAmQ9sfiNgMD/9+Vs+w5sLjJ/
Hp57yF5XLq86Tv9reuKDyS+SSPqadK6luKRSV0a4qQLI0cGQ96dB4EpbApENJEcFIAe3BfbMZK6o
SzdAoDRWPu6EpdNEphjO1mnDEFQDYuLbuIXog0fPnIba6ua/HVUnXCFjQjfo+T2VxLYTiI5lekhb
typq4tQ2YtzmkwUaomR30jIx5Q6FS+9mBdhTRDoL9FQi0ufnkOxrfw/SQhzg6D25e6pwU5YFgQyG
1tzyXaiMHr7UgB9xx8qaNHcxuCRipXfuOotLE4nczoVsryHk0XyV9Ghkx3hVBbQILbQrdUTc9G0c
CDktA6c1T0FveDhaS+8q7HewMbA5WJaUB8NRHbfVzTTlFm2rqcV4oaPfUF68XFYwJLuysoqX0NQI
X4HUsZbcdDXLFJHTAQN9kazqrPd2/qIhcZA5GAAbnPvk4Le8lQLqbGouDMVV6PH+NhRTiSHeVRaZ
qeGVblMlsgEE3RxJ2YDkW+U/avi4Ln9kjtavvjJnexMJgXvPB0/eXTWQUG4Efp3MamFWmVRNTrNe
R+7r+QNp2wkA9NstSdsgBvwKl5798UwnmvoQwyyRtXAwmf4UAruPHjh+XhmqAEsYxLv5pVXJA0Kb
SR2AW+15p1YElZXO5PIWaQ3n7/MN30zAzlKM7/zRUJf40W+LZoRf8c94M0U7BiMGGDQTqzmPFLqd
5D8XXb9GIwTDXS5S4MeUQyzScZhb7N+OTwii6ruWxKfvae6WBnrqhux9ScruwKKp/CMFEfpJuSYW
mNzLhTpf0tsjamMB7poiwXGTs2u2elESqBpG+1/pc9vPrkIoBzQCnab9qCSkn09FjYUUBKTZSWI9
zb84/9SNLDAX/eAl/T8pNIaRmQkw6Nud13CsvVap5SiiJ3Vt8lQpOAB4Vr62A0I/UAjiZjeQeMWF
6PCLANT4ajv3roBw+QDTeW+/Xj7qhlZIX6Cd1qDnzwNIySMoGm9Qr41183iYM0DrQ0XqVdwTRBFe
IXqmiGEunuZtrCSNiXJ1giDrOPKjqgRhyxxdBtknLqxeblHeVx6k2zqgWQsl0OGOs7ijdAzT1fG5
3lXsm4I2HgehjmuVhv2G6Lt3zLODL/jIs8DVgaPnoY3YFg6Jwq+WSULHAWI8JMxCF20Ia1yak6yd
LqlpL8N8bM38iA8cmqWIJ6+KOBFKZBViIIMRHfOTd/kzyVt7y1t/pAeEbyQFnaiFBvbWfncxgZ3I
YVj2mhPHhiUQ1hS/1Uq9WUJaI3Jkf5HFCcLUuOZwstolPJldImyIJGvdagE3XxhcdhSmYHzlSQF2
y1kX40Em7MOilgjQMHEW5I4Ife7q7vd0Cotp3LDCPRtFDaElbUyuLJICd6eb1Q43kqq1PWWie+9A
8QyqhCN+YB5HxXKfwr0Iagl+7SiCiW0gJwk+59AYBO8JCK2fUqX/8/QyflICekokb0zGF8/tuiPE
mHfS3ySptmPtNfNp0YI7Uf8frucpLgvwyOU73tZJrAH+3F8FUOlO4sIEZYcCYYVfUd8IVvKebBd6
FQ/gTNqEYAPKYUMoYo03X6fnmG5kZFEZitc0MAol1go5pNQvfpPBQughT5EV/+YBv9j/jLj/b9cR
LVkMZ7OPmC2rQsJpHc4/S2r3uliUNOXn/MpEENKcnyxrYUYILf4V7zgMwpUeUU/MVK6Q+DhVukDJ
NkEd4nSIQroGyUWF2VY6FElZHUvxhIjoQNURNY3kCQ82ja06dAGwgcUyCj1uteWpc4SEJT3tdfEU
5mCmRf24qLdOYv3f96IB+I1NMuOP0Fm/ul7Je26roNPNAe0SQTgblA2+DxcaA2vO8MoGfQyyyb4L
YJYCp0M+sNdrOva132yqz5PBrG0uK4RR75tAEjpo65AU6maRSxBPF1kNHHQXTNDTLpF2SPjiHmVn
3zxK61M4Noh6hwp3ZSBkQPROTLGhsTawv1HUcQ0LF+uMtPxWz/Njn7F4xd1u1T0OFN20yVdb5DMF
nzLCMBq0xWZID5Boh9sDuyorqIKNmwThDINQENvH3UrC4X9zPxBf+hsxQ8RKpp+6Rqy/e8YDfkbO
UXcOHyA6G5xm0cekV34lHCDURXnao6D0x6zN8d2s66b71xtleXvIbdU8t4Qwo5yapFa9Qed9m33E
4335ANuDAvSjEpgQcVb95vqjBf/oLev0T2dt8HTaQL0pp6HEcl1qup6HYT1mmdP7eIALYfOBT8Ki
02iUcVCgm1tYJAW1VrCvMIwBxbxbW6Jd/T0R6jrNiuSS59JM3Irf9xxbFX9sGPI14j918Mu7fNo1
vFNBhI1gg9/UyXcomEJCBCrBBLAdXKpk29l3+Ab9qcu8Ke4dTUXymjk4+gnoeamoI8qUyi0Rk44i
ePc8j9J5PFLY3avol8dhks3SSiecwE2ZhGxrIHK81U9b/Ey/9KEhjTFi+AAyiTsb74DM1fcrspvN
2EffFQCVvFXVMjSJLO7WIkZOguJ6FLDIRIT+E7cQebrxw6GszO0GjAlXHq/omXZbes9Q0D/fFebW
/fuuVJyaRy0N41aRFqfhjSZwEe7srNXtoKHPnKueccETAFtsOAsHdwAiwNX4cnrN3KLq0cnqKApV
zEGBOT7IFDUamol2uoPa+iCAzw0k46eyWhlvYzbWzIjlwFDfUfwNtbvlmW0bVgFsEqsSemZ+95yA
/QqrKbn08d4jYQvOW6AMRneZJwvqqUg7fkeJ9LPJh73m778Zc8jbDDglVDyAkf1PZov+j2mZuswt
98KPeLZZGnADCjrZLQP+0mDbLZcl6YvbGJNEvHJPYKnHiWhU+Ggu2RXEgoxY+1EkfXQ9vPqEpsaW
EOomKWMyFpeLVFb1EZo90ZrkGK89znPVkCieYN0rIAjopwf/hugUOS+1FDuJK1A6seKh+bvtlSF9
5f8BIhTLX6EXztDm6Hc1V0QZrqlox7aUtNJoRmyx8rsDKPU2HvwglJ4vz2rDfpll61+jQ4HR5C82
CE8dboctzxmVJ2yiePUWGlxHXirKc67gjCjyaiB8D/udNHrRkZ7WUXC5lB4GhoI7IOY4m6L3ylhn
YbRh/nnoq51CLCQKH71aiGn2N556PHAbxKdJoFTetY/0u/bo8SuLbnz1wnEVhaWdcgGO21tDkBZZ
AjmB9WMWzx8JYTRBBYTOg//mnBcU9/dBhUf20UQjzkihu/3j6tsx928ItZlWJrk3guhuHfHfHUuC
qaByldvsAqT3mHqGhlM83UGLv7XIMMzQUw5j8y59fuq2JWO3R36EDM2Pp/yxfkvACv3XxFOYWo9W
CM/+78P7Gnqc/4qruWBJQSbjQZv7dwpsfAUIcn0yX1twJBZ+g9ujWg6NmqTtpP28TBBpIOZ10PpY
lAKy+BxJZuduYUQGaPnApgOr4in8kKSaAVQpacyOnu2+JETpfzfqs+TvX3uTJCjNmhu7biPFsRc0
ccORKKpNwb8D+QQRz9ZXqyNoYp39JnX0TFOndb6Fw809fgdmYUiQHXJ2lLiFb/00FzOwf4YDzcIz
2Ak5ClYglIX8QZztueUzQ/CBewiFFHCqN85DxWvbbGzAcawo4vFI7GAVMcsib127Cq01ZrFRY8n5
U+ovypUKYbedPGEdPY7WKLv4WHN4YCbIRt21UY9rasvvE64kqNVdMCKGG568OrMdUafKVNAtL7wv
il46G/GbKTLAf3wtSyluoLySrXqHqYn9zOfYrFDhYxv9K/cr/dprMC20tRIa4sAoR2hV3iRFd3Bf
CvkuFdKTu5ZRRr6R4Itcp66qubzqBoliJmpR5l+HzuVnA0AxVeN1lLVtxE0YRUtaegrsAYoq8pBP
Ju9u7gD1hD69DFKLagNWclCBUPi8cS/SAGCX48gtCGfm5/ydKyuIwB0msk7eNWVZr3om2h5aBXML
SZ/eTTyACRbeSqSwP6wDdx5+iKBnWfCyKmJmiW0HR/gv6h+l0uXLqTyTxi4mOtZpkHVuq9Fruur7
lOLF7W2sZlNm15QInvKX/GPT1PmbmWQ/h7J5nYIBlGlt7dO6u908awUkOMU6qr5vK7C/xiZzcJQI
obgHDcQLI4Z3euQi69wPGLeZOU6bHTAwUGQRxKw03V2Xi7+kOo7Yxw7vnaDZz4JLqbiJXXmj6s+7
T7kG/C+ooEwxOTDDWtRNDExCNP3UbUPK0jzX4zfDLs0lTzTPtZG8XuM3deqjjAD05nsksVjLjBqj
84IFXl8Xih63jLvcKuDY15S60YBzRbcyPoZ7anKGnkZZsEcSahe1JkfzjRk82WXkodRe4KNfSCPZ
8JkCbQOw5Xj9Ibm6RuraO2e8pL6qb2LfYhrhzI9rYA+H2da8CbbwiFDRLfhFHsGUK7LQXgIVp2R6
MEYzA2z1DWaEjQkRiKJ7iV87bPjFK7x3CvSgRAS/quipjq2UOhv2eKZiswwyot9NcTruOeZElpKk
BZbh+coXbHbHqt6JtpaF165F/eBDAQLBrgrW857/CZCDLtS6kgQVlyMjBdn/1V7GKJbJow6Lm/UQ
g1n0ueiLKtikrLgQKaR2vER41jawoyzot5Fz7lrrzaUuUHwSnv3x1jMawofYquS7nxe4bkBGG1v6
1KwSEw606zkP1TyE0RTKl0SFdM9XnCJ2TplzibLUp8fEMu+BTtDy7WWANwLSSzlSvXwwE4JJ/+xp
WfTM8tAOTo5PFAD5qrco5dxwnRMWvb+aCCHIITWe83pD//XC6tEIkYM+8py8/LJ7iORuW/Cdlqx0
os5F45BNLzIq1Pq5VwQ1dv0VhqqiDQ+XxcV1vN9ljT1d0n7b3xvoodx6VDdq0KfdXKzMVf/Ujlp5
xbvRXDw2x+B1zAyHFgYA1FGiW7uwRw+ODvR+tkBEKNDvAVLwFDWp5s+YOhlCnXdKpE7n8Xzye6l5
QIxHm6TZARg6mas/j6A3ySxIifAS1bSfpviHy3q3ck6pavGh7WY7FjfkjwuEEy8pDYBcOdIfbGh0
BKJeC3KjovKpTtx4or6ea+fTqfKL8iFSCNgEQArbJgjDIuzhwvXZyrrimKFu3kRarN/5t+d/8Cti
eirjqQEARkd/b9/N0+hc7T1ay3QHFBcf+uffqAZe1l+S4ZwxGeGLq67LhluwEx0pvxFoIilygqPe
GptxID1pPFJ6Ij0xtAbRE7GwMss2Z25lQixmF/VvBNmHHHrxdbZEhsDkT6lc2RwVA50I1duUSL/v
H57pp7ZKC9q/EI+MgEcINVrvGlbReskLBHBIP8k/301SO5uJaSnbmqRqp2u2OIdBe5SiPv8e0POD
uyyoYOM3rhRJ1BKtG0QJ+YUm9/8dwB0PyfpMaKZlJO0+GnGVa6PgmVqGYl7tw+Rre0MqexIr9lin
WzDnL7Dwg+AEQi5uNHZS1YM/FAxAk9pT54H2udklPDZr7PEaLpD9Dhel1BDaBTLxfWecX//U88Be
Su9jhoKZrEfmy0EjPmpyg01QhmuXYx4pYCiYdPBdcF+drG12yYCG2mT2GaMMxWcc3kvotjSSlBgu
SP28CqMMTvlnlRvGavf/nZ59gUmG70yOml8rI7YWG+xuAOFwLyvKYuWSMdJrPzB9V8JieUg4YgBU
Iwdciy1xW0rFBd6yrWUEp6YXcWK9Ku5hujPW27Fy1govngr+GF/7+aQwEk8Bfp4uE+tcMoh+MFc9
XjsN7/Ly2I0c6jzzEO73mTfXmjpaoaUPbfNI+0R31f20Mx0C45Gg6Cjjo1CJeAMDDx3Qk+FYSuQD
Zi06xBpcdVt4DkP6d2EFEK9gr4Hv4D/tJSwXIpFU+aosnwu9/PzPwtKw54eUhzCUKgj6E7RGu0aB
mPdeTH4Ipmf2bcKO2JTMYkYZqQs10Zx7capBE7AvX/LzZtMGW1eRNzDHRgi6m0c3lCKkw5jyzxnr
VayWCXQG/SdPFI3sG+E3NOHHxAW8UxI2WR69g8rS7SfMpLobU+HuWeWOGWIPCzMBva5nYD5jDrEo
vzp9wDZQKk5rMqVME8ixjitX0h2uq3hc+BNop8uYWNEurqjDVN0OAPglaCs2xgsWJWF9F9faxo3d
QFA557f9/RXBBy3rSyZa7ruI0Nr6Jvn/pvIkOPJc41F5eTks4Hb+yN8FEF6rrwzm7L8Ozo5G/muq
8SRHjMDQfaasuqt2qfWnYjDnjNUb0dbMOsafXvu82NjnLwWljJpZMzAJuduWDhR4bY8aYLErkcem
QdOhI4rdI4DGdoy+LEoc9eA5Bw3mId/YVcJcvZ69AnJxK8nU8x5LRat2oHyFw4oWq+9Yz1wbUX/n
gT0+e5mYzalyCvLFEGCztKKAMmoiO30x/ZeXCn1+uB64REsUe1uByO+4mzAlg/V0j5ivIMeJ4Nhc
pKO4NfNhuWe5B5g1MUtGnkZacRj+yleUNjyI2A8wsjk/i6GtDRDH+ReXhL91bOuFhmPrLMYhUV+C
pP7Y664LK+bTnYTtqtOxyOrUU+Hwhn2oqUSh4KCxyGHR/1aiAAEmBaoJ6PV5EzLSbBUyBEO51IVO
RQGYkPn1ic9SyExgBVPZuE6UrTBrMsvi0CWlq0Ol6aoP5UhHxLEhKsAoj2na0tDuz9D/6pVxdUHz
ss2ArO6zbJOngB1TkWZor9v9Ug4iuF30xG8KIQx806CwjsopJuZM0Uww3GCPRXMHkQP2a4QTy3o+
EDkW7nsRo6enS2NXHljxNXH3z+u9ormCbdVd6FruIjRK2Tx5/LBFKWMfF7vLn8g6YQzPjj+rKiO6
RRHTn98WRcg3NhF7PIu8ac991H6w4TKdcux9MoMfS6+lt2GXYV67e8G7FbtaqLntnFTDBlcyt+Qr
M5rMve4bXo82NHHXgJ5tkTwl2ScSXNUG83kj0d8S6aGC+2pxWSTze0z/191dK5bCR61pdrJJUz9z
qhzd1HCqxOKz3XTEWPx52LGOKOhAogJzJC5ejUB4V4r0XiZvZN36T6ZUvqnde6BVbfMzV1bQVJjC
Y3H1HikEIjCnrQ488WARYKTRZ+RM1AHNe0tGFGss+VPMjsU1XtMwjRqnrCQnjNj0EpX0RV5yM10V
Ms75GVrEuKdkftt30FjbKcaIHrzS4bvgTo285RN4n1iOjG2r8hN4IJGGlZkTp89HG5BcO5F6Bm7Q
EQ3fhsnhAcLACwtdO8FYHhyiP9IVsGWSx0NBZdL0edFMl3n075pyDOVrrs5v3GOJFBWgOimOcCfu
Vt8Uypddo+dEqkpSwxRO8qePYYmpbHE6dmZIhMgeRz/58C6I8wBAt/P9CdAGYQggekP+7vUtjenk
jBLTcWSlNJmy6EhlrrfH62NMoC1lQnpGvD29RR7UA5qDu9p6vheJpECAEPeQ2JLmnbn7k+H43H+M
PsO/tsX0XpKoxwnbl1wa36r7FQlS9WUIkkVakxDup/a0vr/GTXCbB4Ti6RfqS8PZY8HymA9QPWeX
bzXBB/Du6QU0nSdCbPbFpS5ito+HsZrWmM08qpjD/8KUIRI9ANdNhi7oP3zxaC+5KWSZEluNSYNJ
hmi0amKxQ8Lvc4fxMtLOGPO4Gk7tpYXGu8XvxBh/cOiYiJVUei3/DvSTB6Zc1Zzsl3L4sDH0OL2m
NRy2hShuKHWeOzAm79uENrtvF58LpT2wf+/Tme/eFGbvLaxgVwlazL7lvYDjB0lm7Hy/bIYP8C3t
bBtgwWHRqOTajiAQRiRWEObOhTun2fEeZP7X2rhQJpPkmEcgBzw5pf/EWM7b82KASzNXt47S68Mu
+0KFq2DZJfPR/gCZpd5aJaqindzJy0ZNI7bksi/lD/H+DaSIu9MvAOie1ve+B0hY48cY0yJAwZNh
p9opnnU8smv8eB3Ydb/pR+UUFJ61frA/VdzpIeHTg74LbIhwOA2wyDRlyhiYg9WKzEejZgVvTCXS
BtNxnqfwu4ffgG76zMGvIKxHBAhQUXwkXgPNzKIP9j7y3iND3xY4ZId3jTVPsvFF2ykKdy14jvRR
Wy8n742P2NHTWNm0BjWN09e70IcZs14MgfjPaH64Ey1TBa8caRwZ87JAKTy1isOd6o+ukyWNhPPi
sK0SA0cC+JL8e0VE5EY6xYtmRDKE7b96/QyNTdevGuQu2imFl59C4ReSG6EqhSm3imsZhiBdWEgj
drBS/MlEOqvSWf2UKCVXknHo1pCFYY9fKsIm4SnjC7hjYimUgNt2y5+UUamOrJu9cm17WDi8GGAx
a/xZuhZZ+dyUPY/h2uGi9yI/eX0CQ6gHIOXjggvDy+TUa6tAEwGag84vauCjttpZOiWkonxZyg7I
r3qud2RHH2fePM1BErjw+HKUWGMz84Q1WZJeMf12IwkN3lzkmBviMIGXcPB7mmy8X/evBpwTJS1m
/AEnbCrstvCEdp3lhKQq9UTO2umAdvH/HDKTC/6HNJXi11utIq3tc1Gvbu4NpkMQG99ZQDDDWvHq
hDlyRGEAx1Ibxr/Fc4bKjHckHyJvK2yR7QFrRwvkWncw5urwcI55UPm1+PZJ4T+ug1abgEyUQ27p
2z/LTMIOqdriwRVI/4IKR9Buad4ZzcCMmOlyc5SaF1iRpwoqnRpTZ9NSPn05YVrtoDWNBCdDAjRF
0IOP7ofYGy4rOTF4Nk+CMebgu19ZadfiEss4CpAJWuDpn+B906oVBYp+M7QOZOZg9LoTxvINHQs/
FZfyTLpeKdxyGm5hTxb/nvSEztphwr1qCvx4uPEiv/AevyvcTTYQUfctkmejTXzYK67fV+yRze8b
bnQzne8qL/vjCzoUV0LGCDK7aN2w8dLvGZJ7pFKEp/5Udt3Sf8K9l73tZjBERYsBfVm7yGGU8eNX
8RpxhfQsJC2yPSwZyNjMVs0YInj3Bnp+NzsD9bTdx4gnVSvSgxlv2DrPugVYFeVm6S/cwT/66RVc
sKe2TofFLwO8kcURm2Ly17XjR3whgCPj3Y/B9ps6HaeijglzGXOvl4SqtY/UJfamu5zdp/uNit0I
D1rU0RVW+NsOXg+vXQ8IR24er7cV+iNhoyYVmECQb7mEwEMV/GSGfCkUJrJvxWaLZAbwYS3GwEd5
9gE085+O12l5UJNHRE/8cI/ZLamqVgtyrL/93su7ueiUBcCTAJXRLvfMfOcY2B1lDoUshfkGVeTx
J1OAgqj2fAlidVnys976cJ1zj7HG1PgYPscAFa4zYixXpQTsCB+4wubZvSRroaiz9D1xcCKVF5K/
yzxcX6i+Y418c1M8qXTBi0hQlHKHdaRw14Aeg5zbbU4RXYcKz7wieG99BkBVIAY+Zs+B6dYbxJGJ
xR68VahO7CLq84Npc5KZhobZGrd3TN0Q2iOzNk0/w5oBs9/LAgH9smPqVtFsh0dwVjsqb6OavW9j
usXujYLXXwx14Eyto++fCS35eJ5kGgFbt65Qen93l3ek4ZNdRqdIw3NdXBSPc8RWFe4QaNQfSUoY
XB2sJKWxIUe2/NjtOhhxZcA/DPM1GE+eLpr411a5LYO0f35gNOM2oXeq3aYTVfjNSVI3unpHnJk7
ikgZEh1R8onxJ9xyEUHPXELHd12eYusruNI33sUZ3lDZWq7zFO6ExsrtvDdnB4H9r9g7uinYfRGj
hUkqijM59vGEBiw+Y7uzzxp5Tc4/Cmu5iLOJp32x91EVboN6GSIKOuArjL/GoWEd0+j/K4PmaNyW
vJO0pE2mc9Ml6ZGnL0fuxoz+XoqP0psRRgdZAz3zkbT+LykN0n0O95nRbNyJEVZaX/BGixkWcCxj
b0rZtBQ6TbwHNW/cn2rIeMXwFCq5q9dfWWe4+Wsp3ztnfcMxih7gmR+cIUTMJ+l4KMgQ+4Jb73f0
OTfiYbW92J9YoFwP202FgbVixQ2ouBDMrsRt5MnWMh2ld/mxBRgNKBLFrGHxonl8yw6Umr1X9uqy
KbJcmU7DxusWDzEjy7GFrEeoH3fXIckA3gTXqX+YvkzKbI9VUerLC71DlmX/5P13krfapaPJabGl
oeDZtuhvqAYrFymYVJELD+YKGJFsbHEZeOgcb12hgWCMWs996VD9nIuz4H9RvPWBbRsd5mlaXwMs
lvnSdpAbyfSvr/GGJthBYbXv2s+J3WtN7KFMMPI4pG2Pk5qkXzNG5h0gUqHjakJsnFz1bXv5kN0X
2lFHMurQ0f8R/SHwfi7UYQcIk4pnMqj8Izl3tzzAl+94vQFsRInhZAyJf9kVia6SIm1x+Qnv3Qt6
oteYwj3RC9xlLCbokfboWMTb0HAxcc9JWt5LiyIfh4XV+7ryzNZYJiWHxgUPmPmMw4bntnMjJjPq
M38uwTDzUhjyYCWDuMhpU3tbcQnhgbERpCcRJ6W/XIhOcLXnc26puJvl+ZeRUXtQcBMSOQMul1VK
oNRtXOWtfRUxnupslWKVl1cVQsIY9ChtcYuBfpnS3vFJPAApAlGnHwzCIlJ9NEX+YdQlN1btS4hh
Xlvj60yyU0Zns7e9BHDk2F5F7cwUV+ZdeX9tmTuhekZCmHfRLQFxFRK3VfMy8PZ5P2i/9cEl4OYm
8277i1XYWDMnhoVfifreUM3ZuW8tj7B++Xrz6LgwhRvdo67vkSXHuilbbf+eQLxJKpm9F8waXkVw
tqRBry2IuOGrS06O5CKNreDSXdDvfvDCADx/EAJVNXIHkyPsKfTCMAI/scJ3kxrnJSE8xZHLa31O
El4wQvNzitlCxVMunhh6RDhd7C05R1b5hxftj4e1M5XPh3YLhNqGkje92UmjzmKNO9LApH7ZwSYi
2eoMSZyOe+6D4SiSgXx7UfA+9QsHXkszLxRTBDAw27/3AVzTdnHwT9lGk6uwBaxNUpZGuhULdvzg
ZTPJ6IkdybIpy1PUIB1GxxMz6YLZzvqSi2hJDSXu4q1/bcjx39pKPO4EyQVJZsM7ojtvUlWExeop
juOKMVo2lrnSOMZR16tMCZEXPV9/zmj8Di17/xh3plOHHDNOyhEDZKqSKNhTC38hbBNIEHWOjHy0
/sX+HqYs3VJtcRdYcSEpdkVdwhbck14iPCoRMsp/df1ipoxdJK5wMh4vnfiqRRZ0F/rpJxu/YIWd
F5rhmZFCwVWT/IZ7rBpBJiec8o7K8nlbkaRqXzG8BQIDVpwnvSd0rt70bFw0vbwTSIrgvRjyTKqd
hcRjU2ruVL8I+6YR8PVRnvsZ+CdLA6onWkOO8q3GtX2YmALJhr3eOE1nxTubrRjgFV0R6g6z+lRi
j2y9SGpF1o0Uyg+uYVVRk03fuQfQ+4Sou982kDF91bohUosS0G6O7hLafsW+WCcF1PsbEOabm9NB
7CPGBZeel2Il/l3BcjS01nwX3egzsKY9q4xhZIdNiwvWVLxeXyk2nwjeS5MLAiN6AyB6RmseDipQ
J68HhnUtD5QpHUNlfuCcCEiaz5AyNxRyVcjRBZ/O+zqflnpn6hB0D8p/ng/W+oJFcuMW7HK0yd2u
Qg/7ndipe9A3JXjCu7pzs24GVYfxWeHXmYdLhHZ6O9X+ZUnc0W5rNXQCfkbVP1ZzGE6cQDjMymcy
/5qqNv8b9n0BksWAh1fZh/r+qojO/pH8F5urLL6aCLV97OrqkVWsoWiyxNQKtJBiLG/OSWkEYcbE
EI40SczIsvxuJYAJQPK/TyO/haO/dx0Roz/Gnz2QKxAV7mO+nE5pVzW6OYA1l99I2hLfJhbMLbZX
mTmv+NjKKX+2AJlM5egSFLjFuvHRX90RvfiKU0vCPYuVT8ZZzMEKLqxvFHUwfWtvVNzx+Eodymiw
dRG0EYTvQP10yvasqfupSR0f6yFJp92v/Unpneg0oUlwjZfzUsM6L1Rdt++GzVj/Cf60hn0S4xii
5VVqIVnzuOjLwEiN/bDVPhpfc+mLTmLMIJu5iYu5wPGZuLnHKINzsGPOE2YUTFQghxXG9oI16pqG
FYcW5ba7NWDU7oixjqEnk3ZlM7sfL5u1dU4hCw0j6znU5YyzDXoHr/HVXjF91ySmooV7fLQAgtsx
IeLCrm6oeusd6/t8cv/gYYt95jS5JCFoFNyxZNPDBUAYt/QRWJO+CejoYy8wpRxI1nnsmacw5wB+
biz9xVQTk2gG3tpvNhG2SuPkpSlTKYvOH7pyzll9ysj+fh5rmf4re/DQ/M2WLEqrImidOGV6Q2Ez
j5y8bE+lzwuIlI3m+qfwZw4s/IJ79lTLWhL1FJNELzb3Ojd9NgSRH+GCkVv9yx5hg2XBOKZD+cBs
aE9wPmkd8XteCiXWa+VIGqkmv1OTx7ChiA0RToTFA0gFKeIrg5obUq/O06KCdNsIBpJz7xaioIRg
7ZopsAWuEtsl/acJCEXx9oc8lpglqv8bmZwhhViIKrA750RXw2RnZJCM/VSgoJLInt/UCj3hLn6f
dNJtDsg4V4+AqaAB5u9c7qbj9XKWVgGNw/QEdLwi14p+uRaZhCWjXby2QRkDncoDNzWRdm5cmbhU
O+g+eUwCJDnhJ8s+17DLOx5OqtkEHQ6sYpy0OGUXGs4b3KC/ICN000N1WWap1tk0lyGn1fXmYYv0
M2EnJL54EMzP+5B9SWGHqOaYsD7mARtpxz285LbzRQ/DODIQvJi/jWZapmsPqk4NIyWYymNSDFS0
5DcQvw/fblj7giAZYpSiuBLBhig02o8sqLSwyvI/Y77GwF4OTYLyPz9JfmNwI3ZQ+VxJnKVE85Ty
nkUXjrb+GF9a+1pimAsideayxvzF8fyOYHxL57PzMb4V/w5jEwuwapPigqt2/V6aejxHpVZZyyWu
dQ5DhcbuBJAHqOujHIJ4lLLtGyKon4F2FZOv1L3HSat4h9zErdv9bk1C4S0KJoS9BFZ3iKHabccY
oUfkBG+b8rpBRIusl3pFM3oHPc91QMR86hukKxxOX/+Ovli9CvxcnJkwmGnrtCwCmXXrw0FixfhJ
6f8wk17NT47Taw2VApQd9TEb1RcHMEL9oaqOlAGK4itHot9jEDfHBT0BmoP3oIZ8Z4mqQCDxqWKo
Kbn0wyprwf72gvcAOxEi5oTbmUpLJwD5+j/BSbApOBCnX+N31S+R3hNQRBKT3RebciHzhrPx+Puc
M7k6M+jNBaB8Npsrx+1FKKYhVsd1SZnMqPNjWA2BrMwE4oKKj0l5ZpTXtgcHRGcK5I6qhPdQD7ow
9oANsn1YB1Xjcdy0IvcCCL53r0Kiq7w1oDRVb1724ceKANFibpbitkVvzml6QirbizwM4CgXdoT+
dfXDiBBE12UIcVkvPKsXF+I0rWTxvIYo8lE3TxY9dX98qEjmWODVmU3nRwDMsLE2Lc7J9is7k1un
L6RpwUk4Tm1nvIjgvK+D0U8qtr6lUQZj/jo69MM5krMYhJs/qZv96j38nSx1J3HtwBFrch3wK6r7
gx1yz6AS7mrXoUnaJQ0yPPd9OVYLJGCq7OMtL8JjHrB82SJgE9HvIJMmPnyhtYLsvC652hXULmrk
FeBnOFl2w/wpyC7b503At6ihWPX66O2eGwXHBZeKmSxO6Bxq7+eiQtuWvKmTMo0oUL8uez3hV6M/
i3Fh5tRlpSjNisFCW1X2NWIxw1pN+GWXq7lql72OhuO5YZr/74jtISMG+hsbNpfrxF55p2FdNBjZ
RtuZK0ZAxLULRlT1u3phKBLTI1Djpc74w6C7bjBpopMzUqZ6xcY+Ed8UszePvF1SGIRAl+bRaYBm
EojPi8w+Gz473HxZ0Fi7PrmKzSjEA/MtMkaM5zr1Kan7oIjn53hUjQ5hRTYAeF9cS1SXLLQYG1/m
xzjUpoIn53y9++j2hh2+SmZlyChvN6YbNWMlvP/hykH1O542UP1MJRi0bt7QJw0KF69fhT69vqX1
UIL7BeIXdbqm4owCYbFc4ZqZd5JW3H3ZpaYtyerbzewRlJ8yoNBz67gosS6HWV5jArhQQvoSzxk1
0FMdR8GtSpOzB5i1qSEu/tdjWkuQuZlLxVGGI+WrSJttYfMAup339bUooTywR16PNwA/oYmRXze9
ns1QkNVNs+ePW3JIEfAfOgv/L138o1KWRaYk7dLH1jL7SPg5u5czDFZGd6WaaL6pRJOQI7T9jMvA
wwjni2OdDUNOooFfy2iinIUlgjnYInr7qXK2ol0tCMxneHIVbOvaP3t5ez0w1E7/TMNmjQRw9LP0
3GIkKt5HkIqnQjJun4jQ8ruEWc5JT7y9RiOzpQKMXBGA9t/oz04/vpcfOPCmoFgKxEtpOPJfWCNM
/zqSedbwbxOKUk0I2JH43mMww5P1ID7gYu55nvtf8xMIhFuW12iY03xBUHLyaUKpD1bF2CgUZxLs
aIuAX179qJHP7lKi6eO1Eb6v9J/EGKSQclXoUEwI2LDx5hOahozghjsOOPlRrdHY9GRVaiu4P8Eb
k0uZiy6BhNHNbYk499zY2mfcFNXJiHmnNVcf+VbTcjN0mrvvstYJ0Dte5f8ZbH2I8xRkNLIkRQ0A
99yx/505/h0wCoQkZYkymDLcOLarwS5xwlEjISgt5s4Hcqc01IXbhRuwsMe6wnTGrtm9CZ0lgjxf
tybyhEKgOzb0/rnGdnFkAJl7z8hO1Ivg7Ejy9Ish+HWWi3qa7TFP35oEFYlVzt7tvxIEQxT0ZTF+
0HoJvds2Pktaecb6HYHTEV/q2BsgJ6H8RRFZWn9jfoAxS38Wyo2R/acWRqYRcaFXrwdQap/vjqus
gxOkLOzDsqUMSfKH1Ij2hVkXKZo3/dxDXlgLVqPyn02E1t+Hh7kGdx3de/JblZXV/HbujJpN+NuV
1zo0NCq6DBl0teSMSK1Je24jS6M+Kq/HA/Qz/6Ut4lMQrLl2Eh32iv0pmLHXnl3knT/xpc0kHAZf
4wf/vRrODbR9xvgIAU2PwsoJKYi9ycmDtR/Zn/ip61dk+ArNW0cehB/I8QTooHjzhk5zPvLUO9Go
E34c1ZdpgUnWycASH8b2QvC4kfaGCPFqXTxszg1vF3wQgpka2u4jVEdL1/nk0HMzbeMYwXvNeEtZ
Y7nKpJegchd4iEAHjvGPoBwBQYa5vD/fyx1eLCyl3IHsx0Gi1Kn3l9dkI7MSwhSUiT+eN9DY0JKB
wqeYebJYmLxFI0aaPDeJ+4aFyUnoC5OLDgT3ERc8HQgTgTTwz6q/CnIc4oY7R2UE8sjk9hv3bHHp
Vc8ihvwtt4X8vZzwO1oDEf3oltguleTMDj7Szv3TepkYPZiYJKe59NcyDud2FVfxrJ90CAKjcS1u
mzc+Nro//ySYBPJns5lhtf8zBxXCvuJKDWi7dqOlZdAjaxXtvftUvqlf5D6l/wMTUBG3hRkvAXsx
qIwJEsd/5EVxDiKA+4z5lamBR9gSSZviVlQfmdHXkVkRDNi9xdKb2oMU7JKmwg2zdAKDGM7x2KGf
LprGpQ34FH7gLfvp050pC6f+v7OxzCz9xwm9d1M6D9Y12A3AJMqID4nHLH6DaBcNWbj/MqcrrLBJ
4hZ5ukEfZ8G+1DXChde7rDLHDv1BOPR9VMh248uwfCwhYLanyo8V8YpTv5uXl4gQ6nJOi48ITeto
35EEszLeY2iD1tygM+EoWOeGMlWLvPxTdOD1OU9IvqTdEbAgn+tRbLQkmJn56xD8HB/womqzcLkX
JeV+mIZo+2WBXj6KUqPWHOTs6kpxUkmKNIuLat8uZsTStK0xGzYdhwmeTjhW+qBo7YlvswRCCN1V
/760zQhg1RegbsVFMxs+LpoeTxkFtHYGaZIGa8ktO7L2ofcEhj9raQ71cULzpgsVfzV81IBZlBQs
M6kdDyTz04gbK+2+7fYf/PVLCdGMm9TsBhBclzDA6ExvarPGw8VGOC9/DIihzNWnIkR1lF8jSx8J
0rNO5AIP2M+ZAXJja+i/rTtK5zYdg2fe/f8qCtUR+CIY/mLMZmudbLPmTuprmkl2UYv6XA7EDJom
HlUBoyniW86reMZbD1UiqymSs4MUv0x1iN9j/PVHea8um28zXp5DliTKgAG2waEHT+CLYjGndM0V
A1ayKK2Wn4SgcvhnS4ebc2rpxrooinAn0S2Jf5m+BD/9EuxGW7a39wnDz/EDPX5oorM12rCYoCuC
UuQaMibZLIaxKEyPxlhFFC294OmF1XJtTA7hJHtyprN7Oh8YDbkdIp53ro0K0XJxZ1Zg8eycqnPz
RYZqiIx5DaFTZdXaLRAoYeEqCLa0X3hmtuPHEPCxerl3i2IOAFS9irHozkkta8vm9/69tteg4zdD
9vLNKsycrpVxU8I1BEWTFFT9vCBcC5b8LAW51vYe7wBcJr4e+YN1BdU8ij1H0gr+zf/bKlR0rBC1
ajXCPh8t2jN8bH92VnQ+AcInRwMBx97JZjD9pcQj1/25u8ycY8x6kFx3aw3uD04CfeSGAXqtD5fg
NOM7mMAljz0tAdH4OYI4BpQgigqNTdeI4pJP5ooKe3mDiILpccGfnupwwRh9CjqELgD9xgCxwxI9
75GMoCloMQo7Naa0nCJLGguMH1wOvGjD8B+fEUtXwHkLsCdd7B8vRhJF3GcoLd7Wzjv7iMGSWAHd
/sq3q3ycR9S0d3C6Z8idimrQMtdRffAY0ISRVR8XoCKVWcXWJa+gn/oKzdBOFfvBNC5UoQlLrGVZ
9mf0Wbm3p7S1rie2MQabGgs/19w/bDhd3tWv/kc4vaCyh9x26NtgvD7SHaPcRlh6mdbmf0akgF5r
WzNbBJLh5bGXVzRk5wo4jLaX1zsTUtLlxJRJ9lokyBMzSrkvgK3fxSRGS8Gsn6bE6umIue6XBqtX
umjiajm7FKylo5MbQdwliMhdMiMwbwPNMA6Aj9XdJq8pkm99q82PJqxYFhQ6vkC7yhX5NQiap/5s
/DIIOQRHWomxxS/CPAbf7sWGNeyeDJUl3SECKiapYmlVC6jn6b1GHMOlAa6C1fjl6LHZ/GwiaBh/
YLKFkWfqdZpEPQCbSFPQKYsy5jz7H89fCjoSqA5ocm+pXbFVTh2ELXraWqTrInfxVIoBnDogFShm
GWVxgzlMLM8Ts24CtGtgsYL6UOqXCjqYdevOsWz+4sAm3R9j7tlwTSXjtIT/43fzq+3qBTJT4r+T
0KhwH0VN1pPsCHj8W98mizYn1QM3KBrqlWxarwyAxAN8uBroGw4WgqWP5aJhf0LXI1nQ+8x21Ykc
ZCv9qqQnS8Wn7C0/8tPcbWm6ElC91Fte+MrYcDTefbzX9vdDTFC/JdDI3LZB8AnJysE+70wrJbi+
Ou9L5bvRNwBw9b5i2jTgXmHl0vgAslGIpd5voMLf8DB13oRWhSPtVICtdQYbagLPUQEP72XF5Oi7
et6U4aDKvDAV3cQJCNvIF8cyihJBotTgA8RGHwXsCLb8JE+t/E8bq8FleGUxj+7Pid5DHmFx5eK8
0+GKJ3Ez75AWtux085To7IHHOuguFhvy8J0gppU4/UO5foc5HWqYwqpYY3qgnaZeeOShLaElNbkK
vZnVu4Fsi0C1ZmBaesvfS9FfZWRdNscML/Afb1ObSUMH+RhCP0eOzATbwDff5na5HBpqeS34n9/U
CIm6es8yg92+7XazHqCSScXzXyTuOgCxMElgEM6DAA+6H0Cvewv9yJAHRY+Yx9+Dfwf4JK4Hvd4d
laV17ShkNlqvRC3CbuTNI4X+FxfpnNcHmK0sV3XxvSDRZWq+jFsstJrCPspgaL31FIj6/CG+nPbB
WYFSeLjjk4WVW9eEUeuA7MIOUSGm8faRS8xQB8nqM8CkSZ0sN0+3wSQjRH6j5a2rcTOXRexTFgno
DU4SNQvi1V8+alHRWLgHQRKKPTFmvC1rgCxncIQaGZ80oRYxIIGC+X800+hvhvDuC1z3AwEIP8sr
Rv1/nh4zZBMdcqNRGX9F1zmNFWgzpFR8//yaDho6CYLjYsfV/X0HpPtxJRMZ/hoO8GxI2PuRyhy3
9QmnTtMV4jNUHOsd59U5m9Gm9QQ8cG9LIp/QY8h1Nw1mz5TtSGUgkjHMyPS/3Y8RRpO8xDw1Eo6u
b07P65x2Ml6854TzPGogBIroJBnbI1AXNGdVaQm2je3MrsDpHKXlpZbde1tq2pW7n/RVh3ozia2f
qelCO/BJLRzZkKPBD57CLZ7Se8EpSwChL/1OPMJXR0PymtKcIKRIkDLxmkWC6ZZ2Viw9VA0oP0X9
/OeqtZbz4nMVv/goC521mYaEihrUYPtfD6yBpMW+pMKrgc9B2GZqVdYzVQorLpV+iiJMIyuOz/Gu
sob5I37mpdUZK0UAzCYsoOu0tiKfl2Ms5/U/d821AMlOtKtUPXNdVFLGO6CM8gw1BAE+OWL+pycQ
jwTr8fyDCYdt2LX5FbbbneEQDwvctZeGpIZX4cCAgwdiBcQdtPfjouAYI67P7LcK71Xgm3ygDk4t
b3QDyNntvr82rLK5jiIif4HW2ndwY7Gk78P5JGswq83Rp36wPo161U2iarBFgAW5DcqUHlnpxkba
1PrHeZxH/eFyZqZPTlf6fxw7BX2uLiAaWMBGcOaTmyzIWH/dDkg9fc9t1/zeT5k87jFzWSsofKGh
M5WDF5CmPL9xI94G0o6mgHHAweNP/UUvgdxh09CzVGCOkFp3kHUbyBK7ITCy3GGbMPkzPMz7YRB0
J41AWD2S3PGVhXdfsaiFXWcJkSw7We8P05Y+DSJSmhUyTpvSNgOfPu95gOM8I3+qFgIJCUUd1e0H
nawnA8Zb76wYXXDWaNpSnT+zfJZlcBzQochpmTqfDSnKFM4hIB/uEJKhOOseCu3Mt/RUZOq0Fmf9
F+RgioUTq6+NlesnT0N0xOCzk8BkScSAUVE7jD9HciGV4WsUbGWAqtricC3HEMLS/+lTSFKqghLE
gv8kmiz6WXjE450BwqcufQMxewjKJIIFCIMD+ve+jW96b71svB/t2m72H5NItFVABtBcnLTyfl0q
wNu1RGO9pK8px2fMSkvO9/q2yVP126shZr7kP24Zr66iCzkSupY5cV061k+mTFYemxojtBoRku3I
apYg+h1NZm2+cOd6gLDcjzus3m63OCJJRaUkuRtw12c6k+t6yMPQAYQXupafXVceqKYCfpn2RK10
w/Xq+sUBD0b+jhIr96Uwgj3xCCOBAsIJPWArGB7zMn+grbfiZtFjBhi+ptM4WWVhWywvuI2K8Eie
3D8ymPH2bEtEkVOFH8IZa59NKClafNSMqRhHsB8YNH3jNj1KGOiXtRIrg/qhIESeTVD7BxkIyFRH
2et/UByOL2siM2gGYZy8BVZdOX6lyR4iNmu0DJUQrkcZcU9r8flM2SdhsNBqFry5/O5SZmdYegxH
voAaCazhl6roKK/mkA7zbrS6+vkB+3dJOIARhAeRuNFTP8SBycjkcQIWlsV+X9YyoCTOOYLchVFv
Wrlp0sfshbB19p5Z/Cc63n7j52idaDs0/rxpM3kJePw5/NHTF0jNNmwfIDQfhzPm4o2FtG/fp5sd
rxwY/W04l3ZqqwogqdJCWVoCI3afu7nwSo3fNR3YJStLH+wAgDGvXuH3fBmhDyCSN4kbDtST0uhC
/NgHKlgkxE+AbX7Xv84sHXPNaXmvpyLQkxhw/EwVXAs0sdlTRuBTRRPAUK9E1HFYgc38PcMrSk6L
VA+2mpH++Tsjufa8piUPKSSp4ULUwqCyx/WWl4kXH6FKewicV0FTrPmuRLC8/NCb2dWi0VEwm/OA
43Z0ijdhMhIteChx1RXqydHD41/7niQ0lC/YvVr1jIGUs3tfyy7SJmr/Y65NcsW5WXBvN8e1LSrF
gS65hhiOpyc28ZFLM7N1dyPg3dQ7V3PKDvkFYZ0HVRmOD71c+hhrPBoE6bcScTy/+h8BLxGyM3Qy
w+MVVuOofXU0v/TPeP1aluxeTiKZ2LwhZIjzwz9j3puX2TLwC3dcxEq43NObMRp7tfvvCl4DLZZP
fzUdpxBnQFrm3w1GpcLCZ1aCRdYnuxbid0NMApjIKK9rECPFw0yxUn0B84Wy4CEEZ4gd06zouVwu
4M7vPRNsWHbaj+usUznKul5ZnCRhPzxjrn8ukxXFbFn2GL0z+j1eD188BMYjiLi28hcO7I7Jnjcb
5yLdYWYn26SG7BXC9RASWKC0UY8641C0i+GB2WqNNN6a4tH/zxDfUZ0FYBgL6L7JkdewN7OdvwiD
2YFBpmz4p//yfKyOy+C/FM2TRCmNEBAGq9JXwpggPPytR+b357oCeF9VTddks7p9yoaYFrFWvAwD
4jUrCB4NAuNCOdM2i3X3+fttzQlqqUwAnLYrCjlgVcQzBw4X4LtiMXbzzR2G5ni4hap6Up2gW88S
aF5zDG9oCbKBWynUVozD98eLdCfxevWMpkpo4lGApjj85p0qX9AvzYcmhpqsT7XGVADatEog6280
Vd810anQVmROwffE8qHoBf3v/4mtw3Sy3SscSqrxhr0i11VCM2SRXkeDeRKKnJxJWqFunXHtMQt8
yy9YB6U11V0RQ4pIZzXa1oCCEvuhSFmLPqWJ+MS2JSv6+a9p3MKIPxCOC0dXig5Vj5ZGzALMx5W5
KFondit02H82aF21lC9K6rW9nvq+IGcTlcoNjqFYo4K3aPLwMo8EbBeSFMUKbDDFM09yJdAMMJ9V
eurDvd651u96Y/irSug/01elLmiSG+UKCfvrlYGbJgsSdUlakEW9DYE4AnlM7m5S4xXRKIWq+TY/
sV4epAzdgYkng8VsR4xrYT6OoB84DlLLcJJZRelYOeqHHVWezwwJAnGLqHx0JCOO45GHkg33EC3H
3g6doYAowqGckq/Fku9X7LBZahcyC2RwAt0snT1IE0H0Kg2PMzaVEdS/Ql5UIgSTQZKAgTJSJfbX
aAiKX+f9/xV+ZZsP7wBCKVjrNGZ31n88FqrywQ2c1ySGX65hvfi5dgAr8OzonxJWTiCxwfI4fQah
XQrhi96C9utUwgToEcH+BJzUmumjCiukuBQ0zv0IGfTlsVLfwlxMlQDetTfwj7Mxw84rml1BoBbd
kUNbm4ub6cuLvW/8ivnz6LffCTULlpRSdpyrr4+0PJ6hZNpk/RViWz/NT86WkMeO4akAk5fH/HPU
/pZKAoRSu81CIhFwg5hqkRFruPQtqR0Pw3g40X2d0BDhsjemSPIvodbcb2sbqAhaA4ck2E7cQRED
9Lzk1kCH9d3x78Z9CDS/cqZJYlDZpClDGTE7TUV9bGqsXsiVnFy0IBDDUsblCBprABiwpsIDNoB1
ubF5SPMgZ5flq07TE8yZnjqz6c22+SHRnfZYt8waOkPtFy8vGZAnW2gvcEb2+jitE7wx+Jy9isD5
0xgAMKdj0iQFr8bhcelLTUF+spMQbBIgMwapR0WWYypfSIHWd5TS6kFuiYyAWExVwluTJwfihwXQ
J++ycF3iW/FPMz0Jlrec58AxAP5HHpDTnZMSdrv7NijRJ2vWX8m5iiyE3CGZlcUbmBOJD+blqEyo
lPSsGfpkEhx0IBwdYE0bQqzP6hW5cjuLqtbuZUK4/xJ28V/TKu64/0Z7LYkxwcKtb07o0Q7nYyZ6
1xvktZTzqA5I85GNpZuS//JqJ6vuLuK4ALDgnCFFQGTxDNxW3Y/8UCtfwjbYqHWWSA50kXXg5EiM
KMGqszkpsgDEjZUlI52i1viZBZNwT5t9vaUymSO5nsuzE5d9edC2W6LxbvXsSBcBOL0n/+DgWAiO
uLqrVJ6C7uQIyAuSm2cdeN0fo97kl6Fd0ey1SURiIfTSJ16orFUTASzuOk8LbPc8apLmwEQqjkqZ
NFq76OkKXD/8WBHL2IgL4JyWfF8HpSfFtRSyuOmqHVOaMNRiyROe1eHggHkLgri7BbCexWd8pbhi
L9AdP4SCuHQEEjwkM5nIQa2hK0QpAoYODapxGgyYE/g6s6XiVKJ/VDtpDffqcIVgl5NwCXrc+nXL
dTWmCealh4PckwqBsPAOIQYd/Nj5sUuGaZ+afZVr0WRX+nEYHU1g49TrTt2EdcwPwUEQKGmC8OKt
KJCiSbpEjpq/F/B4OoFni26mu/M/GJkn7EW7bgrFqFhitmfDSDB0DRCcJva+OOYSlWlWzBHn3QNm
lamYgDC3OFBa0lDJz7xgQvDJ2C2t40MvWtPypUT5/ZA9kclf7uJbch7Q0xtMrNa09RF2mMnJLeH/
EL6yqYd3xlKDneCKEJJ6hvnbwi/Jf01274Mf9kNLl1uYjCtC3k0XoMViwynLZDaL8NpYGNHmiITP
S3vlcbzSu1uF+vz8mdd06mQ+iZpD24Xjw4Fozrn8G0xEiIYdJG9Qu00jZON8cx7qNvfgpuIVHYWf
E4yQC1hBQgjfJIinksZSYpQFs2aRpLIquZu+sY53bYlygz43/LkSHxAV9tjMoRndtFmXxpITw9wB
lJGVYd377wWY+4hB4PpgE2rHblyAYheb8Z80vJERO/g/626cG1wf9sDVLvLC1SGe8mRvkvFUc8nG
zVEaResxgbJXkT3u36484RcS4yMWx8vbml9hlkeK1Fwjmsi4iyk6B8b5iMKMSWW7nvxVMTQjRkZh
7ffftToCMMpLnkOxAqvBU2Uf4bliOpSI+8XOMumkks1hh0qOodSEcm79GT4QmRA/i+nAFo4gsuak
98BME52EcA6qrzrDpNkOW+dynOwL+bDgfzLxzt/4wGj1VuvYeg+1NPXHPV0PFkSDPFrbL8J8NVoF
9FspP1NaRkGoNsxGI7sND+BkCrF7UqK6BMBpBVZkoEQO9INIp4Uy/m+tISw/6ooJ+6QfVKDTgiRN
OiCCdqLTmcd8jMXhJsXLxBVEkRyRn/vGXc87hA3EuYHxjKIds5SXnDv7B65Gvy2Yg7tBAGVC8m8u
ITCSTUYrhEbEjPrTk8fEnbiJjB2FDOIBpuOXfx6W4JxQWkv18mibmfAdinStriMFAKT8GzBMIYBd
48iGjInMlcJ5kdCeLYqcfwgtWFA7MLxUcibpd+qNQvoyrOp59BGjJjniAlS2w3x31gX/CkbWJ9RJ
xhs0DTe2zqDHDsB1ybeTQgFfwTfiRlLiG8hYNhgVKtQX7+AXeAlDwLaCZPHVrB+W0kfWkYnvHuVZ
H0PbGpEr7x7fHkGT3oFJCMac7GaGnYsLDBYiLWinA9igEXJXjZgIqQTLB/EVxsvqY0yxHMKIiRAe
a1+CpfSr5APmh9omlntRgsN8iyszDoy9NFAWqhZe3Os2WN5ctm1pii0tRi87ni5k05vCTkdRKMzU
5rNSV9Labapdl4qswRYwL8qiYAziTVhwyRNsrQ/rGUYxD5T0OWwweXIwVOmdDItXfUekhB6Eo6P6
DvcC7oN8FizOX+VYxWZH1V5Y0slYpclL6Y/MALGy9kkSBOgilPvEVL2werM/WHAo6PZJGK/X25Id
IMy2f+RxKcvijlOTXHFaD1032GdWXdmsgeHootPSzTKoFRljVcJpKcNiYCRVz5Z4oN581qT+O1cX
dUkO82RP9tdW9f6AgibPbqsIZo+fyD+mePjRYzDQzd/KoMdLJuaoQM/BhGnd2hxwuGjJ/w3UWrOo
YZoYqCHOu7U7Vu/wXbsHLiZudcMmFM0D2TwYmpZF5NEJfRzY3+B27yQhkwL714M43YNclkZrfqUq
0lC6wg0TKy/Tg64y7PF3fd/a33SwRa74oy8dGoC3UVA/tabp27Rxz5Tp9FYFGsPp6+PDO/SHZsex
29HV+ntvqNzN+uBDpvis52i1xcyzkTmxDc/LO59or3n3BK9HOM9gA8KeBQ3qGdo+/fqlVgHULqE4
N64Dsz3HJYDKR/o9BZKTn1QFbWpEEvMOVDmJX4OP8TdoOPNJwusRbDeD20WK2V4Gi+4g/UPvAa/T
Z4PmZB58bvHtOHujES3t2wVm7jAt+91rBJUMQQ9Rq/JMKaTyZfgtfDoC8KjsAwmzzx5DPr4ACqts
e6vdI8Ee0ssiD6goleoFmWJqrTnFHIX5X4+kgr332hTwKF+XG+WQK4QzkdZZCeYJiFZZwnYrYUVI
qbaeBqiOP+7EQS34uUDuZouWxB8HW+H3y8ravbShUBEA+OSy5Lz2skDjN4VxC7Kpjs/tA2vZPVJN
2Aq2zkPoQkWo/3OMWFvpjBmOVF2A9B5YAMG+sBk/eWyaz7R27KO6bejuivJPvuYc6PzgHGC78t5R
2HbBHXcTJ5UJz7SqVRvCAxavd+T6FPUmdVUrb70wQr1XaLFPw1ZkX90LzEwCGvLarBjzRXSB+PAl
LTnChVHJWk6AsIXf9LLS9U1t8uTDCkRilMsX4fzn/WZZwLQgZgZ69BqUb38iDxUMizP6GRrqE65G
8Pyc/OgRtNn1ZYpXsQyY8IpJ96gJIgYIQoG9tXeyYS9xD3fy5Lv2ln5kBlOvNAcG1iaxgOVBDC+i
rxgpUlYujSYSLErtiIWafaOdJemJkp2Ni/CGM+mu3gUvo18um4hJdYI6rSFQfK+6FLwRa4LMh7DW
LbevrmLE5KyNfW5bf4DIdMrYLovCI9gHOb6sD62WlmgHhnzum1K+EVm/tpzeh8lCSyiIag/eF8bz
tDcl3Z8ruD3epEkwEto3+NN///XXxLwsgzaVBqjEkXv0OJQWfA1QTmOsgJkpz49WI3s7rlTzw5qz
Gu2Mu0pdY062BgxweiCa98R5sM0wkBAS0fnhpa2OO7huJEY5LF64mcMPPkCJUoOxXfd2kMcs6kLK
6PVFE+EsoccoGUDJrQkVv7HGs+Sm6MKNNxVFL+tDvTk2IQ2sGYjxov8SepIhSU93Qpy71et3CIfw
SVfXno7plpqLaJebSUwrFKgSMrmSjY+2yh08mf/coaMeItCVYEdcH0vY44ir04LISdKl3qYU9ID4
rvmWCTR/nE4hv6MBliFVb1hBOkHEWrenYtb7R8kU8R+aexMKMaGXwg+zz+MTUcejJfw8Yn/YGQJw
dC44ylBKANaLIDGIHao8ZMEK47xtqbW7MrliYeTyYo1lpnpwrvf2zBPy8me0vpgVrJQ0DWdFYErH
ePZDgzCk+xnHBERaWEF7GnqAxCWOgPhyjjB7C45U9t57wlSHk36w8ZbMeHU7UfuCFgP27AGzxVsz
jQY1K2Rsj43/M+G+dI10VWpphLc4LZYCJofZqJz3Q0VlC99y3uPy0eikeycP9qQqIRrlWOvX0Q0a
YuO/c7qJXxnQ8UMT/cbEJO6+PKLzIlFVdw21qeKWijGVzNIqzBDUOmdpxsN2J1hoRoTFbr2A74SW
JdhxVU1DJd4TfQyBY2KQ3XW5R3gNQdBU5/dtuXIqEc50uzXso6B5Di40pLqFoEOJ7g7UBmBhkiSK
ZJMFnv2t8efGZJkj3SgIaViot2Jpnn7U5delgh3c/eTCnsWCjoGccBlnkq/dvnk0hm8HVq/Mk/8p
3yXy4YKya1AAY70X4zAPtSycdgm4bDeyDpz6fGGYQmhHD2Y1XKQeA41hIW5crmcqEIxtIOqw2Wag
+zTcuChUKLBKoE5fFs+ro8oECZJVkZZ5dkdtuNOavXTA9h2Z+JPP95vH4b4xvycOorKqSj0x063C
GwkGI11l7itzVxVrv+k8xSVeo0epOs89Cx9X+1Xn2rsj/T2u4cce0a1gCGiQKcYe8HzVTPIBm8HD
ewJTsi3yNAbOhpxvW0FN0gCi4BvzIoNBGX0l198oYhoco0GTys0UrcX4pMqAtY5ljj0X67/XnuNL
47ygSXlnSqLI88T6WDaddWA80mmn04XC6jvx5kRWOJhijmUu/lw604Ntyj/OA9Od1GTrFOwOM1Fy
nKccaM9aXzNn1XmSih8OCPrlgrd5lMa0BmOlvavHpj8i0/PqnLXzWZrWYlaCqKgjvHRUwSn5LODZ
U2nqYMR05jz4FUyfY+WS+YXMNNaqt7oKC6bk419XBrwPQp6E/LAwGc8x3GzfsjgQo2Amdf1cQdR+
8QxBXvb7AywXUg//vU7pOKKBQ3Ssn6sTVv1258/V08U5feOayp+ZLdUXXn5XqI4rEE1kNs44vKKh
SaGSiI7RNueKjYqNvsgxJJmeOFrhjq6a6/RF14vLo/IyxINeoT8lAkpbfUahFatJYJ7ZLxPk8LcZ
78DX8NVd7yAhyAV0ym2br+pJdWtyzn47gqy/6+UWixE9lFPn3wVUK9wLwhp3a47WpQTlLVCIcPXw
iLidJyAmi8ZRK2Sx18il1bO68yEdt4Hw1/ltqHPsLHd3iP/uaHUiA+URKyge0xe14ZDsQFWASit9
xbqZ2HYc/sVIP0XJGdVPbR8uAAh5lH/SZOsmb0MYe5zv75lfRuayt/Heiz784eHewrkifgivoq/N
+uxHA9RvMxfF2SAgmGUvIODg9np8As/rh95dic/aoSP4PuwaETcn9x/heLLxFQCCPF2oauGq96kc
XI3c9qAvMsz1Eqj2aIMJwQXIaLhS8A8IwRPOpshxc+X6yWtWRc3zj+fxFzLVHMhv0JwLBn3ml8n7
ulUi7euCFrA6dkotzCT8hDPObBB1TxLBi06gnEBZr5+LVMOIEaS7FvFX0YaemdATzhbECJMYnGlW
Jvg84eS99bOAOWOeLtyePzK4CzllUXOzWeFkMVtuvBxAHWyHrVaVaxv0Bw6yuWUD2Mnw05g6/SYB
AyOWGdq8QuxV1AomspzIZu1Oj8Y813oLp0qH0ELXWpWGtXzliGePCwp+JiJgg6G/IEQ3jwEvnfNH
e4zgwGVyNN9i5FqBdrnOwF14Rciv/h1Pls9AEBmisUFDxx30QF7fqb3yEi2HoMkXfl1TnHLHE8f6
8A2CEVef9pK2Mm6pYBWZ8R3jnA4f0GsbQOESQVDS58lVOxG/9+4dyKm9SQ4iLWcnZoVc/4iCM3cC
9jLMZMRSpr3tSeW6dvGv+LnaqD0rooaMbpbIhybz76mIz8I/WJ96N9AB74cjf4zFsJyISa7Pje7u
MpeVWRlRza69PH5h3OHrGhhD1Ns+UtYWgof1wZa9gLW8lQhNRDKCQNFQJwCO15lazr3iPRz0oHWz
TcPf6rgVjnq6v6Gj+1XQHYVtXeCnunmtFl0F9G7eIhh0TKmNSBmVXPY6h8PoOOkfrhQjKMFWI3gD
5vOxju/Frd9cwvORxmJ+TYXjP6rhavg8MtdT6AnEmMhviioAHJenNYo+cAu1tvk1OEAF/Dtz/o/l
djOSILj59RkZr8OwwJJ2cv/v179/+pr10qpZDRtvjFwOd0UZckeQX0vXSViDmnrXg8Mnvqm4kamZ
ES9zAq9LpsbMoYA0MIcxbwr1lIqIS4MMdgt1hcsZibEzLBPiBA+BG8F5+9ukqFnAkCfeHTuhsYjn
PNZqqtSGNQ6QkJcOcyWK11HdMDolpgqvfAQv0sXqAF35AUfUIKcVH6VJz1XRJK+G/eZkMoTTejg3
Ly2uURsKnm3cbglVWpR2TgSfm8yWtlgXx35YL9ndSrvE7+hbTiG76sMU34shAxts7G3Bq/Fa9iFB
uDzZeq/BEOQ9FLFG6OZtcXfLi7RG5PczA+7XekYVAoNS25OTXED7rreiVnL1fwfuYZ1KxY3ESExz
9mq/zk9H+9pBFimZvLUjZlCQXjdZJE5xvzqEisk/gZ4Fg/XJGLbqBwvMYISQlKsXArmmI9OKyrZR
fUtxdX9IF1Ua6lBiuWJ13qIfVN6Vs8DbzhPAZFyttdGn0G7K90XeGp/tVnsnFKeJzJLVhR+2jdYj
w0xebMPIRoq1wEeuANFyAKIZiXBhxJZZhhPx55ILivO/FqaCuwbRxwY8qBBNUPUHRGI4Pi9b+iNu
OTeHViT0krQROxU10yScQ0YrWPboqFp1l/LFm2kwtSiqRfyze2TCsF8VxavFmlzLdHIFTfd4MgbN
Nd6o4LXl6MLAN8s+mAMp3wjhjJgnu3EDxbViSaMj5QAdYZjoF9k2FqDaWSftZkM1FeKOD4x/NqmE
OXGtrdxNipMCcBqbWaq4TEctAZagjo8HOJd7vXuwRxUi7tePGW4x+pcP+LuCVpPwZL9NXvm2Jk6T
gbu9R5hVSmIRWUS6+1psG/m6jQt7PvXIZA/g/OrfH1HwnpvuxJm5TINXm1rT7/pAsxO1Za99uT68
QX6QYszfHv+IgM40h9lAKOOZOV7kv9VxiK29zCk/t7Hof7o3sufvomNjEY8avNZXpgEJDWP3rIGg
smDlNqm494Ws7FuLnrMZL+hjC+/YIOgOnhyWy6D1bGH7BipqXE2uQTAGifYisWr1wdQp9fp7raEa
C8Ww3oOGw1RMaA3Ailb+gpA0qEaD4O9iwhGBn+q/ofaYz0G10TAlNh5jkmWTDITpLowrAVauk/Km
8Vc8pgoIZbg1r+mUyzdemrPm6PEl38TrUz/44SjnnyNMnCoayohN9qaUPj2NfGVZSZ3TsNWibq8C
1iVdFG1orvfedtDpiBWVwvhntmu5t8FoNJV5oVTYvyTdJFv4ZbaDip09gOoZA8jH55+H//b6N82e
cinmBPr8EGooCbrgeRR/kv2Rf6ExwSVm9DbD2wtVxJnwrXR4b6w6sbpaO8NzyN1VC1BiIqpkeeqo
esbg/WBhI/LJgFUlvzt9JCmtU42UuO9insmz+++HZ3N70y1tWekzMn6sQprbNGOX4C7pJo78iFvC
3Stisc7L/1kDJ1p5F5kW8ohZ0jCm0WFJXxnveogZeV3i0LVQT2jgKBgxo2iqN+nXXUF+kEbuhDKV
LDOgyIyiSHZTtqGvt4lMn/Rz/pdaulZsEAmpBYa1U16d+oxymjCIWjFesLRKA9tB45sEc7W1Rlkw
QLXC19421IPR8XwwSZguvdgfQHwa9RHQfiiM4Nc+yGteMOrN58xVwCkm+OfittOO7HWT5FDWjxdL
AhRlO8aYSSmcNBwEwWeu3j3DUq1NpaOZYNs9qAmHZtFMKSlLJcLV++Db7UOSNZsxChZ7Xo81aIxe
J5pIcqJ1pmQxAFkVcUQgpH0wOHNUxF8qNkLap4cuU0vo/ON4vn2/vDwg+dkz8a2B20PfkMZzflAm
gT6ZA2THkZt5BCStyLbEbc9dRYuk34BTqpY0RTpigY5v2E1GLPPSG9hOzAxVWWRn1zNGqubVhRj3
Dl+RVd6Z7I3U1uikezZsyqi+qJw4VzUJsEmw1am61l0iCDgFIItdpqBnn/AfLQoQAHfVSR/zj9f0
o1EEZssDCwbxE0CGeWSSh+5ao+9Oy1owGDmmevl75DNgdxZiAhgVp/1RgXCB8/eE6tS5E2mlL9ri
YFlf+b+Bnfp2q8zrTa50K+4+3Rl70MNNZ9xRJfyyDEPzeEa8XNrCTyc78CcFZYnwukrgWn8+yf6c
4lBSYpsdbItqNxOJKq83iNrlbpX0h5NFiy6B0xlqphf0BJKyj+iOKLgT5QeimkJDnCLA59vKZFx9
IBhL/suYPmbrLd3QI6E1Zoz32YAJcnhmJnaM6LLvV1oWnVbRs85zyBBs3vTBuFiFLtEhYDawykQO
vNzzP5h49ILaE3RQSMSLCvI9pEjaa3kkhEiKjA8Nj/c8bs/uskDrzsyLWpto6Cjuj6ghwlkPhex6
cuTFF0zcmVwKIquzRvR6Fc2iAo7q9Ww1qY9eH+F3W6VFgPjgzYAUtEKnO5zdDzyN1Kuhm5/0whom
J3zn9L8qyDiZFjrwQdG4G58f++ij8IIKKPU6BMdqMZjBVoOOwIKvkdnYAOm5GjgcXHG7kOYpOxuI
mykfSYOuR5LrC4SoDTMtqTCNq71m06sWz26dcQGRIlpFEkB/+THEsBk21A2WG0NsV+4Y+A7IPRvK
g0wevAuqovX2KIflkKftrlmAyMQJIAGtE7E9G0zvEmO666OnHT6nyh2Xautzccv6CxVN4JbTLXFE
O7rZScf6Zr0JTDlkEvZg+F6aGCzJIRzqkRCd2DBCwu68vWX3ejPjgaFoXXOuDx5e7hRnDAnuGBqN
QMK/Z+7c3PKlEt5B3uQ4f3V+2DxputxS1rGlsjeJTJ5yz442z1Zhrqf0trYYAoMZ+bFVOqH6zxHN
w+1iqP5EQ78RaXylOr4YGXad1u41wwKFjq1u4OmqEy7MX3NihcF3OJXYgLVaIl3VGfw9nR8RQCyU
Q6sbTMVAwbpzOqBqKxH7Xevwl5Sz4dptEVjNRQfApLW5pNwvrClntQFN3cetwhhDC3VoAT7HSNPG
bWnLx869JtcHoqMN4DFtn+yu0fu2B7RHvK3P2k8PcLANit/33rHrBDLL7MQY/LNuvWIY+Hqy0L81
/aDy4qProfzr4y/6cWo+o0HEY/8hUR/QrVURGGKLX8wRe4ocyVyfObODLoNO9E5gehpp+/Loj4v5
2ueoYj/Aq8ogFIkiWZMWPZBl7xmTQdoidlnmr+uCNgYMUjhUZts+uSB/tllcRFg0epd8wFp+KgfN
LG9YhdGsNh4JHStxOcjIuWWWISsJlWgI9u82SA1WdUOF1z6Dz22xjx6G7iltifbAhyF3i8FJ7Xac
8Ss9B9PDIcJFhdLiuPt0HuFXi4seCXkDemXGT+6owHdO9C35xQGgT8UJGbmlHw8HJBGTdF2YcCAv
NBt/sBAZHfEuWISKbVKmfxycVbKyRDRWKyB1jhPC8FNaAPD9ZQCJUJZLrfb5Cc+o13UIkNb0R+iF
lyJF0AMyDfMM9rYpomKGqWKazi2DkKKvImwrQVScm4/5N5wgvOymNh4k5nuIcr+EB7PaA5Va595t
MhZ+jDpqw7oYUtiVrvbNxe5HuCVFtgeriIpNO2D7Dcnq9LezjElK7f3MB308h+6EpqlaqyQUCawD
7r14oh143FIvqPVpscQc2AmwF8YXV5dkYfXo9j2e7wu2e/VcM7G5MshcFFnZUYpjHmyk0Dwp0Aiy
cnB7jWZ4mMDHgTL3JtUVy875heWe6K1HbvDbedtfP0zwohhD0ddqr7cvltywhR3r8B3bDKeHblq2
1ncgtBPikFgmSIdHXtq9W4vj54UyAj3mMytJCFU2Hqs7mAKRBGWQK84PcgVluZjbgHxOtMPZlnfs
/qoJCcVd4xdLv2TabkyRoJd2ApXDBtMNX/R1KO3u2Ho5U+vmWi/IOqz6DDvyDWJDGLEhneC4tOVA
rINOYNeoKInT0mEIAzC6ocYuZl5ftzC32s3MpUnyOLfCLeqr35XA05lIne+dPS8Ue+Hjtx2IZqtl
zLdfieWHM8FUehainK8NFBmAOtRPLhcl3+XaImQk2HKaWbFdhGWMUHvhzZe7S40uUzUum8m6l1IY
9gYWbTHFgcI1vP4InV93Z6lUQXtpz+0M4YmQPB7BOzWhFwMYmErP9N24zcIZ781SLKvuJtpNONwl
cdQefNBsdd1sxSvO78aDaiMXSGyGGZTg7YhuWK3qG34JyzoBi4gUKksc1jth2iQxP5ckuA+6e1j4
+hV0pHmLS3LXyjno3KMDP3qI7jDyENLuRXJzpzjybeHoHx2kmeoBfn0Ml7X1lLdNA86Q8UMU66q7
0e6rM0/eK+DEV7YVCXdqF9FLw9O6J5ugIIYjd/FoDJm5jFiq1uvAzgLPZKpXqs/RMrd10aTEk6Kj
AlCE1aseFI06O7SZfp8GAiV5Ru+0Ff2HzTuJfVBmy7URkHYQ0D/dPFLg6D3fQwAkEfX7nJp9gzUy
zCqaKCnLZbwdvNj0VDQBqYJEyZKAuBhdlkPasBm8Ac7XXzaMaeZUgkg5fxblKgm2ypcSVKmdhJx5
NNjkkrmudEEob8F/rB8EvX1gYeRMzuJ64JrW+x5kP8KfbZTvrSDdZYFyDAOONGGpEQ21uKwefy7u
33BKa6WVC6BpH8vWBSKfTqsdG5io4N2BHeWgZaKLvBIbl80cFTSm85jX9s7z9/vwotFGK4JvOph/
t5+XFuCH/gkiBEYCDi0LgpIbB43fcqD0Gp86XaM7X4PS+rRnjXRgKdLpvL4o1MyfQVF8ccDQcz1k
qxwadpZ6slGUCj4rtGp4qBppQiNv8KLJCdJJ3HaSHmvQzb09zB8rPuGeCqZsK6Zz1LMVKdMVZ9Yf
hMLRN+/OkZmH/lNb6xnJIkSXDYo6PgJCfpgxnFekzvz/a4990SNqG2y5q64H6E0fpSQmXVy089xu
5ndML7QM/CyNiiVzmMQgFMAt/glD9CAC3OF58ziUnxwXkb4mHftrw3eU9Jz39UKhKm1dMKLkQORN
RBxdQroiiDBWIknAvlGPMZddtLdVZqymWjA67EoqGHea/ru/sVvOs65SQJzb3YvDQb5z7vNDg8fc
xnp7egC6ECVruA6DeboefsFdyCvhfci7tTiMQZW6EgiHc1O9xlRhiWKBJRLG0NgpmxyUQcY5tuxh
ef813kqO/yhJyEBZvU0YyPXOFR746vnsE2hLB0HBPBuv54WU3ZzsfD7Y/6iuD+bJvYqo3dEJU3ZA
SO6uouSXWhqHfdgyCrMpjNu0Kz0uoCKzeY1JY+YBzPJk1hf/kIcj6+Fi0rD7GNofCifoHXcPSmTP
ltN+F1zwdnOPAD/y1djeIyPCWXIIDJutBt10PDgzkCMbWES2iU53x+9QQXGb5tPAaytUMA+Fgold
z1HKtmoZ9Pt3QcO58I/LHiI6aWFHJoAtvw82pXeCCiOyi6ZqLY4cJYoiCGyuhmlXUoOFWZloTOnJ
dV6w6TLdoj0qOQ1NHU5bA7R488r0F0jQmtpJHuXvne7wpXrrPdyCI1JVIIVbQyfzH94Gfo22WWVp
WZe4gf9xNgGsxbr9mY+5Zfg39HzesayfTOsPA9hAy5rpjAMFFNluTvh20+t1JzE6o/6z9bMLvh54
CcxnjQSYgobz3Zr5JXvsMepBevDkrUOfV0KMu+ytGUtH+LTgADrf5t17BwTtN947ioeGDJw38iEL
HMU+gqA4ip/3w3LauGmNJPoi2OkkQpI7o2VfMjMnwSzZAfH0Jt7o8ZqKrH8NJq0MIsyOeQll7W8F
zxn/AzOjaBRaBQ/F1SrUN4/sGyvoIRnCAh4N/feRqzLK32oAuFL20olbQnrTa7HWC6wuJ55W5mTr
Aw4wWUrMgwu6B1InI9zjxOBBedvWe/uP+ItRiXLT4Mg9PEmyXAzGXTSZgedj56FlYBv2YqSoIATa
mwRrKtltxSIAKfiwwZUnWyX5/n76NMRQzlzodZNswMwDqvM6o/GKpZLLNQupbHmxlZ56SkheeHte
gb4N964rbYLRqqMxJ7f3WHRcciYaZsoPivEF/9jyLqmfE+yd+CUMlL79vSD0oNhrU2kFEvo1ZtsC
mbP9au4rNzAk9Tan391Qt76MhQchfVUY1G/H2mSb5HLJ/hDzjA3JVpbtpCjGbnGr1UjM1r1lpB3e
Q8gegfAesR/oPtGfu50isYUBAekS/kOEX8LVLpiZk4Tj0toaYa7zgp0RY+yINPp5ScCqSepnAKgu
7oG44s1DGdsH4FA502lQQ6GYqFJ9MhqKE7KODF0HPv6McJdWRT49OfapbuP+g6KXA4aDZDw5oZxN
nOvodxnT8ht2C3vNdcJxZDvrjskg2Xuc9QGJm4IJVp7h0elXbt4mTddNOpH/7VomglRW+LNm0LRQ
hdX1ApDLhJHl97+agiwgOM/NPjhslW+t+XwHf5BeRdBkTBMqa04+WrYSv2hqro+XRgr2pwRVTeM4
WVtujT5kqg+KiREKe2AZ/ZeAvNec81IomUUBcUep0C4YUZ/TZhucNBY7pbr6CwVdUSkM8INIe/oZ
mFK4GswHIHSKTBxzCpjjDvp2WLm8FV20QXGD1UZIYRVXmtKYzQ2lEiV3/2rYfehhPpOiu1wBNq3l
RF4hmuH9q0fqpY7hjZ7CC9+ygPvE35Z+6d7BKQnZ2AOxc7jwZVFxSA0KcZwcOilnOewBsFtzBdmR
3D02zkWsbZmla6YF960YQlxwpLXRVObwgz3mKEOadheuQHh8yB7fUnSSNQaRWSUWzLBjN7A6Je4r
Q4Rd3Oq42KaUwhECXjNpEGUDW5bQLO4gaBOX6aAufOGJyMSnJ0Bm4bBnxLDYWQcs7kb003tACY4z
h4LtEabAptzJS5dmNTZkRYBc1yDYbjWnvUlgyUrJG8MbrHQaZtnZrAuMx/VvRaVfAhArbLtRYUgE
bK0dcrXtsACY16kR6QrCt9gubxxi1fSR8ULu1fUhul5lQN2Wd1qNpVhBUpZT0eEC4XQJoAdgkwFi
a4NWkPTCe2TG97zqnweK3Azr5ETI6tx7xZsu27ffbIT6JzYQoANp1Vs8tMBEYTFim5estQ6S/5MH
2FEMjlgfn3AY3HEJR2wdlNhu6epCGPrB3N2tImDQjtZx6Rv1wJ8UyoRs7CZ8tsSIlqCeIR0jOAaj
ShXV+ZcAUph1X/jTCJMsp4758Aw6RsDLYzhNdAq0F5XzFPVlcSEm9qbdkF4oDtYLmbV+Q5G02SQ3
aCjHNJ3GjAVvQiDjaihJZZfAI9wLqR/3H6d8ZmQiU8ZuvDISciAbZ/GFn58Kfsqx3ZDOWqdhm1N9
/wSskROPLEmGYZ2cz0mzTE4nZwm5qBXSEYGRkONWBe+tJm5CG3zo9Tk6fpQ43yZ2JjorItHBETD/
hCZK81CSg3bNmae9T21owDXtI4s1j6gYFOXLoRuWWhL0DknkSQr3JHZTemwLNAE1EVC+vMLftR5z
CVaK+R3tJRnKWlOhUWv821j+q9q6N1iLS8VHHrKRtRv8tR7wv7tzSKZN6hDhv0vCyIFpuhDUR+w2
+oWtgLSAnfaGtGHlxGYguhqImvzRFiacs1uamxnc0obiKVQ/zvlIwtwUtVy80S52KW7bU7pdDKbY
0ff/2+Z4Lf8pcTCORhW22I2IEqyj4EJgiCsXGgBNoVkQUHDLO7Z/qAkFdVIiDulZUZgiUC99OKnE
9ydrCjLp9n+sGOX+VyvYkK1BwuxDWnYd+FBCj0Q0UhqrCbMRyb4oIBClRUNSnbZAZ0Pnl4zWCZa7
Ve/6ttbmzCQqz+t92XdZ3wLwn3eN+Xlc9DAb0hZUe4x+ahtinbbiRxNYu/LkfH2GEHFQ4O4mlHXZ
7AVyicOzLHPJPIIHGQW0//A90w+Dj207C+1TWrj7Vb2JHeofR6Tk1wFn4ZTNVOnw/0JGAYg0YW2R
cYIXKB+jrAWxLxxiGQm4E8LUFoYh1ybDfeWhswzOfFYEQ3d4sCrBB0s5qm/hJkFJ5K1tR6mRFzM9
UE32/jETBXNgPT7dcfWFcSX/sFVi9MeDaBhciNjZiqyxp3T5bexgWo+Ispbo1h6MOP6cW7hREHwM
xTonFSmbbSkVL3PP2IidhFNPLL0OVel97AxL4FIssAqhJYf7b3bHndutsgRDBRJf7E4m/QgZgNb1
elYVdQ79TsoNQUvgJ+AYb3xtdP5/j9yEHCRbESPN55yUuAk+mTOwa/S5kuuCs239XyVMIEfHunMc
hFyupbnVATAHdAqub8hIh6HF0qk1MdvP14eGKRoOxL+vcl2jo5Hpy9eBkhrnQUfAFfmpo6tSaMXT
qftYshSWvtRp1IMzK/iPbXxsnOCZ6j6D5ugBhPiuoK/EAf+vIrS2uYGL+deEfcjTD6YC3kTyCASd
pRtqElt2PcbxznLVQZB9wbiu2bleWVow81CUKREMQacuowoE1fILg3FqFXN9FVULWAVPECHUpYa+
5HMPouWEJlcwccLoX7D42DHrBmXMDhgY4I/nB74IWQcUE16VFjUA/SopyfN8pRXsuMuJdG89GGmn
rXWVo4G3h6hs62EX9BGFukbN+PXEgg6fjOveAosPJZ9GocbPVa/z4+ohewkDWEckmB3mDSxKRlt6
hSxm896h/xZigxdxgqeDTQraNWIIdKoQMBFga+jxt1dfvfskZhJG4AnOZkyyEgw+RJ4rxVAHoBpY
BZGUTe5zCyDOs+36tJ6I9q8gs2J/pTUEJUUnIXKFuNAmri5/JaCHnNjsdVSGP1cvZkeAa0VBi6xZ
NvzNQlsBcCiblWUwh1W3xb1YNI8wiA7FFjf87GOEfBXMtBOALjqfXtF8iim+X2R7Aq44JQ/e7LMi
K2EejIb3A+uM9Hpm+CTqSmBacS7ArUxhv5E4+Sk325peoWIPdLUHmMAms2DnrZ0aalKRHarf6gih
fDvrcx6OFRMj13vFwRm8zxd15TG3BC0SCf95qkg44rd4QqdXUto+SvZpp5zgOApCGnzHYFVRxl+Q
prgNPZwtxXxvk7quUKY3DPAc9hqy4uWKrdXksrZFwD/sVXie3LKSdp/aXADzPSsAukMOf8A0hGxk
G1y4BWL3WLAzrpgaGlFgr7FxQ3qBJNG7A6nm/JesX6y0ZVdYrxFZnQ3rw60zSSPplGde/nF/3XSO
Sf+ZSnqhupvq/Er6WkgbtxIjvruJgP3ecS9GExlhGAxqElGvrh4rvPsOuYUh+6iNoqIhiFDtGdwD
QlX/KMo5kWohZ5jMsAWxylKkLAZRY0oVmSKRclJIMXYJcDA8PWGAJzG2UtxVCDiAR79MaQRMddg4
cSWfrgdZCeoqOyzoX7GjIKws69ZlD5gQaRTMUBLxySOz+mgpVWUBc8UCXgeP6L5lyYOxws1xZ37I
vZMFMrwz+ZbvgYhuF5bk3ajDUOj6K4ttBcQfDHO70l/UP/RBmkATtvo/q3aUkzRXgJoSql4Nyg8E
qfUZvBAfp7aj34d9jcW+2RfcsUl/CNPFPmX5l7v8UYvirxwJWRBPH07oUydGzAITqp/53zs6nXAu
GZ/QJd9wL5yDjvqG5mGCSSuksoPPo/YCZJJbRNJp7Tvab42PYpjA98Lav0Ykd6oyPqhMbfPzB8cc
z/bUj5aVXhr5N4JHqs8iZbqk7ojzOLi8UaLz0pRCWNq3Qibm+KMWCXwnOkyW8a/gG7nfdZKLqVMQ
DhVB/D13IpokJ27Tc34AJ1hM2qp2pJRp7Yusq5Q5bjcsgtxdx8T3WQkkN8qBda5b4S7LMjD7uBlU
/koWVjojCiqa3xIvJrGmGIF0BLM4fNS6jD6jS3AC8KIzWsZSYnzDcxHW767NefMy9HilN2i3cwjB
IDYGCufaGAYgfI2BV4NmdDOtr8OFtnS6syt4um6KYa6yWUqXtiq2Y6L3tIs/y2/XjtDJxnFdB1Zu
X1FSwnVsW84ONcKhpzRuMpCwn3vk+jCOQcnbSfEIFJ2aL9AqZWlPBS+6x2Ft4Ny3hNBty3zo4at0
i+hOWBypJHDAVfct0jLghO62qLlAA4joQ9/YkiQSzSQRWMZ/Y3bFj+TwxkFMA7WaUMVjWFkCSdV2
nrCAjeh/7fostgu/IHKhxLCeqsWLCveHp1F0V1Oy3iHP74sUQWU0Z5qsSstuPkfU3DW504xUtMwa
JmTWCDsiPH4cpRPxEDjbFle+VNu2axeQXWXuZ0LI6g4fyJ8mYzFv95qbcijl8mI6pa4jg5gNYPf2
TDK6M0DjZV4lZEwBCKcV0NmV+bYIccZ0K+dccM+s32trhBelTCudRXI0O/o7jtNOzDI0yswtdqG4
uwpEvCVobGZviveyNMe3sDXDIYAE8VdblYXbS8Dn3SmHvs+4kAi3sa2epkwzgyGgQaap16gAI6tN
RGkU9Sp2lW/L510Admwi66k+z0usgMMftNNDLae+eSKhR55DMSTNWtQZBr6fu0dsQ2Ckmb6GGdDM
uq2aeZFR8Q1BqTxO/ohEB+DAJ9NEmie9xeiXsEM9Rwt95ds/6C6OYCjeeQS62Gl3P2hmCKpf1H62
ovV5m9/olp7d8KboRZ3r6aAJljU7EI4YaYpZN06rAIOhJuSIjHvkU8pnW1kmcTd7FxAf9rI+8A8T
devr7shLjKZgpGLi61KKuBrWtY2rkjNzfudRSRCobfM6WDdNWSDunkD5k5vmjb8noFv4zMleegGu
8LdOTJvfK54vsMJYlF5fg8oZ5ABC2KAUAUHRkzrGAPGutflpmBodo1FT6XUmX0LhibnsoAvRWTYl
XKGPHDNYL2ZfYMEza1p7B3/wlNfUxvQeJRUA73CBrd/t3RdoZLxwUPDLTu8Ue8Q1w7ua6ddwMow+
depEz0WRHi1SFpUWkze/gsOvJ/bBkGrjTnAg/WlK0LVyltn5Vzb1IX9+rtIpzmy816JANokswU9g
IbgMK3aSrg+8+zyzu7ipPKEEfH3CGblzZGVH6Mdwaerhm7JAGdNozQTIFyV0XeLI5vnoTnDFPxwL
zuOYKVZjq/ag+k6RcOi1b2FMzFrhv4XXNxMyJLxlPn/1QqG1prq4ax2PZmxs8+BwyUhbc39Tsv0p
Pwe4IT3yz11xbYmDTjSbsfzktr1sV96VD7q3B1f2SeqRindT+NdBiQQm8M1aWhMNqG+4PQUNrfxR
4cz8Nx7jqQjVlSQEwmZ5+iT+OHVdTqW2+nPQqt1EcXCjsQTs3vxBfOaGj9S95vNqlyVwm594JnnO
cUwLHAisBOgeTBIgeIg9YNppYY2w6ots4dtXJYBUgylCrjTpUG3jdx3xmLjWV0d96ZGYeYt/bF/b
uoUNQTTjrR/hlvTfl53K7tHvnd/t4lFIK362n72gxu/2bNESiX44+lin/4WKF/fem63u8WqZX3zT
uytRljNyS4GjAqua8er8fFqy0BOuVyrNwVaAjE25dPd1/Qo7BNj5Q11T0D6HmZvCw92R9qkJq6xP
5XxCe1DUtnM9OrPMkmVgmxguuqwTjpPOXb0cfVTsTfhfE6o2L12QhcO30rdRQvQUUN1DWD39j90P
fVasu6WepETU32HCFIm4Jlh7SgwUHT85woFGd7ditMcp5cxaQ1bdZBOmRBa/fwgFzJuUJ4xjw31l
EsbmMqnYw/KEjVJq6a0jjBam0uB3XzCZsxn1j0kqy+dk3FlfuT799I2ymTlg1Kb2XoEKFHYjU3ia
YjncqrsodJJnOWHvRP+PUAiTZbkrNhHnHoLFB3c5gCHilJeP4/Ew0RMn5a6KHj4Gj1Ck3I4XEeqG
19FVJoA+OV0nXCP9jWi73PooXxkrqCGxAY9PiAkWE7meUChYsPf5r2BRCyzUdiHjIk2+yVnbfj/J
aCw9v0c0X9LEUi3+RxWZuZ0+Uchx19XXzhAFXCQbHYPasLTpQAR4LRStseDHDlLo8Y3Cq5xAgjWM
m2tuE2b9COMBHBh40b9NeVI2XGt4i2KAcyay/BsxO4uchTmbfaJgaSOSQhwlGe/ZcCvgehW3whlX
414/SKxOlDjFRORcyqVSx3q06oOxM26DmbhYqwBEDg58WLLKDnuhBYnSpp/eAgJPg/IaxrPXTFY7
j0aJoTXM6Tjj4ScUErSfB5K/eGm65Xn9bihpYOdSbbAzk7YR+2CuL3OiuqyBCAnh6uSm72WK88Ku
9sHJHghRAafzwlwLgYzdic/JeOTk6vfc3hvFYQgkL/Gdc1y8ZL6faXTp09UNQGTP7Ca4v2+b5TT5
jMTqc4DjTjL8tMVQ4G7Nh0lsppa+hJqFlRk6fS8tDpwIpcpyu5UCYpV2LMwtMBoUw9FmhpVgb6cv
YKZbgTrdB20d1kXb7n2YdQTL+3uRwUWXPjVRzPAG45Tz87NCne5m+/CQUeLptzDvf2430VXiYevq
xb2z8yafgVm9IipWDtSQ3aIQ2W7eBl3qd2saMJc6KwgqYnwFeJs3HRVWF5LC+31pwP+0NBD6/DrR
nMeHhHWM4SLUjZ+JUhThfF4edTBoqf+zE1WKOjrdlCCjpoUYhQl2aL86gi5RypfisY47xGlgvfF3
Et943bCgrF5CaT9Is4HEz5Kfc++GxpuoFYE1nT6mYR9srL//yGUs54qq20NRtr2Af5uhiXOgkpG3
W275RORA2QgvkAxjj7TqJ+UqKP9O8XyypIhs+jXRraBTdZxlP5dc1CtJOIZrHKEd6y+6bDRfabKc
E/zJU4519YKwL+FAzD1QalpZnTl9nKPhPHCXds9ViUmO75noedvmrMhU6yzEy2RSNdF8BLY2kqsR
Q0jn1MHxKwJUv8utRwH3fricxWymhvF/dc+Us9V1sUzzoWK1OX2VeWEOk6mMdshRF2Jh2CnSd9yW
F6s9N5y2aTa2G2Vq3v6pq7Tcl3xI3PWhghWpBDZrK2cogDmQRTU0pYAErsskvZf5rqLMF6xwl/Hd
jNFQ3hVPEcUvj/or6LWyUK6VGICVq9YqZpUM49LHmxTU9AoXwPsIwap6YeZjDPxfE2lsx+JyJga4
sOAB83G4IGVrGOHY/Sf3PaYfKygOyAY59DL6a/Az2JC0efRJZFFvnRTGCmJqBOJHj11UKWLJp1h7
4QKKg4W8QL40IICUHgEQFJACBWnFBOC4rtB7oG6JR7qKCMxkLU8H1bRZhDU2WVpbZ2UqYziRsiMF
XpAvQJFQfsAxDAKXEnK/9reEARvAOq+6xM83hCJbj2smM1Ur51kMML4D20nlu/biPGnB8kTorAKK
IjCJqFqorrvOyPH/NjIHommMmNpPF4kXVZqmi45JJ0b04HO/PvolbgfS+2UwW/VfR7MSPVGmT0G/
DemDswXHPfTAsXR8eLdIjMTRN0jMABuGrtzs93hdu5Sk7cWiPhz4IIu2802NBzoN1/0IJXv/ft9G
fwLWdtmHZpBXuea5nW3pmICni6Kq0Zk+zMWW2byzizwSdjxYL9DthBnv+vS5CuB97QbVfhGoCqkh
iaau/3XB4rjWySWabGFaqrcGMZqBp9Hy4u2qHZDTvwnW7XPkZcR5jUScSEU1Hwmwr3eDYjo4bs0E
6u+40l+s+SJeh0JTO1lG+xrcOmGcUS5AmwboHkdWLj3MnPSeDKHAzjjOY/D/V/g9W6RcngXDSZ6h
wyId9eiBbDlMs/Ayi1BcOjZGxPdYk3pAlttczwrTe1AYwvzrXdEuDLrh/YRXRumdL9kzfrBgk9HG
labm5XKy9LT5jKLs09JhVWl4GXr2CJwMIOtSpUJ/OUcOx72uic9M8sSmtWoaiifh00rtZUakLOZN
noORQbBTHHwgklxTvdgqqWpNatjbV4yIwkn3eQDzZ+C3pUWC0UvkaAodmBsKa3RB0N+vuN/WNbXg
meioE391OwY5OoSovsbepZugG1i0LWzbpxgVjsjjSB6jkPFwylFgXYkfMPDLFj6ALKe6M5wxls7t
axlbZApMv6/2KUOxBEW48wseiFMLbi/9n2W2tHkSo8p7fIwD+qXCSLpFvc++a0uwMNR9tbYGkZl0
MX0VGL3n1C/qX/XVBXHSiQjpNbSTrsM8JnyWrFFqZJGzCzBRA0e2CwaDtfpYfTQ6GtGBXU0Rw+Of
2qS4i3EHaSmvbx4ZAh+MjJ53iQBtRrryLuFcamuNVeQ64G2wLC7itsjkA8rQSvhR7XMGvdJwkxys
xp5KxqGL3IL/2RILHNzcb/q9txoY9z+Ap2toClShlLUOQoB6q7B4njsLN3BZo0pytjrtIuUOipze
zhl++WVl5ID4uQCU5iQEdZGN8dQLlI30IQgVCzcbMdulhdDhZf77KfpGtvzNqW5h0ohdjuUrcFND
HqAS4+L0zQL1LmK3VpvpJpjfDq9mQ8025k+inaeY58VL2qqeOykrUJbeXrXKwsRzsJ3++9SB1nLK
5n6aCym0rwHj2exJKnWgvgpbv3YP3wOs4FZgMN4aasjLrjOugRw+TgxCFAh/w/N13y7i22gDF30C
c/RYYZVy5wmQAJljzm7WHE/3uBSMDIXDCtdGJxY3jbgHgVy/kO2oLM5Q8oahLPl3GR0MXr7Y8VDj
jRtYbhvUdKfHOL6tKEjS9EU7kbhsSPl/Q/aUE2jyCY5HZYX3JXv3FGfMOfda0knS3xZUhPiNw7BL
Q2gexFRuqDy23es9xuRDx6KAE1rUQIqHhVCYN8/760dgFsSlXzzs+2r5xT25jm165hs1lzsNmHGa
sqtO9ZGSPP8ahfGZ8M6aFcIBfyoGkppSCF+8PaKIUxrqlpMscYHSwxrhOKtohoaiOrpUD/Z2YOxu
6KYhWcYwFJ7uOClgxzA4oKLFE6mkc6HSighoiOeoIfJ1sGiVMhGPwUAIbFdSTL7jRzwnfRwYLYWo
zVuxIlfo/A/JoiEmMyqZoZXZZQeaYRSpHJ7Ns4nyj80qgJ6HuNCdexmdeq2tHD7V4aSphj97TbGE
wazx7FM9ewowT9Krn/EFsoPBeUBTPNU3Wc2vQrTWqZ/44lCGQSN0O2uhBHIC2uvEAOAiLmqyq5G2
R0IRxkW1q30LxOqC2NLmxtbuTChCr31Uzl28lGzJjNuQK/uSonV+YcIlzA6pPu76k6IFxqcd6L0o
OwaR7L3od1TpkumZ9zSa1bzVnu1pOvVJ/1k8//OIY8tDbB+8LUeAZRnzy24KgGC2WFz6vey1vyoh
+4MsrhdabD47iXtwYvM+IHobKW14VAmOsnX/QryAbDx97TE2m9pENTr9VE4GKW/kwWL/K3Tm33RC
alm5bUbh4472BzA6ot/D+kXnhp+fBSC70ROUkoA6M9XXfMZkWbg0aDFEnobh7ijLlbUcQboN1/hM
E5pWPhtj4S/amcwv5R68yeaCa3aQJX91YKYQhFn1Ev765FmdkGf4SfZg8EmsPL05EinvWLqm55fF
7uZMc4+nb5khX3u7RXGAe4KCvDFOPxa9Yva0BiS1lmkrSeVMtY4iKeGhPK9dyv/MoJT70fkl1ygG
F1ODDLFwaKVyDRdl7O4ShshyE6w7MHIUQFAp2ZKj96oAkGPO6OScTJUNISR4ZSyN8hPwD8VH04G8
To8EW7ZzOAlWeIENxVpn00EMuhzBn7LPbbAMA2X/b44UYiH2SiuXMtEJmB6P99375ya57WmMN3zS
vKF1lyq3eIPn+lkeW/GF+YZaA3D3Y96AOifVrQ7ZZU5IucyxLyWt+u5UiTTZr3vvv6azNerlKU8n
Dy4jBCFMTg7I9kSbW0EWk7e7URcB7YdNtRcSW3GxMn4hDaapsmzIdS/7xhx39+sa+12I5lV0w69M
2Lk8gKdV2W/cfHCQKDCyyLOjNY1+y+Q05GvZSlvpcB1rY4/cL544jJ1GGxK3reGSLlLWoFb1y/EX
RE1OaUDJAXlsTUsEoVR5zd/oH2f7y8PklXcGnjHx9vDu96yk8uvqOpRI4nCyIMu7dtE4uVMyv89k
et55LXPu/7kRJrp9xHJPKgHVodphhNhmKOND1XtNXL5kt/bb2qpSB0qaPdbQ5W559sI14tw/TU0V
37hNh7TCC6IJlZOo6FB1kehM3a6wMyogGvCBGZd/R+kdyD0JqEIa5ToZ2NeUMSzj94iZlW85vWbO
jOjSUk24ozEcTiFJAy+hLCn3sagUdKprOXS4sh+hEnrywqL8VRxNaf7jcg+oYpqFBS7RuDcHjnPC
GkGgv8l3Z7kFacp2lLLvPTsDqAIfTjwsR1u8EVS9sQcL8UjRR78tz8mLmkOt8VhW/7jKAAORu63X
OgmJ1YWwCS83VUKNvi0LgPgMW0rvTwzP9Sa6qc6EV1KzqM83xXZcuJmeTXuMqmIyq5zeZR/ndyG3
vRY+49GpYeveiUXfDLm92RcbAiPXCG9kDbLWfm3xd8qu82kQIs0V3GBmdi4gOmilKSTp7M4F2WUs
MPhylAv0G8kJUm7KkjzjR8sQU7CzDaPYZMzQ4hHK1c+dnK7ZhWxaM5OXQgmrUS9sbjZcCgvCM9d+
F+lgHdasMdK9XS5L/zvhmaWL9QVUVIhX2KBEl8etnb7zYMiYI6SL5womsrCyWN0fBWPg5Qco8nYw
l+BETP8rINOtLm+A9ElIuZQQ9cUL+j4INK0uVhwnTJBAyw8lhrCAhrdwaXs/ZHtfjopBF+pK+L3q
cU5p9KgbQksB7VoGQXxWJmCL8vEYZTM5s+bMvcUFaAJVq63Gg2s2r6XHb2SDRKzMU8VWV6LjHcNP
zaVY2cJE5FUqJ0mUOpX6/0HOWsEvThlJ1NGs7mWxIvKI63WqlPFCRmU7x6ghvSv2N7t+f1yICOkZ
mxJaWMVJ/VcMVNWPl1cUvikgZpVO6YfqB3skGBd/GIJ/36oi322IkBSl05V3mTPgNS8S6S9taB1i
FhKHjKDxxec6vcpOJK/q9jtp+jYTQJt3xG8NLm3Gh1chBr3hFXdpP7NFAVRJum4jJfxV9YuHKu6q
jfQaeq6R/Uxddji1J37FnKH6igWr6/warSbVHwSVZsZe6f/5ck/EoomhK5m0/az9tUftlnnzeN61
owxUDYJNozPAAC9l6sd3prE5QO2WliQRm51TJmhVA+KOYtp+Bb8XWjC6Rk5lQhmaIz+oaDmcwMQr
Rt7NdAftAg5vDipwl0g4xqsvcQegoNOEbvJSgVYfyWW/GO/IhsQHnIsAL8oufsMEpAucrnSU0Vpu
gPxRjVyDIK3RVUQkszXDM70V0ehQdIxQRCs22CMpLraco41BXTGotUw03wFhMioPss/sXuPVOFDk
Acrrcq5AWCbU3eM24z9+CY2vqTowOk9axu11DfaxUki79V7TLuTuw/fEEpdKeTy7WJzqMGifvJGd
N4PgpA1MPuq3yZraw1EjpjRK6a17V3dlT75gar2uw/wCjrRwoy74UdO8rTTlESwXemOkgqSxPuMk
Ygprx0rYw71itYBxVJhXs4BphFBPoDYjmsNFIgTM24osntPVZ+Wx6SFVZnsmkX5JYhXRvSeyG5c9
idBgohlr5RpumB1HoVQbcz6xtpd5FyZ7x1v+WX8QTQ/CNndAQvpT9mTViwZa5LIQDjZPqbsUyOpd
DLjVwtFgSQYoOdxjx9hW6MkuhjWZ9XRM/fKF9MC68b/2DZHWw0/IC3VvFUsA6HWaiLq2pbyBDdYJ
tjpNF8qX+47tdoieYB/2UlFfnldsDMJt0xttXN6UKPhmlXbS6S89+I1f0W/gS+rtT2zYkuJ5tDL3
87qfCz7SpBq/tBTYJmPj3PolcfN8Gu+RhAPF24ZrslyYyoCnGh7chgyZKY7eCNUN8wYqpdTLhKx5
ncnQiaT0BBPhfTJiU3BFR3tEUJW+e+q1Eb+eXK39Q/YCK4aHewmVC8NjvpxefaNu5+Lgamf1nK07
imU21jou/zzeVC5e84MoSYhBbEoK9F+FUFXUcq7L7pOoJKob0uQSeXTVLTAWe89Fu20hC30RgCpA
ezpQdPv0cUIp0Ht0QvG3ne2HkgC1lp677wbbFdva0dvzGkfzmQG5jYbfYF96FqLLwdXNwf/IpGls
FuvzLD/qNQpNsR5xKjFw6a31XOQifpkG+ddsYpA4i/307/L8KCDXy0+pll4tFSdKqC50VBfUqO5c
lR63NHk/B8U7qcDAAu4Xgni8b6lYQ5c9+MO5RTWSoncN2GH7XasfqNITSooqkrktX1UfdnvUGPab
6jVwGIUmDouep8Y5PTYEb2SROEkVBYiO+0oe9E8TofwUFoicegrJTxdC5+wLXnAlP6iPSlOzJBlF
81eyKwqJnbnzkVvsPIwkwTrYnUerrAhaZdRReYJaYAQxT7c62C4tUTjaCpA4Q9tdPACoFNqzTq4P
inYEw44VRSqNs1vT9VcGbnBR0FAlLmkFccLHIY7l4r1KEs02zgg/bkbQ6KhvtU8EfQ7cu8ULmiJI
KJOKNFAtzidYxkNIH32EkGlW2EXSzk2aAVtVzc2Y5/9qUBBMAL8tB4GNaN/8TscrNuzHGT4kzxjd
aYQ3kqnU87cwlAzQxx+/N1MzX9j8O2jLXNQEIR+5WcenpOFmpG1FwwaYUY2pWxidj5OqR77+hykm
A4by5GsQhXBj/8RaT7WifxOSvzoqv8Ju10tRUWpmkP2wp0hj72UJZv08tXBvYvMsBwVfXb5keELc
JvfC10xqcipAwr1h7MztyDTDRWX/psJY3HvH21c2xMSq43BfvKUu+jUcIP+Va5clKQflsZ0JgCJ/
EAvQYLapHaAXFMDclEB7euH7OvuYvH4BCs9VFGcpiiCiX+7duE8PHcMcV98vpXWjSxJHat1j1N0b
3foQXObHnyTaelX4IIh2ThcptH7O1j8bjjH/dKZFokmxKp7N7FsbwBPzerxRJnA1Ovg7DbMzGqvM
/7Hpj+k8KKI3uhJOkFahb55Td7dE323UUihThj8DXDRDEsi1KyrR3bIu/RPXKhuCZS7Vo3oonUuh
0rM6thQDOBUZSkMsWvNoGZVgo/hXG+5rLqa7QzgfTu2ZeA/UX/78TPBR+lOuXltTOwuZosrovli7
he+EvPt9/tsF++iKX02uOrYuOpsP9lkaWGZ1Hx5B9RoruruoV3Onx1+lsto3+29nXPCCHbLVKjyR
d/6Ts/5pDaWPBpyrLFE1J+GYsgcEAqnVQVVjCROj1KD5K8FE5e6EszjkVLkndqEZdTc3lVvusdSR
Gtse+bfQfylahnkMpQo4CIKETdpb1mQj84F0ZWS17cNLAvXma9vPxiNbrATgo+/3HDfs69IGD+pT
LoEUoSeSKuBBhhkFKPUJiu1QPQDAyUGm32qiYNaZ19kz7W5mbCO6fnuPE3CIQ0k/CodTDvwXNtFC
pRwzdLbMqnFHgMqaJHVGjKfEpxDCetb1GgAAVDIPyAUUgKaA9xVxCBua+B+JQ6ysv/vapFaDJmB5
ZBdPEU1yFkWpFAH3jnXHATjIbShPWN+VvvC80ettRjtHnSvvUuJVjGdMv1M5dg93w+cxR125bfuA
OKBtacrT4+g9/fgORCZ3q+JB3uKXb+aRvyMuCQGogQXkammsed7B7k/b7PqK7r/IeOJLoYnBjmMd
kTvy7EpqOs0pqGF4/r08pY5GVUCRcjtijr1hZ0KCMrkIJiUQTFQyGw10fpxyRy1Z+9OWIc8LF8hZ
fKzOAzXKKN2i+MdiJ/F0PZrFoBnkHtn3o4a3T5BQY6QKzRUhBdXhNZsCjLZJsoda++4LL6SHObrT
+4CbRDKHqaAChUYDAVN3lFrYLVcSXtl+Me6RdKuv5POsYv8sVRzlnaf5jWaybs+5onklkcsf6R7m
bZdR86JT5Df3c8maU/oQhoLe+Q4pjtjPcHjdJduimdOlKU0D0qqnZ0e/g2nB7SP/9NVJu/w4XhsZ
BoDnWGWyY0p3yP8r40viDkLUmdJUKgsx62KP0xUD9Co9ATS2DfGvfC0YYZ/oQljrYk9F9K50OKUI
r0q5IZ3KbEgPd8IW3dku+nEtmZQkC7pR2GJKS/41dIOjtuPNY8Xt1NO78TYxEd65wi+ECOxDTMm0
HEXsPbIklk2RdVaWZvLG7Kp9KkmrdK8cQFI7YXPnqTHaWbDgb9J8n4oiSsR6uQQ3RvOfEXEsVLf4
KfJrzkB30a2ZXOgfs8SQ9gbZYjFMahVtpxuMLxCXNxaSnjly+pdjRTALiEZN+t0zWmdaMivZjWjH
MsW7+AaXDPf/EVFkuWNeUKEPDtPrzshYb2Zpo4ChByBK/WmTFk7Tc0lzfFc5suJzNnJkQZDaPk5p
VI4sYrLdUe4Sl6fWZFYAoh5YJVnC3zJ43kGDeYruULQHWoDhmsIGxwpIzL7Kyd9uj6OCIg5N2beh
OpgHBEoz3cGt0Fl2MaYEYqWaOAp9mo14gi2Y4PnCnFZj+LkU+KKZnIGK45y1SSNwl52BjYty1LwG
w/jVy4QMDwXYmfEDgyFm+Dq7Fil/eWeHyll6++L/DQr4ZNbn/4H+i8f6MoMiMbUKPZUR9B/HK+ZD
pIdexPf3BuORm3+vqlAjXrbkwEizzxtQ6ntIQs7K2HHM5wECMsBqVuBCUWNsnsXoNd8fq8tNIbBm
68VpL2vj5bN2/vOlDwz+iDTYWDaPV6eGrw4+49drwZSFa5aIU2dcnINZ4zWnoWMXOdGNAH+1g1jM
xWESb05b3Z2gg/zMF0fzIm+rrxYpC0oCeTY8lCwhmmk3Qc6jDyAfu6+F9dTmtCK06ujrs8iaQywz
NNRvlpZmb+6PPSR1QGilSm5Ls6qwnLCc2hk6m2osu18B99HDi4Nui1Er6OLnHNyh0JmUABFe5/Qc
lqH79M6BGia9kIoXiDYwJpvx1Ams7V+qAkF61OM6ikjqIBc+U0SxOuPrSHqRusIBZi2LMFZ6Kf6g
kevxTnM05m2pAFOCZPoPbxpJC5pprRDAU3VzPRmDk/EeWCuXmZysYUnnl/3gTvk3NRq1lvWqItxa
0qKDGl3cZRMy1IOKkMVEryiyO6xW64s7qRb+72QHh4TdPjDJWmUSC++5pp8hky+ttPGs7Oadieh1
PHZJ/DP/slw+GKgN7Tbr//CdzZy+IsY9Q3MX80kqlMARTaYtLqeY38MjzSGvxZCXQOv9v7C5TK9G
XHPwXRTflhKfKhmQZK2nyq8R1H9e1tY2XIezFUiHSFxxBl6isiMkkeLRTXt6mo9zW/Bb7hcgS0cX
sqmVjQyhH3cfnjhQRlZn6TSM13Y2sXQnylebsh9QMNWKsSPfGqPAmsTEV1G/hH9kEK4kxMtDwqb9
oZ3VFKFoZTiIl17O7at0RUAwQi3I9wvDvKCGqP8Z5V/DwRSC4qoZvNnvwPffHZ+dcWlqoXBxPAu2
VhB59GL8lUwFXFklUvJVCFZmif42xXvBONiZbP81M7nDWqLYUYaSTi3JN9cUe5oKxPyxlPyM2vaM
rxzYgu2CSxRN1dzx6K7GbaaSeo6spkO/WkoBENekb2l0rxL7d8FqXtCx3+L512X3ie+d0PDMzNhC
bNxFDZTTakSICKA8xzj81C4hJpd4RaKxcze/mro2NFYferQpGnqi3WX2FOKDyP2cdcbUN4MiMLb7
72HWAs3hzAsYPNJpXdZsE5k96exX4J8xeaJE/jnLuXO6HKj+fkrPDpjVjynbmLA3ep+L+vXFNZvK
GrHJ5wx4hTr5XhnMXtTVI42puZA+bj4qBbnfAQGTkWwRjAp8fAvKrXifZdZFoSEyCV68RaJBGCaE
C01VVYzZYVgmn43glupFc06/cOXxiinb26lCSWzbuqhTaiLl/v6OO5+QR914+N5yyxHhmTyW/Y25
usY312aD/Mo3F+4+mR/bzrL/pnwOyjyvXNj91of6ZbhT3fTvWZR2gtcz8JVVtTlqKSyv5AFScKaR
LajKXI+VEfP6YhUVPJ5CXHcJvL+Ui/vrj2j8uT/85+scRJ/yXq6VvOJEv78//OBlxoj7c5KW/GHQ
2bCNSHNx/UIWzaIoHtconY0oz0q2+6T0nZo3KxTWIS31QjTaOfkPyr78tBEnnpxJ5Pjo7ymQE7Ks
d57mfOeAzx7DTh5wNZh5xb5Zws6c7qifG9XxMQ6BapDL+3zVbfDmAMpnJfP5m9xyMlJ3AG7XZTts
xmTnjSXAZw4xj6KrLltIqdBADcWMI5EWoPq7TEhvRFcRAnt5YFW+RMzeOtM3g42ckmenumIByY0x
QjL10ksm8CErsTURsyxjP387GTWaLIM86P4tww6dlPhDh2LOMBY9H5CiyEtSP7tEDMSrXPiadjkh
y4ZhUs00eNXYIrOnHiYLl82ZS9zh8VUyLn7rY4wkPC9Oeo4PsHXBazHIc00FlZ7CkUB8w71fFzhi
92Z7SYBDo9wfmp5UyuqDGY+P+Qqhdd/l8O3q+oGfx9fSpYo8Hd6Rpe5ufAlk0+nrnvv6umNSqctS
uTSPp0hyO5zrwjkrolLvlnSB+H4mpOFqmKjAXYWhOK78ImkUjaXfS6l28ecA1do66yg/tkmrQJTb
/99wiFu4UcIeBVVXoNKZho8XHMJaM0ELR8auCKLseQpuFhRPgugeCC6R84StvXD2e2bhjluZhOWc
atKe0P0hqQe6kuQK/bSJodHZXQd56jcKVnsXuBNmOC26vKg7PlS8BUJP2d0CfmQG9HlshJZTPUn9
qNBpbKkS8uANzDxir1RfQLHjK8QpKmSSev2bSS/9cFz63xoU2KgIYT3IEeRqWb/YwPT4yuVu6wJP
NDDxeNqWbsTkRtvyk67xKa7rRm1hoV1Flk6aDIzzEn44urmzAXarand1UNnw7IEdp4aCAGqbmpJc
fys8Vum8gYF9fHuKVCliNSrdxkfvPWAluW6uqcZs54kDBy3mwVKUU8oMLFCXvguxlQL5qX+CQilD
qG1lAdzYdazGaO2hSjWozHaE9Cvciy/zJwvO3JYdpk79IfTIzYdYbYo4+szHq74DWSxZ5ubbtjnL
M27PWJngXEWpNSwtoP4kdSB985gGtPBoeiZrPmyVhDVKA/fubXnRKLOyPC0er6IQf/CrzbwUyxlL
QeOdwUb5iLZtyyo+AA37uaXi/sq6DIci5yCAj2tV1ht4HSYgU6cUqwcxuaiIY4pJse5iqy/Er8K9
CDTd8sUcP0LTjDqgrB/CKe62jJKswuxbz8wyXCU75525TQWNmbnqwAS4hByrjfI1A0tMmnSeSI+J
NUJpQjfLXphsyoxg52HHsT9yshdaaQlyynAmhZdeVPjL/8b1+IpTih7ScVUk3yaSMmefc1SLNVko
4xu4v143eLF7V1rN0UY0wsiT71fES0HfQMY57b8pb7y+nDshOoqsw7MM0l4Rl6mzuOuBpa6ANDup
Q+3fE2i3bSaXKlfW3cn5SFV9Zv9Yc8hja1tmjRtnzpoW0lmzws0s82Bxh4m02y5jJDM0jKQus4z4
h6ef2/RVG+vNEYwmWLCaHH7A3yblBcMEj6PQm0gvPF8rt3ifm3LfwO99YoBvFF0uEApAVpubJV4S
JoAjXwIjSAU1jEkSKIItXRChAZhUYE1biZ89ZPp2PvS2DxLlZi4AD9Gq3cMVjhQpKO5uo6iIcwxn
1Y/Viuhr/BiPXqb8/ivW1Zye5enO9vht0b95LsJwgEBLNc/xA7kTwpdcYVV+7fqm1T+Kgk01kth9
6ZqDHOvrinrHOLOCXKFtRsRkIiR0OzO8SsuTblJvydlfdXDTMWUyKafp9f2ZzNqsW+msNqBE2dts
8kfgEhY/DyvV2xcyM0eQBkfQm2tGrTLbZoaH7WjiKN78l13MUMpmMIfOncDUmE8eFO7o9qSTAsvd
PQ0crqDQhk9MQz/CLayUgP/ukLDiLK+joP5PKeFNTviKbXeHx2adqjEmdNnbbVd9A+uVAGLhayut
CtIjhRrHsNvRFIGqJRJVIyRWwyBlGpqYzntB24VZW0UOVMY32No34Q+DxrrGagMB/AFLLAZNTnhH
PlAA6Kg7axYNl06B43eYYNTiHzo73c4SVoT89wIFNVtI6DvS+RVZPIGi6ZY2jogQoXcLEDYlh306
X7HwCVx3q28A9OuRi0BXmaUz5grKQ2pVIg86Qe3/DBiz4/RZtV9+arECVRVhf/3iaebN14pqLfny
wT41xQwj9Kkw+4ZJmUevN18+NHWiUD3LK/NcwI7P+FV4KAGy/gnj++hBB5TmMMQEZQs/Tozp/uqB
vByacGKSv2Kgtkb6RFQ5xyAYgsOAFuLX0ZcBSRC3O4Ifr61ZCagjCO0xszGPFaI+vXxBiS1jh75Y
raX5MWOJ0rX+vTOo+Z3gJq1AWNCgwytXaWRjU+RKYK8BMbtfp5N1UVltD/LedyCKCLtnbQSz+6hM
cr3N1KH8to4DuOFiR5b0T8IowdrxKPga/6KIXOcJy3gr1ypHwWzlQRPwnaHEZ1bFEvQLsfbHuXGs
Opf0v/R97v4q2/IoeG4nEui30AepC/OXAILa9COyPloZ5wQcyvxDojU21PHrDKFaRvJyfqcM5i/j
YLTLlqTJce0gebYiRGEGHb7q68NAahuB7pemQ8shcWFPmelvio55GqvidueqJKU902gs2wxHhYLE
c80bCpzgu4exW3oOX49wCIZ2phPNIbb33fCagUeeHVBUs16XyV9ejZN0aphh5HLJqLQYyAKBT+tj
MUeVYmy0r4R0FvSz7mxciQae80U1wloUAySZdw1N3+BPk0sMDKWujRE1NkdaL5rdnxMK/QdEp0Oh
4a/mgYOmmTXsixHH+1FFXo3OAnFK6zYG/nfxEPMurQDgzwsFTfmCVwcC0fc8yRUzzYJ0C6gUjDTz
gkYRzneH0j/3e+KV/mlhsAhl9U/IrJZKdvvt2aK3iy5/Clq2e3baI4gKQJFwKhPZwcqxJAZwqmz6
01LG+XbvHrH4mWXmYOGI1tKjCtNndVlQI7ZgVefrYqaWWpuUwa48j4z7OhodnOIPAWCRv38+6MtD
vZEsKWppU2Dx9K+wE5qMy3GddwMyTHWn9MVIrCW6aoaWk3HVoJQpQSkevZgxScighRpqGNN4vPqa
+38tXIIsd2fKf6ZTfMtnElXA2G30enlT9QCY3TezMPORlZ4vbDKENfCxlwJ+EEn2WCDSy5OSVJ+o
t0ZX6GvNwpD3voKTd4ZloTzWhMCyQCQ4hwn8ut0M4Zz2uSX9s4rPl6HmK/jlJu244jtxtG71jghD
mi79u7pv5fkhfZG0/snX8FsT3+C2Fs9xnzltyIH+xgqMYcJeiMiRY4RNlZMV9d2u+xMNvjNv7i7c
YA9b3rYG2NMTpGoFr2LYtoeexERDWD5BismPajgO0MOGn0wOga6dK0y68Rl59TsPhnRnlaQM/MP6
XuUKhvn6oCMLvOZjZTpkmsymMpBzZKVHqHjV9/xmfrRGa7h38kUP1KIo37SmzdZzx07qk0MH0l0K
eEuaLjK72u0RRc/rnQ9me7trbgT7+chZNCJL878Z9b19XKlC9A6tu3ljJcvplUj/5hIgoO2Mnemq
liKZpJCJO6imZMLPPLbWmdwftjW2kIbF4x42lA8ASGRLKZVkTE0dvGutADuLVUzerNFiZuUrAg2r
74V2XGbHjxJrMcnrgMk+pqns2V9wadNlxTfPbjSuJgxWQG2WBgA2SxNx2nk+er2N2ID6DMwHQ+bL
4TYWOy+cWx3qiczbwh6J+esQJtSNE7fvc1Any/AN8+LEaypZB6rM3szqi7tx9kebUDnS2zD6AO3J
x2p/TAIo0GaxOjzM4Rs8gRljjuM/dyN5IEYdFtm02aWArwg1rUdsPGrCajk8e9ysAqHSUm05piRu
0PI5Krx8eQkhpAffhiGB8kTUAdpiSov1WqvGour6BWcNJmTFm7x23bVru88d+H2SpY2nrDiCy54J
5TXJyQwdXDpBMQkRpYjpOsBx8WUCLpk4sOYWFOfDzQ+R5piA+CHYrM86hyIjDZFEXXLcwl82F5IA
sF22joSZ+Ra5XDUykOCtCYaI1fFZwuBi1atISxjeIX31BhJMR8EOMhYzQRaWwkHJl+hWfsmHgGPX
cPBfr7Si4yuMGfc8Ac+FkLB6pscmic/GQv4xvMUgx/Gyil/vsf5gjpYKFYefB8YhQ3y7iVJ0M9Gu
1ZaumjswBCYT0BtBfzsE0zeEAKZCBng9LaO9eb9ySb47TmlMb8ixdUGdvkfp8OEgij7hI/mXel1m
m++mcSpKIr9bSg4aX0cP301AKj/nUkDKyzTZ+vmrsWJ3w18HRqW8t0lrX3yK/4bEL3iCQyRs9K4U
KqZxrM9ow6/H36v/16nvhsjjKS0r82oUzs1e+8nypY4ybxtlNq+tiZ/q02Ia4bp+EBLpgk1sqcVA
Ks9vybEbHoQm72wcDSs3MEWMGGa9K2DPcPgVOmgMOI1zyjQ4QqhNB4w42tTzbDUhLdX4VP38bmBN
7lEW/cOQAkJdCPju46RIrz7iN34LcalvKLBphGGviGZeDUKc1SmrueBlVKzc3a6PE/k4uhSwoiTG
vGRLFqmj5vjJ0zo6MTkS0pHRAj5ThnjwoVJL5Vh5B08FknFLgVg/mRPVgGGDndJebWAqgGBSNxH5
9iqqq1K80seyau2iW3cQ5zjn8syGV8OaAdzeTzcXu4WUu7+b09RJYmlfOWnG/K3Q3VULkfybLZRi
n5pluWHBwFZSf7fYx3EC9sYWRehshvTVz8Z6okDN9YXJDK3cPlgERfcC4fac+8kWLUZB0Sv46Yvh
KcAN/NpV5XJffPugp+BacI5vqnydQQu4RhZn3wzo6T01RJ5/zmqqx6FbIhoAbIws2Rr+HGpcQwom
Gjens9dIOWxiZsCSV5tZ+PQODSr1kktxjYZ85YwozMgowGZUOAWMu+AzO7DegraH9aDYV9X2MKL6
QNjCHuWXPKUqgp2DNxY9CvtL8c+cPLfBsOXq6zqE9UwsGrW/qrWUn6YSZkRJTgtLtxiNDTROaGjx
xpR6pc9Zphkmvj+VAfGWduE3rF6M+LVxEGQX8PdauveUYxwLAs1UCdSNDb6H25mcMTlIt+bKDjse
SrkFH26wSaQYDRWTha7EXf/+dUCgQ0htBtobrMaQLBH4KYuMXl/O2Se40aAQIr04ENZwGa5AwxLc
MVCt6OW53RbC6ljhCwBOgHwGvJN2deI+XplQYgsf0ct8/yb+IxHTtbxt+WjOSOyLg2uwi4yZLLCG
0R6q5PMEmMPj79iDnoeQu/ag0rem6aJMuGiwNo9JWES2MENdHzczFLMgRfDFdQtkAJ6r5g77SNsz
XwKl5J5bmOOLvtWb9rSeM/0CBocoM6JI7XkfThNUbRoPMCf5lIEvKbzDfG8vlQJQkxBHgi/k2ozT
Jahf/FYDcQLGlWcYMo0/hqM4mYxOf0d9nIywOGxZon6jgEzn1SvgZtu/3zMgpD2TM7lOXctnAYd2
0hrgdKtJAVrn+TIpX3KW6S73fiYrt8XTZ/O/kJql579p+vnYEjQN1sZxICAo93z+H5CdG6qczqtv
wprRJgeJRWXK/Q2fAU0RPgYXsTxIdXSqkPyMDCa8QHZpzIsN8CdgDP0xZAKf7wbGTsBBg0ZfU6Lr
Bc30n8ipe1Tp+AkTcWaplyx8YUFUlG3olZTUCb9cAqqxiV7aCKVDLhz3LffR6N7jH8AnilNkC/zJ
O2O7FRVp2gMfLODFpEI8bAduldsRbR1YY+4g5ugSrlzL7SJgmWLHFO95iKw64GIZ7nOZ7kaQTU/s
dBOSsK5ZIwZoH5pmH1VNEZgYKNjbR/DqHF3QTbeXs5QnzkdSYHM3I3rDmR8S+FoY51YM2zOnyNVc
ouKuDa/oMn3CFL6ZN06jY0jalsxKdrapUNCYDwMp1wZUH7HD+aKblC0oB1CryVfP/3O2jMP8X7ah
2COkQp5xY8UTGMMTTCq4sHu9FIFSniD6sLK1DOcy+Zs0ia+g+hzHuwVi1132oxzu6MzIlvy/Mob7
Ib6QpvNHBxB0nwisEGg8mUHaUjnr7M9UH0y1ixxqw3537vslkzqQ/g+4BFnkDnTEB1CnNjBk60iB
GpqA9hegXafmCM/MTPhcoSq9UcRXb5NQNKzJUxS8CutYTBcz9H4F+BS1XqiviOyK7lbFDg+4QjLS
m7+2phrrJ1vNXJPPhsfnJJU5eaqa/YU0/Nf3r9pzHDuVtLorM2SyDbizt5doyfOCjMGV9hEVUBdR
k72pT6/M+5t8SEeDof7jqzPDhAfWu/Hm3+Rtg135Sl3/u7GzpL+KdGCM8sBh8Om/QUPRYJN+iAXu
HjENx1tJrLHIe7viEFBWNQ1jhvnjdlvu7YAAGLPqn4jWSad9bH0VhjomH/CkZcZPGvsE/Yd35PpW
/if7+K24GnXhA+shqk0PQDR2rykaI204HtmHyZDmOR+WAiOBNM+IgrkxzcE+bjZ+JKhUQAFWqDb9
sv7Ca8JGqWemvDjyx32/Li1S42aAb5CAG1CoLcnvDgRXWkgHBZMl/rP8VP25WhUfJnQizKAVitLy
2yIRgvALzJuTXlRWhWBW1K25z00gK41gI/M7LEf1oAwnG8AuvesoL9xMFCTsFOaOVuXEP+WO4IUP
IQBI+b7O74d5b/2JosQtaTZl/fCDedqPIVTMUjzCJRRvSRyz0uyHpX9d3SIPXbUhKVljcsWcyTBQ
E4MINZZETJWTTyBcOKy3NWdVqsolYS2IEIHDg4DLEA+1lvjrjhxHEarJ2RuNnVOD3OTVsLM4enNx
6dgBrHBl1Mw1ScgC3ES4wyGe1w0bIkRasIbD77y4WBubFIH3Kv4dj2lAliTovpYhhw9MasktZq0k
Gm6B0/ukTSI++d4S9/SBahN8CGyORCXDIfoaOL+SLj8ou27wnN7ZqdqXkgSRvO/yu+OW75DJmGpo
ywX1sNJ5EwxZ6WycSBW8Thk/rPl+q2+dmAIqr0TgvBtKuNJH4Z1ABZMc/JSjXWtcppCAbIFjqTvu
1/rKLr19VSj4/PKNkG+erS7yQqTh6YzR+CnIBZ8Fysrj3oyVdNfz4rgDhiPvj5G38ELwQ4xTLhIV
3N7w55mybWNZfRtQLjvgFVJCbjQ6enjG4/9Uz1v5u9afRWJVxq/f16iMBlapL9yv1zmwzsdwGA5R
MDCiS9lzmmIx65M0ylqHm/CQqDq27FCJ8wI+KjjraKRnYc5rfqI8C63Rqepy3cRIx6DZx6adiqk6
vYf779yYvDmyusOYHCARIjtX/1Mbw83tf/R2aFbbg787TQ385OT2LSJ6XhzRkXzDDYn+xxyBxR2o
oi3K7rVQuvxy0QpnHs3W7PSe7keW7zGbr/moShQ3eVq+XeXMzzL0I2MKfFdzl30JPZYTrInznDR0
e0/lbPbtnm6y+2YA1hGQZD5S0lo3yEDSWeUO/TBxDZ4i5kYphRkVglMd5ojv3W+6+P44OmbD3fhA
pIwxy021FW+9bKvXsNlsG8281yCTD8+JimGOgyO4Tu2NOIg6e/fKotILVKk8UnQ7A47FAHrwfnTO
UJwVJOpmuXao+ZmlYW6ikHcQoiRQXhPSdz2euvZtJ9q1Z2pA/xjtEsuE4ByB44ksWumjagndqzkn
zBrA46bQR62qlKXlN5F/5QjJbEH9w4OHwuk2EiijRXWoeQJtaSTZitwXZowIkIhK7URURtR0+7se
2++XFv0/TeqfCVJsRnpAP0SmdmylvpvjXTQfgPmhgnKGH0wJGmAgVkaZxDBjjk3U7JdB60S+g4C1
2O5RYoWq2nAe+6XitwlKlELiyPWXMKmVKlh0Ibg0Nvkz0RBfnY5Wc+iophOlwyAevzXS1NUnPtz7
Ctv8Knflu9bZUy8aD4rIH71rSgBW+ddJBUFaZQK3RCm8z8DWnbBFAzDdQdC9s+0Opsi6H9TjrjR3
ELiu6SCwDLarx7IcNSf7tKQezLBS6fVr2dBeZowK3Gw9Dj/mJJdZhxru3N3PKnX4KLux3D9TDASv
Qyu4XtYET35+u2CM0rmyAEG1zaQSgoiXvhh8oM3IiD+Fu5Smm3qDiTqRV5zQXjjFJEKq++5JxNG7
MuhqCxWUb+KKwltgbuBYRruSsjvYrgFFDz3b8ia7h4SPbnIfNDBuxznxlthurOm5xdyo515RE2bV
XtxMOncrOjs0OfyJ/8Mka9cwj4Ef9Qwz6uE8AYzNwzViiNjKPu10MVkwX7wO44U2ipesBAf0uU/Y
bDAIHsTADF+4VUubradQYalTg5DO4+tgNL+tQjdiOOyDGm+8QTA9DevmXgn59cYMTMfglM28b2tf
iIpPeLC0+aOrArZsFNsrKy02Lt1+QJF0RjQPQCtULoAS1SJiQWM3i0wZz0M2p8KpL2uzT0PmbeS7
W6mF6zBoDFU2IJUKgbajRiy/tAcIyKbYaHpSdIKf5yka95GA3Lp/3aMx1oXEOA+VQEsvqeXC1jJV
XNKJSPEJ0r5pfudo53j+aElPkzn0/fALV/9XR7kxOD/sw5nAy9xQZzDPKKM/7zRnttFC29EIhNHT
IB8UCC0IhLqRudFc2NaryfME/ccsiYyH0R8Qz+x8q5+0FvfHIlT7JpnCcZ41f4oSy2l34yd+xqQW
Mn4W4xeN0w2ARGHbqB6tw44v6VmnnY3gIYLINo3acjPl1g+tqT0pxHjSvg+0oYP5l2iZD0uFhXec
SvoqqVLAXkvkjT82OmWc01yPUztNDmGEd4D8OYetHYD5XyhRxEQLrtka3IiwGUrS3/hkrjpRHnDD
8Tk+glsQV98kvpKTmfuUOraUeEiuhZT0SR8fskuzaL6QNAUp6ann89BP9noAPTnk3Ag7CepwZtRW
Fr0KLPH8bLxrKcAYxY9vkPAbwU0bwNjhFfPVkUxsWNVMPgkowEwBctKgcsWLRGfuvH+nRU654NXd
XqC4HCXKkRGJiHR0l+3soCVs1oBza7VnC/2Xf97ULxVpoOSV6Rj+xJQpjyUGYeNyxtDotWxeVyj8
PbAy4L+dwiQF2E+MGwZtPexesRe7+g493W+2/jsPkYwkRptWpTnklGHZe01jh03RjAl8MVLMg2yE
BeRIvUCPtDwk2aYW3UAC4BjV3+bj0cCgUhqgoXYuWQgnJSqiUj+BWsgqniO2QYXLlvZHl+tT9wGY
awXowYe1fnufJ2y3WM3Ttpob1WCUZr9oorH8/ZHafoTSF6yMlceS9E3nCBd2jgGkki05nX9pJorr
sdQ/IL8a4UOCvAK8fktRZ+xzT2ayXKVWBrEsoGJbqVHeH5eVrIzAHIKLEyUtod/oJP0iuBC/MqLj
kdsEzAOQi1wiy1G5ZnqyE7tvV1jhwEumbGOVPEsFOI/V08frWPr6HmkgwpXPvS8g4kH65YhhDtex
Rvmf9QI8uXwJPvlbJSOu7dW+ecXNbkAAuOr3lOQE5b+XDVAyK0aaiAPZEWcf+2hpl/dMwD7qiMIp
MWmAykmKHAkWjvWVp068iWq52ky/xRdPyDXzcgTuwETt8ajp6noFwtWGBPiBvNLZ9IjlrqL3x+/Z
ajHHNr3Ex3BBMrGz7YY/uUzmwjLOzNwSpvyOjuCJ3JNFCjQJ0GoYMXwPiIFBQoSntOeHJ1iKMWzG
MrgMsBx5Wrtwli5FVpgbzcS5LMi35FsgzxuhlATtZn1RTJXuxLIPJoEuNBzuHzpjYE15bIe/p+to
O5mn4088Z4pIPLkF4K4HjxKvrLlhoEgKdUZ7ElOTPlyqm0WdU/yFVDyrcq0Lj2ebFa9Uk7yeS9hF
/lC7SSJf/r3plz8RidAUH+pGWC5o2kdVHaURM+dZ/bzVptEP5FSh7Tppq6P8bapb76hqC5j0c8WO
PXEANHoSXxwRJj8+pZlJm2K7kwkHPTjrtxW20xlmleVEnfWeBt4y1hMDTU1dYrtMFGvhN0gXLTJa
uNOTDCPBluXVNfZCNrfJF4+gONJ5f4wjW3cHusJPdkWDynxxKuU7nxtjPk8w6iwbbWBFb8tc+QrF
T+jkOIVZ5X0zHH0atP2xqSl7uEUpP74gzjV8WglKowscN6E/BuNMPuerGpJgJFo56aIfdINJkHP4
NFBixjsg1a4Hn8kdB29CU32S6ldiRGHqrvcGYis8KPS3rUsPmb0OP4QDpRy4DUe3VoB9cq/UMKp0
d/x6nypLbsjKPB4skkMhCHHwyGI5lglJxNCV9VMHHqqzwwcs6YaGm76LYsBf8qd4UC1FIH9NvUHZ
kecLtMnIUkngMYkiazo4P8R2lQcs6/RmVq1IB4Hq3v+aFUSwReXxx7fKOCqvIzYERJo0959WYRh6
rHWPRjuacg78FjBWdv5r7g0yq8Vp+gHOtHD/3ee8Z9Y05sPXWE5IlrnA8AAF8vI+DxK1wxHNRX9n
F5UDqBSQkJEhZmGv3bnynO2SiK91pj7amVUuOMRjMUGrm0FuMtxvoZNGar6mie1gPybJIPyG/ZLc
9ni35OXCzMkkj3XJ5GWhGsrpe7XO5Qh/xOSnZjE4m/rPcBnovZBxTNcbHQdIHlSCGmJ92Hwftc40
7bT1+SxhX+/Nr6ClG0h+4UKLBfVSwElss7+RcHb2AuV2fKpXS1aMTaH1wRL14jgjuuIChUVwqgXf
v98+YOl+6quIfE7MJZVxQv9r11KQutzQCBnNipp4cZZUujoT9j6UhLyOCjCxhC70nkHMIM18ymDF
ztUjYl6GHk/EpIjhaWlPs7mhZFktYdx1O4DQBBq/8zrbIPNzdRj8DtyCnS/ZIhe8lgROtggbbaDD
uNPEj9CkNqCwU0nSBjPnXAnOFlaqDy+pqv9VaOkrj3g1t8ce+pv0C7+d7yqyhgosdjbfpmWC0ICi
sZK42U+GMcB1sHsZTj2xTDwfvZlTKUZFe/mkjUJQPrP/KVjCk4urePyO8ebRSf1CiveStXnvwAjy
iVPlvf/8ypJ6Z/mgy/r3Bh24nXdiDvwC1mx2TEyRrqbfFbu3zxKhtExjJ0AIwnY+81ZgNr57Aj7a
EScj81YUPnpm1ULf8+ieN4IxFkiYxyPf2n/CMPWIZYzPTs5BOLn9laaStBtFiF44RFoSj3kePH6s
g4b01Me6S9ynLkJbvBMWM1RxU5BE7eQwA9V2b8Sa7RJpWJuOyG91Q3oWcGsYqWN5a/jNcPNx0vjK
dJIIxzyeMdEU+prA+j0J8wBff4v5rMLWKcVkPb38GqpOXhFOu+7fl2nnSwt7EmNpC1nFe+vOetsV
ieNaX8e0e7avkXgpKvP4K2fnIyz/n6JEIdhqcqhs9wDUFHdcn0T+pAVljl7q4p+YRWSp6IqMk4Di
GH7ORIVj6BRS01gh8GChtZ3w3E/dPR4Nc4h/m3DLwvpWi5rCIgL9QIDfyTTriqgqXmJawH5vow4i
v+AnqHUqjgLkP+q9IhkQ5BOJ/iIz7TVZKV+CpKuDsiCI5hVtIcSMQ2zYhl/Tzcvpfj7wwC415Rau
1TrnB0Ix8tR7uQA7Kcj6D3D7ACoWTH+4BsojBI/UtVpr3P/Es43lD9sA5Fwdh6AOS9ljH7IQ9jk6
zR5GbAXctC1kkrVA/at9zMVaWvfAS2VhKHrUnwftpbKXAwZFTcpmuw63NPyXN93V+/6yYk9pVPsz
bDHySlBYCNIJqj5pFjV/4Pl8t36FyZFruIT1Ay/zIsovfHpgSCcwx6G9ybuD2D+IJ8ehcwTgvf0v
5vgEOPY1XYHneTCmkoU/F2vOooTnEqO+fGax6WlFIXN68phECO/glbeyHt1pkZBs4KOuxMwhBsLX
lFyLq4n1wUOAwjrZpWfm3gpZMhMxTqqhmnCojHL/AziSJvTRFgvOB/tPSn94I2HIMjH1z+Wqz7BM
CjZNv/+virISvmPKRqbNzA+Ute7c/jy+wuL8HzP3Oh+YkJQs4bandRO7Cvdz23xqLQ/HtLs1iap6
TBMb4zel+p8eDeYSTfNHAoZvGmddDQYoL3UIb6ZGa0/gVpoArY0aGYVL3OcI/mJXrBHrOggQCwI9
S9JJ6d8EbzFhtOOHV6iVbqZJlDvE6h8w5xeNGte4AkTdnSdgj5Y1MyS1vcsdstSF7cdQ1AApAs8o
4igGlhgZaFCjvWmg1oEIADIjE9cjdGYinNGj+dzHPxN+NtWki3+Rkgk/vvCQdeXfhi1bOx4/XgzB
tq0FUXhm5WA3U+ctdzEGjLf1eS88s7LHn4zTKxb+l/EtUxBsNmUkW5cOdnYza/34KiM3voF/TkzI
jCDZxZU00Xt/xSCtvu8DEBDwfMhUATgvirP5MYlzwXJJkdphntDU6nk/WCx5DBUXzKWpBhZ28nWR
oBJgVDAzmTNWW08nTMhEBqUU5q3vB3d2ggqM2hpxO6xmPdbAwpgSE7KgNHGdxhRmli29hQMgsYLA
JTvKmSvsEmK0VCVrSOhz3Wl22iuMeBjkXWM6Al3aukw1LaXFoG+UlKYsHsseDmkxhrIymaDiFubF
+WgtvnPgjCNLB5iFvwvGfOprn8PfbyCWff6Bc6yHqK5xbLcgszUwgu6IuopflF1oc+9Dn3px20Oa
e2kdpWlWHKvK0gEKoSMUFUrTBySjBtDx/MlhznJWo6Fv3QMY0QsZz+T2l+4hevST89iRyyllnApb
8YT/PPKYX007HHiVY+lSApMdWJ1GzDxPFHagcwp6ei/qqlHqGOGPVvvgm6QgU6eFEHvLUA/gX331
IOUTZF/4JNsVJKxYuDpd0TjIMxYSJN7RHnF8hc3qaxX/RcbKG9OWbanh83WgL2A/q31xWhBNHb5l
b7sTGx53I57d4qgzWk88zunuCmSgDGCPe37qwjFsienRk4kAd39453tEtlc1rO7N1mW0cpmn0xAv
DqXn2u0ZUrqouOLa6huWhlJFJDmatBNYBAX5CppuRovhZTEZFU+iy4926GXg1CFudDBhCZfiV7j9
jp+0B6SwMzBrx3qcjpaMmoAaZBCHAiwqV6mpi4fMXJ5mouJYm8WSqIf9hftgdmh+VQNCDx3BXslP
CI/ZQDfrVX5Se3HwZ3/nn3zNXWmVJIjZ9ZM8qSUtbZx03swrPUEmCeX5Vfd7sjA/Yd5ciBOsF/Ge
ILlgm6VXosAI4WW9JSmFYbiHOhs9Z0RaDqun4hZVTeM52xUMvMJxOKAQRUFlRFwitHfT3F4spcqU
W8uy99CyQhRNaxoeWlk87+B5865581OiCrgTxvR4br/WTPbvMCIvjH3SIXFBh8A1oMmWdgrcsUNw
NUvDWxghWheHGpZxXNRokF4rmJDoyvzchwGr8sBunfhM259PVCQyTM/L/SXzV7I4Q/aTPsQgZMdC
8RHcRU+8g271v+387Hd2dd9kFrVX7/fq/UaFxz+RZawCf2i/kfHrnvy8vVE04oBLsrZcvfQMHiyL
JgWYoDzCY8lO/ACRa4Fj1xEdbeRW2X3Or9K443VH4Cug0hkOhUxNKNtS1A8Zxt0slo63tndcP6ij
ekzkPnX44+1IWblRZsU9hYhETfmzK+u4ur9GD5VxA5WBx+lO0y8FLXrmdIy+G+VgZK0znvjMtl/6
lO5YR5mnMnNkCk1hX0o2KSQwLlVNvhLsfXBs+qS6cxoB6YBl0OZfrWP37n+gbV/P5La1cqqJJJlE
pYEx8QCQuwBC2+9FhKwrclTQRXwEDGkPyB8K9KPVib1r0p4Hv6ikzUXdK66v3UJqc7sKJqkjaJtV
rQXujDy/N06LzT+Rj++jHmy8Z0BeS1s+5PkGFkxKycSRsAmoR7I1e1QbdRQeQAi59s7iQDqKnxe8
Woa0myBdbo5dxHiQiL/4E4xWTpqZ4Ss6DZBvsBQoGjQbOD7D1J3DFxdDpfL5ypvIYhco0geOblUn
GgJXwe9Yy04ddQ7RyFC6WZMzCqhLEIKpatmoLMNwuHS+7ALlI0+oC9LtDH+Xr1uUshl9x1aGaIEK
GL7pfQvr2zAkpUdBWaM/wNQsgNXydx/Ayydxb0ONyrSOWcBHotK9TihoLzJA/lsn9gl515B8SL1h
lmvkR/YHMwSre+hEeKsTHF9YLmYlT6mRXqyEP+Ltv0wn7zv/s5/kFDD9vkOziCPoZxxZdpJdIG+f
XRKnvSG2gnnQLPf7wbg277tszzdza1FuOUDge4UY4KsqmKjANAfqHEd5adgMS4Ur/cGDTRm72iPh
TyFk8z0fEE3MNG+k1tAwz7fimpRt/Ym7pc3G+xzY4zhh0/bfVyG+imTvJBaWjoOpJmB44NHRdCYD
Kfvk5uYB0OXMKtClwwKvQ0oPMFneHvFJI2Mw5kuO/yQbnp+NSLFNFgu0EtLwGhDrLSbqv9GwDxe8
10PBgysC1Lzx9XpArAu4sav7HrwJS7N0MD1N/IBEGuxfz1xDGDrYCxzd1sCKYcupL3T02e+f79iV
DDFaYELJHzZ8CKSJlPnFNPnK72ihybpJcxGFk84mQoEy9K9noVtuQshlu7swULEH5cfEY5mJwBAW
oZl02LOmcu+OXurzFoLP47GpwQgzh4aeoXtigH+pG0OqkTDxNsosqgK2hHBnhpjnuX+hWcbtnwtP
eYvxxhj6zFFdKnH5YVNlkGlPx4MeoPujFiMJxto+hyDlhIJfNiLsfuD7NdcK4X/05s7un09XM2wz
2lkGJu70GxrOtfcN/8B7sXo8NWz5TrFCz2yplUGAfYdROBTJSPT2UW3RhAElWJ5EYRmgjrgNephX
GlDHUBTr+DU+mGplYrfV338oKsQ1w4t54MJgGXqTNeMkzQpRH3sKOGU0srq2RBWyn27c2LnN+9vN
dK1ezGBpE3XI/MAB+OwvVGBfnT4tM1wmJtXuSccsxTHROfBIO7Pa5DRvVSKUdOi3Y3huKKXi6Hxi
r2+N/JIWcOJdxKkaawBGYBy3Xa5btXzmttb48rEOLfhvi/XWnOOLD5aCj9pgCHOGW1xiDD2IBhA0
25NpbjnCu4mavH3VGtBl296Wl/TTaZHtU99JzrIjpi33xs4Ti4iRwKATr91j/pche4ga1yYhyoZ5
yGCRi33J65u2jCySl4o5fRCHg+cxxRCxYOOvUkOoTZmOYcUiTfHa7rd+ioq++YfZ9cN7dDu5DhY7
rE2rPq8CxzIiPw2QbKnqrEEBFaJ6ko7Qj7n3fvURc49khJtvXpy0H/N1OODpADPjA+4YWYYugp0X
zLGgnzu8K+6HBj+L4yFdkB/4G2gk6CLbN06CMTU0RT1IxAsLKTlqtrDdn0ibyDhcQeNve9pQLWge
UmVokGRyv707JzCRMywawoOmCQ5ELN2J7pUyVmz/zwH0fFix7NXQL2JN9f2G7qEizBwTW9ojlJo1
F/U/sTKGddbYcwFWlUyEnIIDJqNEy3WWIRC3lNsgj3T8IdjDBZUkBPdfr4TWCFwFFW2jmtR+exdR
EvRva5SZyNLTmLNX/sY6ppaxmtHnUEiTLBIEEqhzi3cFpsby6HPcgW83lXIW3DVoQETZtm69mBWO
E5TZwtblau+oDh84GfIcyiJxVncgvRX9w8uC4D3DNPl7LGdBFq4v/SB6B6QPG7ZICYrljSVHYXgb
DU5I6jy956vrJr8sqT6ZlIxDQmgeK+gplW0Xdaug1i5ie7jzU4SvocqoH8auWOQaPUDiJEvQ+r4y
LwuClnnFWI9qvloeg/u7A4vD9xxz3J7xMNFQNpryI0L1EOcxVlzdXNDsF0bao6KfTeRiw4TQZIzO
ttRMFTwrCN+ZlNHuHdASZzXzspmP3DRBsCPLgpFzXrwYuZ7keL5FuA9evEUoysUJg+Z//GJjjFUx
mGSGYceelWpPOXAwBQOyLMHVr3+h98RHG9GotbNN8z+d7q3vWf5yaBYB8OQbF5xPTfDxtNyCs+w7
K7fgIzT/xmCk3p2pFiLX4bQJJMS62uKVHEDN87vgWNjluSGdt8/V+ZLOn5JUzwhHF1UfGI4CcwUh
vJU4yJwwaGz4kpSNXZ9gkmLBmDLCrBByTp5HGIwsJFI0lZqX1PzBkbd/MgAddIs8CUOZaeZLeJ2/
+K32M/rEBZ5hF1E0qFu2EMivc0ICuFJhYhhaZQA2E0DySe6N+qwMS8xucNGeF6TQqV+Pm3QDTwUC
ES2hrTwFR5Dpw0CFBt4eNYsOfyI+BP+V3VXA5/UCy+4sDUOP6Db/k6ek5nPQfb89cmPhznYQHNYn
K8M6yPt9jq2K/sHHyGC6Bog8ieIelvGyOaCTZCjV74bzpa4VNE3KlxY4HZ1LhesGpYQOCSyoOVgq
FXCj8VZEUnX3bFtwe9keGYYE9blMpyR16/Qif+GZidTAZbEUo4BYdXQjVnyRHjqzwI8jNUWvksGt
P9/XSJGvUZrKvIvBXPYbmHn/MnEouRrkxus8voh0UkeEF6TnDsU1e5crDJc9dch9qOOXcrtl1KI7
ixNxAPaEkIHvQ2QSByCI8HxyCkDQ4QPm2eefB2dU0LWX1nJSsJoheaGzFzEnGa0vz8fwQy6TU8Me
d6Cr2ApUb8iYtCRVu4n9GTrOUzwlsxo0yIZrQkIK4tbMSxMc3WnLSsEV76ETRWQGwk59CM2MRXHU
+i9yTKB3vFbkuyYPvVMBnr3lnD26vfDqaK4aNalyquB5YhLd9p8yCh1+ykF26kq+IOUclBBzCpQ+
u43cQNFSyZ2I8CzAKLDkd5xH0Njyf+0VIXUeByDkL69P0vIqrvj/FCntXwzr+JoulSn3zwDewVmr
g4EiQK+DGfD6yfm3pLdu0Qu9GRiOT++RConulWkFjczXLtTEU1Bt2wlhUewsywo+l4oHi4wtYVSR
6iVQtDkr0OqeM0lZakaJwNkcxe4Mhb7ncIneCp9LuyGe1xoUIm9IKHNfUKaiRBVvgeww640shvxX
Y4CQ8BaS4yl6VMjviJeFR3bTxCYR2bDbRiCmXrLCf9VyKCiIoOwNi/tb79tRhbxPG69/HGIFYHBG
nRt35lUeYzs12QF11EqR+KqcZrSd+nWCjVys5F4P9B7oyaBrcXkRvcov2DzVWiQOZ+kVGbCV/JtZ
fxAe04bzDRqZdQ9n+tYr/R09Qyrr2Pt9d6sJKxjJsVv90TDBd21iCCYdJwdoUQ1uZP2eFQHOywOP
tUncuG3v67KOe6VZ/h7vhHpkuPhtzttpLscP4Zo8hf0rRKEJiFBlsNQhQ8tyxs1ZrHsX6IlvbVe2
I8ws7mXiAgKWj9YE4YHd53k+MAUMmoMFtCEhm6wY2oo19v00U3JdskKx//3726PgFZ0CbeX26819
d5nK1Fo3/0AK1mRo0RK1kfH1UAqV4NAl1qO7/14zJu6kstfItiQBr9TovkpwyKirVlu/WpC73yTo
52pU19CJL9ygT+3X7EIvlQQhko74xmtIWbdUnF62xeEin/qVA+qbvtiDs4Cxt6lnoA45fnEyIFzK
VdhLtybGBlmB6QLgVPMn4pelYm1i235yqgdxmGToneAuZxo5gs6oTyowwsUCfmtHydX/iAy/I/ut
fk5tcfEocJXsHNgMwPg9F0mi2/5Yb7suzEPx+gQLrbu87ERD4UNqzQgk+JTQbZbBDFvP58dO2I2R
+t0HNrFnaRBhzpdlS+NY8O6IDQgY4XiRSBHbGYvl/uGWe3+MEedKVxEB9up212p6OVtTvvB+YIzC
B9/mzrgzRzgngsZzbMXELLbTY+GzPP88SwKdTg0zj26IdAL1dUoQhfIiwGas8h61m8cPO6piaS3V
VNbWCn3MJ0wMZ9cGcyL2beESL/BcqMe8MxTHc8rpfJg4STjFt/nMPBjXW9YdVsNWhYsOEZhkJTjr
436iiN2ZwJvCpMajsS6+/EkQ38sn5hJEy9GqAzqE0oV6FDSRHrXjLSrOAOJjcSg7vWQGCIYsEP2Q
CbZP42hXElCAgb0Bcvg8mxYQ87SeaQb2rVocD368sRrbIP3Lh8phWtXLVcuamkyScCBlodgYHjfO
hj6txfDgM5JMW9xKnVlzpiw/yDB7Xzvsvl9HAZp46jNA58iEdGXpnJT72yp9gQ0T0etzBQHnNDB0
xupQ3QWjwXAgzehmnpaNsn502zO+1BGm2wZN+uNP2MjXz9Q44xI5ocktoOwk+/qSzHJnB1sWhHh3
DD6ZESVUUuXPhjsebHxP96SbrCTP0oqUFBCQYsrsMCh0ZdTGaNML3lyeuiFwMsbnOJkDYH1XeGQd
+B28d/ydnji+b4Yxx8US4ln78gWwp/Vaf+y81mz3H9MkZvKvcMTdnvfS/fJEBDT4YjFVw19kwo9G
H0vMhTghQhIKQhwO8fIhjrhUckXzDPSxUtCf0GZAzryGrsUXm18r8JVFsroHKARLsX6CBzYjY4sZ
fdUIz7+WhGl82vsRG32QFHht2Dsfi4bEqjJlwfCjbG/Lmvm45IL2rWytIPRRpYskwPlP5noJ3YJc
2vqcWEee19J9vrKYWxAc0a6vTDPBZmkr+8r9i2a0evLlt+NycO/ZcSxFWsLza0+l7wMxDMZtSYCw
gjJZZODIrAy0bcUzJXwCYqLeZp083cdzz16JShBYFViiYG8aMeaFzkedia2X3nowHUAY/L0p0odU
rH9DvBBeUteg11E5IMrp/fqrFAf+eC3A5xKdBtej0IeOPE9LlpnR+TkY1pqhowREQBg9Xw9C1Ysj
S45gRwTe/PgUckRpa2FmMhlej3YRpsoWueq/p8VZGODmAQ+qA/6HdcKB8t8Q8cmjo69tiV6K5tet
4jol148h+7mh+FKdpu0qSBJGSNLw/qGWzbgr47OAFgJkqUf4CGZLifVKqwFndrDNYMTZSm0Hatn0
CNvl8bAFX2drByWpkHfVjoNdvtE2VT5+wv/1ErF0ZGb7QUMRH26XXu2hmDx/rbwpq+SniVnTo2sc
c8kPOfMRKwdqZ0FHFRvw/iGzT23JBz4GT/Ay8oDVIYc+SOLUjVyUyznsiEVW/f1/Cj23iHSl0cmU
98blkv4qSjcP+DwXsbf/NX5bgAx/X40Js9uVgD7yz9Is9bHYcdZyD7NHd9M5cJTY+H644O6zfLNZ
OBu0+MkA40ApsGufqd0PNRWTBPJBNIv7bVuo9swDG+T6TQBAw0EM2Y7oneJhkWBaDTnK/ml+sEBp
HivoOB3No4NnzQqVyPOHEUdwMuTN+t00FTogGf5UzwilDPcgcxwYps3xIzdA19PkPZ1352N5gTbg
UI9fSC4d1E5P9yGpn+B0MnbU2ZDvUSlxVZLKL/uDYaxKzd+PalCKBzm/utT1UsgnOB3JBE5f4cYi
Vf5I+dR618m3Y48fe798C53Vp40cf1ShFVub1CgAT9Qf9NiXIWs9T1Ki11qiZjCm6eBbOS9t/3RN
X8QKw9c5q+xlqnqX1tmcn/3ZFF1gA8PSicgVfVZcLmI4fjJ0FqPGYDAI6EN0PWBYL7vBWtazObXA
Hi2+C1VRxL6LfK+XBN+QUFQbv6QBhpj59cKlz8vIRjwnhpzKEbfNPvYYeKLAxLrchXdttubt1eaR
jOsbHYmD593CSz1ETkYV1Sgc3ZYs1yUyb0MHTSYwsYx9bJSch8/xfJk5M0EBoG/k07LCmW1yTxb7
ycHsZ6uTNTKNeoFM3oLCfTrr1J9zNrN/4o4I+BZeIdIccNQoY7t/fN2E1FF959IlexhrjEXQYqj1
Vjs5qIdURCCCPKkEoSNwhsZW+rs/1GdKsiYb16+VNQk7PBMQ5QgLJP/3tmIyN7i6NzA0ZDc+G0LG
6+cFyZ4UJUPxwUihAe1HEBHRxBlahDf4NE4BG9GeMKdjnbiXxp6lkaCHzAAw3l9+Msq3AphKkNRK
2QjfWBYc8FfyHLsza7g/xqIopWj92rtbwknoU+IiKtza3EKXxggFlZQiW+3JaoUniR0obm00oNrL
iYkFcDV31TB6VHzeBwspaN9C8dD9lJHQAomTIgn60W3Q/txs31pLcNX/S6hujDr3kCMnPKZ1P3PI
WcO/xe2IOEL2Vy8dIS5GQprlYYjnRUimD70SlYYoJWRxxs45YA7QObi7WF5BKt3X0mumHJScUB//
BAsEgJEWl+9ocZmQJuZNV+BJbjXZu+qI2S32UYedbqM2w13tDM/0f5/RhiMyxmbxzK/pzNVZY8Oz
XQifZ7rK+N7P6ANwUbWVnw2HG6aMp0TWwdW9SdX2sggjPbsh0ILQg0ktkx1xydFFdVgE2Rh11ry2
uEVzuH+BttPlvRpcky1mFEdI+5U/kw/Pn8J0eEhLO4uFD2FGFDE8ou6LsO3UORhNnMji2Pa+z3c0
5M/3NL4hLgD1SE66OXtwJ7XaEplqT55sa7I9dEFvnYBuD4GsZXjqR+cQXAEc8oy+vBga1/b7wRYp
4b6b8N1h++p77fausy6CXrqwTHsAJblrF0rlkk9qVl62MSK7WF/vfWtIFsu+B+ZkgB89PNmSRKuh
V5T7abR3eKe7v+g1igURDTe5RlN7SjFJM9N1Uim/BjMEP8RQHFcErDCwmqHt+C6QUZZUzwmjLb06
gUt6WovN2umANRarS03eT6QnCYdvROAGg1ima24zXN3IB5tsz0lhmz84bBITw5G00Dg7pTfboMUK
BYzLg7PAv9WY+OXUy+JfKCah0NEUJ58khRNpmcyVZesLy+qD0Mx5MLg0DROvZKrkuypDJQ/OwEZC
67EXCBQuUDteyNit7zzso1lHqSJVo75q4KS1rSpNCpY2YAomFqzvpdM1TZFXYZ3h6lS2tevU9bN0
IRtxWc8nYecjjjuYiDhL77Q1ZPBkh6KAQPyaxIFdC7G8qWXert87QqfXF3p9e4Q7HrF+WRFd56VE
nZaxQ/rOFg3ujV5MLyIjzqZo21VKtGtInEXVLpDyaZRHjXFvdwH6adGAeyeKJZoQ8cSnrXuv50E5
I7yVRz+w4tR40jcmmOqr23HueY31idwWvjHjtDRLqSrBpehcYf753Kjbtd7+MEON13Xop8ETO4rD
xuCM3DorOLa0L/xIw8b0kmdGPit0kbKuIvdVsiLAIN4tYjqze4TUH6NcMs6ljLbmZew9jP2APBFg
FrvrfogUzmnxPoYCXnqdFBfSssshnV9tYNIviZ9WxjZYjUWzBMdM4PCRcfN4uoKqmD8T+p0Jf1WA
IW94MJwWwS5SO3J83N0utRkarwEKA3RUvCf/+qnlqvosFW5TX5N+dWQberFWfG+Zwgn7IdXmEY0H
54bmqwtQz/euy09RbJ8BKTYg+B8PCvB+1q6bDHNgW+WAG2GKa52zd2nBw1waBsod/bWU1hv+cie/
WxOg9AZ43yBDe5bMKyJ3E4HGtika7rrKs0Pox6c/YHsRvHvRvLsaFbUR/lT90qF98sBjwcO84mIC
ZxDXYg76GpgLswihwUvmmKcAdyNfgualrLxcsCm71Gf6vu6921qPyT4dGZKjLsc8X8Ncydb++r3K
hTk9B98rIaCBj13gN339GX/wjLElC/A9f++TP5kRhbKCtYXnYxrl/Yg26G7ib2qlQVDCcNJSF5SX
5VCwvEg3SLbaOr0J72ktf5YYi8wbUr2UIIze1G3Z6Rf+w6eYQvYQw9TSNqE5S0vEx+CV/5XkWUIp
WGGRUQ3+ZFZKqnS7NKRT5xtDqCOnUR9nO/owRzS+yhx2ZDXv0Nq/jzLcc7rJlhTBeemNWQ6oeGjN
WlaqLjsRv4lduzUN5MHcWygf+hYWjh5e3w9noQNhXlTRtjRHFuzJvuRT/fDPA9bdFh7YcOQ7JknB
2qdjG55Xx9XZy098X7mVHnmPKfjVONQGjqNfl3ZzcAAPwROO6UkbO5VyiJrhAMSvU3J/WskUnurO
FdXvLAhlA0qFudmEq2QDcV1EcOinYxtDI+uKi3UARG+2k519RNEC5LsteONLrXPuqzATtNP7PAX+
m1aayXdieGcgJu8DPVaV0dWaofY7vrKcELCMr1/6wh50Z7xk7YelbnUtescsHGZwuI/VvF88kmQC
1FpuDClbyE6YlMr2kQjQhBHVmNyJQqaHGVBdZvTo5jvKGilL+NaCna76Dclthc0mSrr03xWAFxvS
WR+O716ilLwBXaaSzn0+K0mKszf+uuiBnxq93+RK1Eabgrw4wQE0h/rjHA0H4FxeStWH5efeAw2s
u3Yae3PtPSWYGyBlqOYSLwkDmw2Y3I9qvc2SLPnn1YL+zLZQMM87CJo0ZfFv59uQNID6bAjWkaaS
z/mwpH15OPNw8WJk6z6jXnsypBIWMJtNQwYOBJuMNLWn3BpS/jaI51oBNwMH61ClVqaNzBodPXyi
/IK+DIxIBjyIy0wQlRkGFp3HkSeO1Z2bNDQn+ggsCXUXy2IbENkOSpR9y2OesbBPXWvgGeKbOy40
L9IIlQ8V2iPyfdNoPwrAK4vVG7LljK68h+QWjJTTH91dmAf02uhPI8BN840axnuyDJVc2TJwS85K
8Sxu3LUp6TR9Qv19+u+TYVUiWCXyKMSegotf6i6jn2iLe+ckM86qZw6VQ/6VOQHJ4/MC17b5LL+l
kiHJEEdlLBw2jyRaLiRumVmi0Nu3MxdXejx+qzrrgYiLjZk5pOFNIE4Yzq/MMSAEVn/oqojZEaFQ
2hLqQjyF9PnrqMYtkAUHVWQxZmTUI0Pj32bz9e4fmvxI0foBz+YlOgHnz5wt8iYGYtQcPQs97vhR
lQnB/rin4slqtrR/az4i4kn9AJgX6okeWrsXmVVk8bV7BERAocawnZPDpwdqUTRSFMmKPHV6J2dI
POfI09CLJi0HiUoPVy6QvK8Ka5jcHE3gSvkaDfz8RQR3/pYwm3C8N5LJeQ/N1WKPhHiczVzs/Bap
rD+EbUtijO0HWXD6J2mF7ihvwzw8mjVOr4hdyZJpeYi/T123WgAZUOew9Mqo9NlTHtmxnDxPcavm
YI45IzQsLnooXF2g8zX1mZO5PlFeDyUQuET+CLxVWARpp7p87x/1XyTW5+NdE6H85IWNIfhJ16Nl
iFFTVtTNy5q301c6DvGsL8kYBw9z+IeWQJGdENCKov8wmmaS/qPhzGMGeQr2OsViWLKLlOPZ5z7C
d8pdbF9U+BIXviqx6G9WWkoKEbPJZvw3/6LmNj3WbgAH/iHqnfIQsWAiq+RrjU8HJIyv0Hd2ciIa
k/lMqeZLsrvcZ/xNnVLd3nosLJ68ozwsVDtwtS49MWZjbff4Ds0dq0F/vWEOjATPymcpm4MsvTYp
XF6yFvpHx/O4Ifq/AevgphPwQSXwvAtbO9aGuwcRDlHly0sr5Rl+EPwb0vGXMDVGaBf+qNhLR9Np
41GiKZAj15Ju8aeTsX5FSwWrlWvFjSpLLYdQapjkWUq/0RD0Y7RkGe4EZKyXHiHZTkLUwqQq5Uaw
JiVjOAPd3mBk8IgP2YtzIRrtHtWsSIB7cq7JOvZocXtpoizxwZAw4jL7UJahkOlSNZAVmMHLaFrc
/VFZECdv9t2hcXsaXKVn/gWGuhlv3VirRDuofh0xiJ3FTtsc9ie03Gw3D9tzbhVafJz66zeIHRiT
aO8kmNI+KazfzOemaacXv73Pj6EPXni8suhAyMAYnl0tuc6lpiHbvOHRqXq+JhUwD0E/eE4inyA/
q4g5BeAJ9S3x9Qmc+wKEb158Zd2vZsr0F0Tm6Dsw8OWYD+tNJWCIUqT2By1tEXXMavKpdVOXEaeg
cPH1Qnw0ljuA4R+4s9Az3S1eubyP0LfMn41ydVzxrSB2wagxn93+3auxwZ84ccZjVyNiru9256JC
3HrGJN453x2YnLssV1vUXzursdYEgpcGF42azaCVUzCu5vNP0RZ39W+ZG/t91VqwEgBeXjZBp5w+
CB5vFhrpBd0tn79ysm8wR2Y1d55H7mXMQKw6mReXKIsOtFFRlJ9X7lawko3tp51+dK1y9hpxm1xt
g7PHF7sRsXVp8bVN3JxoJEG1bC5YlkPsUZGkVvjPIYT5jkkWv8OBVUh+RA+VcnpHQkXw+JaFpjjT
5KZMh7FyshZh47fEpjykXe3ErVmJe0nLbtGIJgOi67xFrYWAJEBwtVYPpp1+Lv3fydHRF3JVQ4h1
axcsLpiGBKp1aN1ZB429zh3r5EKzLcml5goPfI7LMA9c3prnCKhY1ADKfHSGYQOj0XixNI/ypY4A
AhYdEskevc/0+tK0WmJwIp7Qsf0+16Y10il2OPS9Vti/hUJN2G8YbLp34mBHGXWsXFyJ8+egmOgR
DgsReGame67kX6ThLKGG0l1oxgKBw3Oatkgj7WWRQif9HdYoh8Q3dHSTDYd6HD8ecRpI6mlXONOS
2FztRqngXxrmxeSFKfZFUi12UXlNQYO4J18loVECdz8oT3IXNMT33D8+4Td7n0zUoBwcVGHYuLbt
GI9uPG8mDv22DFrmOBs8wN/WmLJkbp59PAZKhpsOqx2o14hWNaseB0U5txyfs/xgIkQrTb+iGyLJ
YRzPLFqvuz4QU+6nmParP3nPxKML5lQp475xPekBl/R9ExAYMqHTVI6bpvfQEDk6ZMhnO4PIuQLg
xbKp0tKzohi71Z6qD+TmK3ExME9oy6KiwNuZtjbzRK1NjTSCe5UgshDAxSawsVhdMJ1k4bnYqrEn
hGf7oBiotdK0T1lFe1vTDLo6MpxKLpJERtDCNj+Eef6HRBrUF/FmXG1iUoNfiL198eYjLhH8zsW5
W5kBjhwrDe1+laeAjlqVTp+SNSa0Jldz3QSYhik7KpShdUjGyFLYWjux50FdfTy/B5Acrvv/9tfF
65/nocKGqog37AkA1AHv84m5BKA6g3u8vOlL9QmLq1orcUUGSiNJC5pEx/vRdSkgJd5NRYvrLLOg
TLmn9KIkhXjTOU+ZKR51TGbZvWL5XHO4/9/Fgmm+Uznj+RCpaNsst9CX5bvqmzNH76At7cYwrSUV
mw70yidqZYg79uAnZhnTG8iwtOMLluk7Lqv0uQEucDzxP7mK2FG7uCjzO2O6TZ+DzADWNNFGBEjS
ZqygXMiMkkJrSzaiOt7I6Z7JE0nzvUYcHekKfi7/wugT1IUppMhcEWW2QI/O+FObJt15/nSzlmbt
3SlqLVIfpw8FC5NbZmAimgDZ1eYoZ6IVWX7LjSDbGjmByOn/P72fD+QA37er1BPr8+iETcKRDSwN
iWUsGnKFexq4rwF+YGUg/Vsj2b79p5OXexSpnugUaKA+2LFcolyr7jV1lfCGZNFWk21s93IGaiwM
IsTOagCWMhUA43Qxu0u+oPEL3uhlwwQOSi13BElRlJXQYPuw8c6fEe/3KSPVzAS95ZK40hWIVL1q
0yWmr8fpyokb8Apu9zfS+HkDushAOw10g+XDPzRxjS222SOrUyvYM5I8wBzZwFfLdNryT9y6U2uI
3tVM2f0uY/PWh3y8SXZgyEaZ/d/PGFV31f7sPqIHF6ALsPyZmWnEUUzTMLCbLVHHZfAz4wLowC4T
81EU1ivvEHBx8HWRkiffU6+sBseD3AH9q6UmlWp2+JfUaZ2zkpejA+gI5wdI3hE6mHUAxTtx+BS8
AR+bjsmpfoCl0zR7R4X31BoMO+CoF11c7YVnYyi8yru7JrIab4WDYrwADwVw+iKuL2i0ZdNI8JBL
eNqf2/n/GFugy5ndOCQRaK2FNhI3AQ06FgHuCOzYK2fLseC4SIAeImEcktIZkE9XLocBgfF2kf4P
Rkvbr18TpiU3Sb+br3pJ2ik/vGRggj9XoQplzVOcfgXs0BMroLMeo9iIUWU/NmQHsExR3HYzb6OK
MdM7MxSffcCdbkwSsOCJt1OmX0g4yorkVCk4R7jE030fWFH/CXYvWjuNPGfHqQtOL0WnZGdiStCD
NSHl9d7Lj+neKiuCbI/HPInO+ovXalpCM4pj//wA8G/iHwKJiELmOb+Xp2MjLZczJXUxGD/CBSsO
kAO4yLnZU8pQ6fYcgO0QjKv0HeqVZe+2odJLgkT7qGiYadZplQHf2vm2W2WGkGs0XqNDi5JFfmT3
ZL67hcjWvm+OvIvie0cotQGTESfV5amXkgHRsjbQ/Px36aWksmN6iaILwouO3kuZLBjHLCl3l3d0
+yeRUOfNC24SNITm1OO+ILt1WrwFi4vloJbrc4TD+X4f7R1qdiXEEACI5yUNdkPyqCOLwCl4uC/K
0PxUlukC1x5+r4Hb0RPNLQL39Qx7rgdEJ4mNF/6XVKwMfDM2gld/JSQbxlxalOwkHeqjVDhhbGFO
3dORd6xZPXUfgYCiT3RSiVaNk0qtB3FyS44p2IcC/CfqJrKUgi+imtwlw+4W5dTnemlcUKLVOLao
dF9OU2legFLzdYSjxCXT9HZlkeVYreScQYOrQ2MaVOJqN6YkD3rynEmBG4/m+vnnaWjFdCMZMgTB
USuWorTmSQ806UQOPh0sBcqOHbOT8uhW2pWER+oJRRI+TSNHbLJQ7Tenkh+jquJZ2A2LWMBWItXJ
BIv5ZbM+f9oWfQWvaEMWSjPlxXEFf+1v6l81xNo2EePG0qCw4nBmWbbcffNFWgtWMCUFdM0OXdHj
WNm4rUWvNmVI7NsMtMMCxvY1iJnBgs1cQ6x+Lv1T4ACFVUpQkCK0H2STIDnTO7mn6nEmcIrhWHnD
DiAZJsxn/k47iZM+u8qfpQC9lX//UGoZu9hXlSo4vNpw9HPnf6BTMYOhOGsStgNbNWbbMIthlitC
OqVUI2/jTs2l0Nh8gY+7RZrsL5N8/yuqtsx6TVictYFpO6GEuNBZ0dzOQUvl2ku7A/A8RST4c1cl
eYx1JiFe/JCyGcmvn4YOff7cMIK+5kNjDbp9/bdMvzhbYJyWiG3mLNqMGaUgH/cq0StbPbYKS0A+
HLsooS6OxiHUrevdIaygit+f/wHiZl/7IQfJxD84Dl5XNJBeAkFUZOtakjA53wXjobDgI1pK7LUg
2WTIqW4T6n+tIcKJm8sACumWhAG48fqcsBKS6rVqiOywXjbSmHJHpjCU+NuboBDej4s/A/Ty1FrB
WrqWtkfT0siCvRqMi4Fi37lWp5jubs7kni/1ovTuTK6lQfGFXuRUpfmawrM0Tbi+GaI7Y0FlozNJ
s9cj+mm//mih2V/bAoAA1kuAQ4IRS09s8nYXQlKQbDeaHPiYNdrAU7JyuBBvcoc8aqaK9jw3XF3J
biP6SFB4O4PRzHvOEZp6P7CzzBqAqk3RlH9kwAWXfoTTy60g4E6/gTw2vddfCz8v8WI1vYhAB1fn
uWKOoJefQ01Ch5mlohRdmnJy+0TtebYSDufqT2VsRX7w+emrLoLteJKEcPJgOj4PmOEEk98RWbvY
eVgdWClp/0ceNpf+2RPQaGxrlD3evRRByiEvqGVPIETJoIwkxjvgWknd/UKQ5y/Xx5Xa+H3QSxw5
qLVcNkJGhjRj0xd6vDetcHW101QcdshORRiiKGpuAjsTKsd8GWJ08obxFPTW4AO32RKO8j4VGQXH
v/0Kbs0IltUWhBtdNMA0f2VQKe30sK4bjwTLzY/A6oZobBT7EbosLxfoBloLRdmqy52LGw/PFFxl
jmkSwrYuSPbcop0bmvMpq1kiKsSV8c+i/ZcY5d0HQuXxG4wmWIoH7DbkOeHxczIxiNGMGZaMsuPT
fjmEU9iZ4XAtmRCWD7MwjATJA/jPQjcswP9JE3CtewDmzurECQHdIKMx0z1kkim5oOApdjRwF+L+
QjodVExM5xnQZFsAPfjilQpy5/V7CYm8Oh/UZF6YgR7Aamu+j7tL+hEINEcftXqxQ7Nv/MRWDKea
WcM1UJzi3xgkTFZGZmaYtlVLq7fZ5m6wv7lVk4UlXig+Es3tk9sxtiVzq4HDjoJFc/7O4KKs9F7T
sIZzMUPChfjRSm4vaqYOD+EZZp3DVINQxtPcsFYsClaBB9IdhyuyPEuHBrb7hvj4yFKtyuRrpEWe
HOdpxKmQBdHcUycpyhiDEO8Pkf4oX0/PYuVWvr0BNmkglaBTeDH73EutNe6cL5COJQWLmi28EDPA
5RC/rfDu3cxZ0gBZWyJhkzaE2NbXQsJsAjo1oRntuU4sN/HFTDS1dC9ECBr5DIIHa/yuXArX3V8d
y5sDCSMbFxdKjjkkmABpB4+KOiG6bhiLBTeIXhk2KMjF6MCHZfEja2Si6v8K+UC7CB/oiSXdkikm
z+d2qcELznqMp0kFwK6ZmDBauDC2HOanzotCCU/zwCx/sGKg5MFaojZxzJ7cOse24vNgVNi4znIG
lKZEfEw6D22Uk8+UbKWshGLu1dHAkTcDIbiBI1jvfmHzeUV2zvRlYuAWms+1zpVEkcWdDuo12oBW
Yy2lno/cZu+faWQBP2oQD1JXJU6OJUwX7SzdgKvymxH0nWUlGA7qxFl2EGltYwDAAD2iazPAUTRW
RlNbl1vsES3qBEaoliAtvEcO9m++QnQd3vHwHFC6ZvO9Bg0xCU8wWWhPgah5HNBgvcXjK196qxs/
RgHanCxDqcE4QNiigLWqKG8ylEcLrXbRNboihFxCptt8yZQkT4w8ih3HHGORdc6TnY42BegTVYo7
hB+iInmT/JUNpXQpk2L1MqUyM2UAC721fSLVR2Jfy6wlnM7DXQ5QdWfVuGwwIbWgSZhUtG1OPoHq
dFd9DBsaXNDsaK6/yh9pFjWkJ0o3QX1zddk6d8nhKIapWk0FG4ETIDOxdUT4G0tpqEEi58PVchcu
sxPAv7GtYLrPvIw9W1QWnjwv0VdpvLz8GhoukNJ/piB4jTMm65zZYwGnwo/q5O01kwUugelQGI2N
/5UB9exvoGWiwSEnNvfgXDY2HRLZi/KgLMzzU3JBfXLk68W0EZUt8jiEjghsscvZ0qAj1leXaD/+
g5nKy/AooijqyDkmGMzB4YU5mjpRjHJm1jVaeaWi30m3yh4RczJOQ3kxLoeNvlUCU5Be5KszWjtm
Y7mN62k8Agh8qomGyLnCJVpfLGyJl4S7JsgHinv26uCCVceJc8i1Ha7IBRZrEnYjoztGxtnUpJJl
vFP/A9a6tecGYKiZtd6ShwV2S5nuG/dTPUJ93713QwRKMNDTVAGv4P9XvJyf6kWz2jc+gXMdFw/f
BBHwOR9Lym8GBQwcCMK70Mj3XBGF/ldMTtxVxWAUkzH1P1mnEKK+KtstA2emru77TJolyiCGWuKV
f76ACa5gXNwWiy8JHOHqwmqVZvV5ZbhPenVa4nii29jU44BqIQXwGymYd9qtrRfKn+qrTP5+ObkF
4B9XgpYMJitRzocyKTUNwOe4R0EjOojP/zbULN45CjE8kmKs//1FIk4+ELjz9RAgrSz9rBbdq0Jt
cKEMA03rtc0dZKAz5wF8fk9dSu5jV6NijrNjoluohzJ8xTjpaCIbfdKAlEQT8ws9RkJ7ZDXiiYj8
C9I3mHGuYwrPU1U1WXdcCZ5EUWaTn5h39ShG/CxieCZ6SZAmznFo0IBOwcpagq/C7ZLMhxOhKecr
p0tOtxoAd/096HCZgLWDkQcc5WJXbHRkOz5j8d1kQb9Hlb0dg+3FNEmIhJCCGez1VVekz2ueF9JA
MPCmnw8Mc+dDssxz7e0tKBTBktFiU/cY/B/bMky+RORM+IEFmtKp5TPhZuVaBHwAWhAAjPuF+3M4
d+5+Vs8AiTAC5tWk3FNoCqs2sd4TLmIJP5MKDo9v0phWJdaW7I2V4mGrGbfeQIhT0PISJdUZtVnc
W/k4AhHDl6SCh6JtAFMgCTjtKNGbjrd7k2A3zsUC9igKqWOPbcrhuFGMf/u4vWDlhgT/mWihWLR7
sph8tP+PvIIa3YLqqEJWW272cbY2gnsMIVVlMF5cbZRib3hjl0KaAcKI/yHJJiMjnLxY09XYD5y3
iJoVxnq7IIyvpJRu3zreeptbR9U8Nwv/bBJxB3ee01BcqhObatLRxFxXF5Guj5RBjKjhCqrlXNyD
zcn7P0euxxSS4gzxgWL3ljt2VreN7wieu7WxHePHKe5TRxKLQQp7xiyDXoI5C7Tn4s8mttclE3el
X3jzKwYYihYTVZod1sGeJjE3hHtckW7njPRNKgFdvcVHFzgGgjRCtp4aszIAiC0WSc3LOHzkrZYM
Bu6ea+tJjRL9YtJRM9s69NofhAXzQbYrFjF1tKiiN+DajplsAt14xMxd3W3AN4tkOtN5G673HZ4W
q8PNZ1ckWl/VdJ2yjNCjbpFgazGq7jaPv38qnxkT5GdraImdzF9C0ec3AbW3SWuAva7R0gAPvHeL
iPN0sTEETsz1C5ZoZY4dfulCvYSyzaoLI6ESICzdEYpAp+27AgI4G/WH6Fis7xR8T5VzPrLe2ymz
PvghBvDgOp7RgFOIrRYNd7XizdtE5AZqw4WWrzbIOf6DN766kQpZ+I5xpqYSyb1/fYk7m/HF9j1N
BqX/1g3RhjcvoBI7owPL10XY44XN3yftJFC3rg4pJJrzzEu8I8TM+BsAeLXE9sQAsWVSJatuxQcL
YoC+EYkqecSPULCs3UDpj/m11aeDUZEUC6bY1JNaseUOFd02mW3KYk5rE7SUff8BS2wW6SCANoBI
FJWyz1C32bRB+uHqtFxxvPqMSYPvpsn/1nAE1SEH+n+o3DTdJdr68ghSNYdCarK0NkhxeCMaL/B0
Da4m54y6wJm6HWLjDr5gTOtFJO4OwFDwqLTDei+HCzAGDYZxXIy+22haonu/VMk0bM+Kk9RzjRWg
hqcgZQK0ATG5iWNxv3ayp2klViAeglsVg2EXN5SZJHT9KePRUBFKzvlfDLb4wcuTPVsf79YuA2qQ
1qs935+3Q7THLtcIgzQnDZavRQe3SNSBFu92hVzKpuMwztDVtwoSoYm6LWfRKzIEcggkeJBP/K+K
OQRrvyHUFs/e8IfhD+mMsF0OFWzkuc0N4v8mhTardr4YUuPzryDtjEgFIBc4H4A/Bs5QvXXTmQHV
v6UBjK/VUl5UzbSpgihwloeCmgdmjoD+qnDLTqL4QQsz2I34gPj6/BlUDsvKCG/sSQgo92j54+cX
dyFK0sRsuuQebpGKbdTzY5JBdiKU2HRwJPyqtZ11yf1GHWdEB4lmAbi9wglxPZpHJJzsOYU6r04+
FWeDbFWJq5FyWHGn/PG/v84WRdaVZ1tPNixdmDRGbgsxdcjkZKnHIdqBt42TEZTeEzV7zlA1hNPH
6knVehg+T3J5Fy1indUgitXe9ZBuz8EjWMlcejqNPa9tlKfDgU2UNyZr1clm2e4bQgHrtqgLyCmI
nr+08PpYwM5RSphD2SW/J+tpgtib+8aZ2m5f4o9EXdJjqyLmiNtkuQWvGTzkVmU+2CPUV3GOkvg8
YeZqCL1X7m3rcljetsncKStIOQNu47rGt761P+ZJKeEYD/ZZF1Zm+nu6C3rYGY5bIx442eKXARAi
QkSM2xlcwAa3vtwrB+pthI+qrWLLyiKbHqesHdtNPrm7m7Ob5poxgelFCt8Qe0CQLhbN/vw+Ytu3
bLI6HMSP1eu3S6KNMWnQMpVUQfqnHKaq+hSqkjmHJte5Cat3Lv06eMWMZzmZhuyrgrO2wogA5Jjc
3C/ef+MAo/fWAHCqfAPXpw7n/7uWDeGcBL6gmZF2aYe5YD0uDHkbaHgBulA8OkUZBG6r2FmsrEfu
vjmkZ6m06nVfDjLeNGiN4xJ/c+HV9FXm4ed/Cj8A7Gy5ObSMUmaEkihkRjcdgvqYfD3aw3HmCWDD
qatH4iG4NqhgyrP6thXSGI+YAtKbRDkFs5ZCvemctZIHGwMMQrwlPc0BwdCS7rBKsZ5OPUq1fA24
Dj7SQ/XlyIyleWJ3TE1n2fts1VSmAcM9GpidhmNtRHjojiXbHx9HnalS2ncYo52sloa5TKiQERBy
/BZxrExl4VvhpuD+DxJdHH/J3KUO/t1uARNnHgUnhangOBn4qL+DVEiaEUo9LE4PQpBWfJ+JtHxZ
81d4TS4Q2zKDajbYZHd/mknlSF6AfmJNUrjDWF5aIIujwZ0Ql/OUGtP7f9yOZ5hjWQOVlCCANs8N
8eAIYtdMDJc5/+jXYs2076NgxtFjQgoJKltV+5zVlLkkKYZrQtqRCeBDw6Wx0/JbNMb9x+qaE1GS
B5cUU52f602SwlLflyXVxVsQ5GV98jIXTJOTaF3Kh1gjxfmc5l0nxf0s/aJu5ugWe0hnAyvZiw0Y
BZdZWBKQfrI7pzeVlVdUIeHglUJJ/ygFll8d39PyGGyG6yJxWkq8hRh9uOMmqNQh02TZHd6fiN4Q
ZA5svE/VBRZY0dyn49rPDlK2C0s3TExbTf6rUhDE/ik6fNbEG4bJULWdKE4paVCvFnDRrqJZ0zaB
XHF0qrSj+U57Bx19N4lOdRdktw7i0SJb6dnS44xKFFAzH9xcRlId/x/gjIUBBYDeVC/arwBerHOD
K8HUtBPKMRW04ZYgq1z1Bq4OEo+mhnL2YKHKUeAWzF2AXUjpwKEiycbWam4AIe1wsWVVGWQqbwKM
F3WMa9HdxKQycA/6YOgamVpmCnQ098KTqBtj4dmVh18pPtiP6u/YoX2npog9Kr+ONe8mbnDkjaIO
sar31eaag+4ohC6Z3TnKoeiiHCTPxdGyM3HBiMKM3IfTbjeQ7ObsX9tLy99FJrIUCJkafPLM9WeV
2UFJdIG3mxi1qXCFnlAMchf8Mq2Pwfrgp7kbbGcAG9e6GgGELapPEHiCWTHVRcyLljqaNpt3B+GS
nmJ91WlvFGSeVBbE52EHVL92wsPKjq7QfnRnSRt/9DqvtAP7jnW7UcyrAJFSZO0CM42/uYkoMB5c
bsg43+No5A98zQ8mSW4RqYMN19N63AZHl8JxbotZ+72aJmnyebqFpdcGj1kPHerMmRqknrbw6MS/
RBjCcrhmxg3U8nLkHw9Lwgb5oDGPosmhp7MKITGV9VnNw8AsU6W1KlxoDvcFV7tRsWVC+qtrP2xA
jegFns+7vGKPRqazJrl2zMGwx8J8jYzakKmPnR63bdIDcy6Mfj2s2EXBBn1xLupfP2JG9kD/2DQ/
lh9lb58/sZPzvY7dfzOo89YQQBfNvYnO1dzYEDxR698zpkz9GaXaHIy31QHT8N1TafKFhzQdpSvy
0SNKYkz1cqN/JBLubDgHRKn+rUo/K68ZTKS/WWJ8NQdI98KE8/vIGWZzpGApht3kON/YmyMHpXUV
wAbQ5/kLtpKGPfpQowmgJ3exevao9AKdqiayWr+ttFvcKTpUBp7jzL/An7A+hT9pYa1hcZ5tVfwH
738zF/7NezIMYIUgrL7IY5w/4iDqbRs7L2uoQA9Eb5cmDQ6qCfUHkTaAqmOKjgeBOJo5jh3VMRPF
j1AuamQABmkEC76h2QHA2TwkgqT9JjwUSPtjpRImNwOxDjdlStikX701NLyjUsI1VoHEzJL3R88h
ORhtCdAw4ONbKzO0Mss09V7ucbYqXGF2Rv3nFMFL1k1lz9O6Ivg3Cl2T0yEJ9TX54gMXrWTRpiTQ
TlrQiOSvz/pZRUI0Keq3lb1ZA10Wg1LQ9S+whl6s+m9EUKUcd/Zot+1Dh3HZEqsJD1CrMmTxDtL8
eEx6Be8cmWkY4uGLHCAIV7fqIVLJnMI1MLLI2wtd1Nnj3T9+L+Uo8va6DwDsOOaBBUCietJAO4Yl
DiT8oI618AD/D7YqYDrL77BaFSW6+EK2iWzU4HECsAfvKQT/E3w1d/Pq5mQTAdJMhXscUsEuZeez
ttQQajcF6m55F2GDls55ev/u8R8rQUgdKKPdhiaKPPioA4xmTL3opGndezm4N88hQ7JlG6iGscBe
DCJT1WJkmdVhZdzrT631O3j+onp8LVdlsT61eoFedTq8y4b/D9LfSLdHicU4QgbTJOpiMIfQPaNW
71ncFkIvkZqmVCRH5BKJu5GeaH80KJ2II62k3Vvd6GWO8zMql7vO44b2U3EG3fEzEyRclV98mUF6
WJiK9w8rg12ov9bwFVNExYQR1G7kFqe2FjPb9i3nWt/TVFZ1i+ev7ceUhIz0TABC7lgJPjd7pUzz
nvK7WQvhv6DDI1r2LfHoXAhtRInyD1FeV0Z+oARgG+y8QmfYgp/J0anKSP5jqQGHiDJSYydkdQh2
dPRzkqPecZcChJhoDZDAmrYbgLAAgnaDY7xUGbJCanKVNVpQpnMYHOStRf+B/TsHvRwJBCA7sHkM
0o6g70O1xr0Fg5KkgCA+RdnFo++eAwJ3zF+ZJD/vkOIg5rqxWTqZiI/Ib+9WyT0cM+pRBvwljX0Z
biKiX78jck/zAtyymoFTko/bYpvkj8sxcW8bPs3ByDWquLMNKvH22HJCWEv/aahHBrL98E4Y3X4f
VbNgv5s6xANeIzqRVgoL+bSmdTgCP6SpUWqQ0xY4jDWS8irDyUOr4jvJ9bO6GDV+uOOI6zHzEJG7
TIhSOin/bX8Kpqfnhf760kV8ShTqnNxFKYy0KcXc4LD45I+tkNh7BzbXI24xBzVjmbcdY1teChn1
ijmSXzpzinWP7r0UBlO2nuUiTf9NU/qb2U1bXyg7tFk00ubBhfx2xi3RaWZ5ODPezgCuyKx1cYCC
WxIZJLNB+GYKN8Qzts128XjvpcTBEGMTet7azfef7EMOW7/qvlERoYXwOow0hsUXmdS8/9qcZYtV
odlpbKhMp/Tkgf9YfXMzarr7u9dB+LVicLlStNHvHUxdegJ7H6b+0dpopg963ybg2+KSnoRysTs3
cppbhtfLwErY+F31/cOTnvKcU5xg7paw/cLvWij7Qc4v2NcX6qzYz1G06FWtiZyiMWgqB514x16P
9Vh9PZE8OgWDVTd2/rnIyXK4mc1KmBZrUho+JqCJb9pERpdC0hYZ9Zpu+pOe08RYIbdngQoIR12c
TqHxyp5rCkz7kvzySAg3sBdOrUHXVqUdmUtSnebwvby2TzEh4UIsNg0Z+j68KwUluVUC53nC+fsQ
k+jQlty3KEluLFKmgnzcCVdMKIu4vgwI1sdK94QYx6Jz+sTjU6BG7AUAJ7RP2uXxEJ/hd2mj9q/N
tm1qkloRAl2ksdi5cItdISXluA7clDEeHx+hFTAmmbijbIPq489sUFBqTeEnohSRMnckmY57HL+N
sAi9R1g2fjdJP6ce2Y4KhMK+NQ1OVfuOV8joqOYpr4YaL2vQ5SAR3uAljMy6DXipCDJz5sORuYmc
8koX4Et93Ug/k3MLvhP5gk2OdE0Ipq8zsSx3qZTEOHaNsNmX6g2NeYgcZTL/hw1YhSF4aeYyPIDI
nB1z3S0AFxaKgY7Mb3uZAhpyn4QLUEQCuhjnulCWPOx+abkN8NGvsgL7QfRJMsdBKuXCe3DtQVd6
bXa87trgHYTbc8cidBpGnjgGlP7+feJjghh2XmHiVsusdEbkftPVjUiS0bN68U/FpGPZ9ICfoBQg
fCf7jppOtIrZP9bz2XxjeRnO4qXczodiYyBQkMmf7YmxvxFWeEdh1tioQpWIzYc3fwhDfYarhoif
2peUg9RkzI567ykq/TlLShvAjsaN47T6u+upkHoD6dYPSMwjhACRjiMH7G8bCvLXcySiCUgffmf5
XAC9043ASoVn+cyiaHsrCNWeJtMBMDTyySaIPfJpWIYha9LdcO03ixxtu59HfaKsAOKOZHZKFufv
1vrPQEWTex4yK1OM6mqEYhTLnh0kATgQ65otiW35PUOdfib2NXd7ARQG8m6TS/feeffgrxvKvXaA
m5ntfDRM/IT3Y8BsJpesFdtk3ZDGPTk3W/GEFXDkAds4H+EOq2JgdkWChWOmLoRT1DtzGhQQbJOE
LvJKrGslKytmpj8Dm9r8LMck9/gG7Ahj7XEkIYTrVECAV5JagvzghOPP1+WZrjOx7xkjVQkJUWq6
/EmN5NJUsqQ8SbA22LcZeDAI+HmMgPCwppG6VjaotBA01C8N/Sv9NvCjI/geihEsEmciqeHc7tAO
QIZSmreBXb6drVUK83KDpGx2kNS6PGuVh6n0myoI/XlBnGxyDq12sZ9H4TfxzGAQdRNPTTq5+ZlF
0DmI3Z9E/3/80cfCECS/A4+X8GSOCaD4sqhr1N1NXy5jiN1BDC5H1h52ujwte0uH9lZy1a7Iw+Lh
451/Nxh/eAUmgWTgqJR04OphGfKziBIPsYwGOcm7qO2jpWet8RtjUuMnvBQpr65AkhAvbhIR/2fQ
Z+tOnP/0fyFZGNznZJNPgra92wG3V4J3sZ8n/KkQ1Ji4XsFMvhx62Q7K0mS98r386Q5x/5+SVYS8
SF7HeiVjxQhXyoh7Clz0V7eLxBJno0qtNV2HRE1PrxsqSffOCXJF1Gs/AYQSJxQTbCBBh2XKvmf+
Q4LLqP2h7Rn8cFeOwDZ7ODKoooFZLoX4imHRJmZRtBu5+vCYPd/2sOetxFoSs/21Aqh+U2WLm77j
Y84KHnX9VfM9wcpE2k3Z/FfR8QsHLkxAHsewl4gjqkFBH1yR5XAhWamKFcB0VV7ql3j5IpZS+ALT
eDsqOUuKWs1Aq7ulhjWBDHpLUlH6pBgBdk3T7/GCxnBZc3Gn7lQFW07fV6KTpn8p3l/q6pnYR52k
dVjHWqgxwQoV77mkwsBo0ROWOcWdfG4kVFmVXd1XGBomcXVjkLgaEaCVquxvDMZWkeqO2dw2nNdE
SL8AKPIv6Zxl2igfV3yxWGgMEi18RTQrRbu1bBfNm4466qYabJrlXzQ18KCz8cwff/SBfbIgl/qh
p5iuUtimQZmjKgNWT3GovR2alpdpMK21xJ/iEkB5xeS0ggJnzgcVjs2coJF+xJ2B8I6kuYxe/3V9
97AEuv7r+jv8xKIbD8bGOB+D5A/Izj/aIhvWQ0JBgK7DdpXF1vi4HVS+bDOVMC9bSHquvyHpe84I
OwfQMPrGocmO0XniXLwpUOwDC6anKsDgonKxyhV3XEJVGAJTV1t9YXu3uOSvsZklpWpm2/UFp/WR
6ICiPfeRgvktNE14ok6+OnkquhlMkAg8Alf0jBk3YzwVaxVnMC7GfsVEy3l7VsWlkxFZaNX/iUVt
knh3g/5kXEOzmVOuTp1ahbo7HEHDbmpGdk/W36t7MrYxad8e1hbzf7B9vs0Q8GSvvF37gycj+8m8
ZLVk13UqnOaBWZTkGSLRVAwehd4SeBFEbM3Nqn9FOize4qoLRcz0UY7pHNLleXKjsApXLDpJvSzY
x9b2LmYQZ/34jDGy/Xq1BtYnsupJcw+qBw93ppBbrlJo57zORxEYa035SGBqXuD8FX79yR/30Du/
IGja3uBwJVAA88JZhvSAr3TxFZYAioNyWQc/g9qqajcew/Z0Pj4+IQtc3jcQgSyU6Wz0sol0QDfd
HsoBhCOCHw7Htfb16JQ8Jx2B/fLEGOc56zSx4PkvMtsQTxcrbmPfpzci5tRfWc3FV25m0oQiRwBJ
JqJQ9lpUCbOTpOjNR544AFAi4sEhRXz2fVU/JZr7szRRVI7nly2hJF9wz0CI/YIZdfzkOJGKdrfc
NKhqqtuh4tqXfFo+UDIaLBSCo9JgT2186yk84kMf6IkLZiKRskoLTqj+3GSD0R/nZKPrFCLRyrSg
U+OCwr9YC0lFSbOFq3Bg+ptugB/n7kUeVyKSv/Qi2UNeOfzyR+m1A50dMAyHrNekmQKuLZjAcmww
DSQwfwfVArfP7JVTBbiqODYI1anrNfKuGV2yixmhKGdOH+lMIf+MiAosUxRTbwZDcC8UvNmU0D53
nsmUgimxcIj3rbvtBvzv3LMGv4d3UEFovmf/JJ3EDrj50/ccCVkXU9CI3NYEXFyVVh7toKsrcg+J
Der87g5gjuysb2WAWPAi0lPParJyqf3l3kcWvPRWvn5ngX3IlCPF4LYLLjpIk0ntGUcaSS9Tlaso
EOnR1s+VPleIT2PPdobMHenwSibl+5efGCXdmAlYjnbtQgvbt3S8Fs4rTp+gPIklsWyZR0flPXkQ
tEoWuraVga8r8kfOweqxRYVsPQgUMhlPUSsn9F16eW6GHN+1wFoGD4eoO/TuCllSWpdnhfG4WTc+
LsQurRTD8DGAEHtvMX7gxLZd+doVFCfM+2vcTaBp40ES8AKCvWvknqAnThRtxsgOOZbHVu/6UT9j
2o9rtQLnqI62UCBbE0YCQskmkHdcQxixE4tt0FMb+ghrFtZtUJAhdirUMy/Zt5LVGe2qIQcp6ao5
TF5mmj460ed3gHPxlWro6ALpeAaf2UrUSW7nlkFDy5cvMRXMV2CHjHTwwJt8/RpUNuUUJ+CqG5fl
lZOeX+zUhHeGjWhF9b15/6MzIDIqV3sFhtNTu8End8GnYtelY0AY4bM8kVvv6LFgTZUxdBL3DLde
znraQAHTimkdRjxhnKkGvVMP1Ft0UgFevsGLVni7zJYQvytXoDaqFfKTGRgNI9rrlal9MkfGxyhs
qs40uksSQcu9PLeKFRzzH4idh3O1QiPyd1ORNJcysPAinwcMJzRb5riXWKCehg7WNC2KWbufUphD
GAY+i1OyxR8E8y9Bro+PyZjcF3xapf4iQODwlshiuvHe2XPycAZo0BMQYwAK2XdQ7kZ78CX4zBSb
g0H215m9eZFvlCKl/oRW9VLXm3TguD7sLGOcKplh93FJYa+BnGCUWwb9OuGO5gG+OhqEdF9ZBBin
P7RvIu9nOADEF57bgadQXzvzcqTz7Fh7dZHz8HC3m20LL/SCNAPM4tE5KOpVA11Orw2C3bcxGU3Z
FLAXb45dbs+VKLrJh15JUa1KwFyknzoM5Kiq3qISP9yVv+8d5+MJLSP28LgS7hvXZABarD7wT15y
4XMIHmOkTMnqomnvAJN6ovKJjPjcrMWg/VtXzP69WPnfLZpduQyD5rYjciaSrzuFloPs42HiRnfr
7R/a8b3V6Gfy5VpZIq072fvk4iMZEjfo9ffKD6yQS+y0Nx5fDScpERTok54qOnohLI4w8x02ihUp
93daxwkmK8HNoRr3Y55jTOIJ82jy6Tqb9nbqSl6DYFHdtA+gxnKcAfR7//317qoBK47+j93EaLWa
Y82AqNIt+h93U4Y+AAAlwRZD1gyWJBFg5vf3927bPABcRFDtNNExQavje6QBBDVPpB65OGjFRsNY
fuN/f0xxNgHM6dDykDbj0sNVf/2HeAeJcrs8SeCu9wZ2kmW+qlHgYZOJ5+Ogk+OH4x8ywAUUJF1B
U95OPmazI7jS/JWo6PCMmi09mZIkfZbW0TwR2+tG8L1T53O7BtN+MI+nakVkQ6bpNZSVLNkqpLuD
uV02pipigmh4yTm4UVH0wusUO86StnUJBmpUeLdxGM7a0tI0O+eNfYJttaRlU8iSdODm9/0od24V
xgpj1Px+9NFEolXSX+15aiEHmB1nCuEdGnX1vNw+kRHAdhRId16DMTZhKo/nGdh0Xfpv+EEQQzzT
GRQ4tfB4hb+GJ954c/BbCHfvIsnG9V6bw92Ey78Rtfr8XcdC7hSW80ZtZ8JcjvLKjoaDfXyeWk6X
we78lBIqfLiJ/sJ/UHeegEqVAy1DyC270pp/fEgcIxiuL4hQGMURxYlqqpG3/+47fN7fIGSJZZLF
e8VIMIo6PlapKguK1oqPgCFQfAK+NYHGfCjxBAbIMScNfmIwR4YKOMn2r4zxkOqefb5u1BSENzNo
PH8ZqRlBYV9843LvxPmiWnPiu43uI3eDscdiyQd/pNbFlDIUz3nGta8Flyrq+vqAP5yvd1QR2pSa
ECpv8+tu1K2aM1d7fRsEeS79CfVr2FyU3S8JUL3UgTFx6UqAHepxfvZnHepCp1pJlcg+CczTjRkc
U4o73rEQBiIiekany93+XchrhekdnjKD2Wefx0KsBZIZiP9S6gmFiiOmKySTvCGN8AK3LbRlZajL
RQ+CizFThhoWdFTnAWWdL2rVZVI7R+X+liHRan1CE6mopdofn2v0dRi3T2L1yDjl/RPEN9JaAuf8
FrQCr6S9qwlkXuCTPYxiwt2rYsgpb5xAoW9fdO+yjFPJQW2VbVDVM8CKK5TQy2ZcYqfqNDSXVt2V
kG/AwxVRtWqcvPh7SCFCmNrX8IkXnm2UV3g0svTglV44P3fwnacBQh4E36yePeysI5VvRa4JBhHD
3hKP6qM8BD5CFaAU7oKCpo8/jWQJOvkGipv0bS+SbtwDyNtPIT/Ky766kvGyw+9e/l01yJTBWiny
8OJkzcJyAKcV8xgh3f/TEeC9TKrToodmvZaBewMRaNRZ2U0WM3L9DALftXpt2E7gnfYzDNXvkrT+
H0EvWZ+yiL4b0SjtSxNDIxVboORGfAl2QJ+FHCOMIidSuf8FqvJb1JSbYLqMpEhBoRLcn0vK+fHr
Zxa2gdMusqSP98Eof53y+4d0624xfvaXlar/eD6NQ+tlrace0sw89Z75OMJFjYN7KTTZsPJeBRvt
i18s3OAF4WEYWVVTaPN9aXAzbge10PvtyZs2T5zCj3ZVDkEG4PTtU00RBJgKi0xJsg9e18oQ0sTI
A1291hER3fIphgmMjqdceJFSKuswPF1J6cI5yNh4f028UTX8xIp4qwfhqej+Pfvc+lt7kTlcplLw
dFVdJhAccZ0x2eYbJLxXyUrcGmUDfdvetN9IAdpShAj2j9G31woZS5imRBkbWq5bAxWanJDfeLhe
9C/BpqtHgCgoZr9TCBYoY/ze04lZ/lmENUlhPuXx96qoqe8Cv094C+pK8hh4Vc39iDsdxj2psEDi
CKfEDvDsaldu5l1vA+Me29bqSlHNucskdc0tsBvM2tiyTqYjwaHNL6LnLqJJznUk05x/+BXUemSR
8zlx8NshMEZuNS1c5PceFqshnABlROq5fqgcgm2MAxdo4uD5RETjl+kf62D+YKvDpBgLWd3Ia416
qdPPst/yHdKaEzhd+A5LPdgsTlHHdk65qjqBqP2NzqUGjzn0KFFJDpy3R/1PbrZwI+qx6L5elBh8
XsYKq2qWB/W0ILybF6v6Og6KxGEXpto0UmUPZAnQuJJ0cSnYb1OlKhVHBNmTz0v1UmgI8EPJGq9B
+pOVHLfVQrE+p8ZW65Jwremb+ogn0DC833umlGGsaXr59um557jIcPuRy1f/1NBrb20hFv82w7uf
8E7tvbU8cH6dRZFvb+wLu+A2kqE4U4INAyHhFFM1l1W0ZAEyh44+VBBj+I9Jw1G5/WeHA9+l1Zt9
ARfPUVuCzKPLZKRwETWgdUHckAg1Ai4yE99IEgf+1zHF9KOnT0ANn2QeGzZ8mqnmGFoh5kIVXPNb
gwG2mEf6TLHWq/dTDSDXR07i9rMibMlxwMcUkNiOIBLfL9lGEyet6USlRmTy6tUmLPEfoznuSRcm
sJcwoQt5FJq96mX03ZWw8o6PQrv7IBbNsXoPzHKs8OWg6nKJKqoONIRC0l5peOeBT0+PHxiVgA0I
l+7QphtlCiNuKI77XCIQC32d5btAmwwEW8GvFCa0ZGe/88evNctW5hEkCkcMWoheOFaVZr5q8mnN
46cQFGlUFan6i1QEzMg+jIv3qu6z9lJp3xMKZ/GFqOv38TQTpyLPbTsTgd1Xg+iSKWbtzX+2DbZV
LV8NwnUOh3eAFTf0FcAHY+1Zx5h39DD31KBZiMEzzQOlyrTpVxNsdHhO0y4UfFd8xKEryfToHQ6l
sGx7AObyh7Uzb2c66YEBm0rbgS8zaqJXVGI64PSgM6KX2MCcUGtQCr7ZACbbV9ksc95RT3sdChd1
dPAm4XUhJZUiD0+QkIJT+4ISfOD/hT+IKbrWazfyeruyY87yr5JqwZbX9XODYjqWmC7st3bMCyAs
aLcHEvD1eIz9Pse2ayexROq5OBNWdMVnFXcjGq5lU1Vhr6Y+ECIJ5R7n5fnXNjVOu5dw78RufL2P
75v7sNWy2i4vueQzsuaaOSvYO4Mt/62XRxMlrIv2lB7FtiwODRW14Zs5PQQs6JMgvm7fcsol0/c+
Un2tF4ZzuhIx7wRrII7NkgEGk+vK9qOOoS6KcvPjumiOfhUMgXPXTN2nSqNM+QoFfg4mvkai+yXv
v4T29D60EUr+3LzyxeYblhooJ5ZIIqH+Qx1g/kkl5xNZithaBpSZxLQWQm9KVTDpe9GPZMhLZNB1
DAH7Sh9iYPsVqo0hm88pb7HZ64GDnSrXogM4vRXsPdgilsffW/e7Q4kTBcdeOSx1cGBAWPEQ3SDI
ar/oe/jX+9D0/2Pi06In4n2sRPqYQXOZRwaCBXyA6iczs5TxXeKr1ozaKvSoOQvS6nMwFRhdObI+
+tZFhC1GIm2jq2+RRvEfDkevFAk+5SWi8sjqjjCb/YX+Yjk4nKfKqs1s5MhPW7JwWotm/BolIvi8
rcCGz5xqKr6uJAJ9b/ba5lhMPf8+qcNVsm2scJfSV8GIO+oAcBS1X6Hz2UtjqCeC+fd53KGGH83R
iHIvNNATOO0ZPpHt965OUmrZls3Le4HEuYVMIUW0c1oNpLi1yZ9gAeCSoZzAonRkQ5uY/7lOiN04
QuzmGdY6ivmME3Jy4V3Lu6Omc4jLVsokxe5UTq+08ItMe+v6CYKG6pM4fgS5WuogiPH2bg/EwDfx
uJ6kiJgQYZEPJokiacyp8UD4CvYk2RRJONjcuJ3otjyjTeHvNpYJKmqP9Nogf+VJOD6RpSYMN+yn
r6Jl5v0dJmc+VEz4RESGgrvSSuZ48caalZYE25mF5KOcUD8dVaOwR4+qrhLuDiXqIADuvlhm+1Xq
CbhTwLqDhSRLm8VGDN+h/wymkSnGqltB9iLG60JYrxCQhShw80LvmHcrHYsj8ZqgflAkRfoTjDkg
5lLYUDGiPrTwmvT56uIeqCbi+geBYgDuHspX+zXqfry2oBGjJiSZbYuShd5g3sFaPFfpjEZE0gQ5
Kamj6gme709/9Ti+EbTGkgbpAKjbSb8b/82wehv+el3DRLekPXLcHiGgWKNcPd+KGLzg4Ou09Ts+
maz2WntPmFTOEPTU+xrQrn1erbxOalZRrOnVeQwbHM2MFqeYnDib+SZyu9G4zSC6qjzgi/nqjUGW
/crYNrRn6gJ35J7tX22mBa8PTL1ohcaSc6sPqOtjzeI9dSOySKpiM1RS90p707TX/JgSYoI2RF0l
nlMqCv/StgeMiWHV8ETDIjUMe/tV75ak6ADTYeiE26y8VTzOBMOG5XfHy7eS3WFAvTXTkJWepVpG
r+MbsYnRgGE/fZhSNuctpkuY9Ea7dYS7G+C8YfOVpeydDZBbBiUbSAkpHNFJaxNNnIVgBkKVkQxR
dosG8qrQ6iAPiFuUDfehX0mTEXKVtReLnR5zSJq8BZH/5p1gSRyHvGnff9PkSESohjeIlQ2T2a0t
EEb39S5wUjJxVkbTFTz4MqQNRECOh6NXaIRimIcsfedvCcDaCtGVU6aooqSP9lFTjfUfQgc3UIno
XvNoLHbpex/wnNMoHQJCeEXZ9UL2xbhjqw9zzYDJdviFv2TTYHM+9/6V89exhLlzG2hrGcK7kA6A
H7B525FKXqjRUFLx6IvRsKsnbY+kOUF3M15hV0ImXcLfalwJ3UH5fTJvMYWHg3uX1MJYD6CLEI7y
Z7RoSYNpL5ClpY7c5PKnU+4Oe8HB6kuj2bO9/A7D6t8HsISkyamEriqUYz2fp6EgsK6RRALC9GfB
KFQmTGjCTaBRf3q7ML/Ab/87ziereuw5Z3tMSU232ohBlpA6TsepG6gg7BHAKfOUm//4FY6xieMV
a0icra6BrwuBuhhd2i29wl/Z21hFSGISxrJdB8v0tkUOvYdFQ0kPCZJBxfamRfwAUBKvzen1Jm2G
5rT3yfIhXnenZjCxA9DwxfRwh0R7MuZwlghjU1rCpKBloJcpW9J29Qa8ort/CldqHdIzYiDOgdW6
yONBkdKJB0YGmkkC6JNF27xIxYawgkc7LaZPLX6Lv4YCaa9cbkIWU4MwGwUG3lT/T/KVHGZkbW12
IEKQy2wd2wHjYVBockfsfu0SaLOscJsaZ/mox7FvF7SOwaBZjwg+5VZ2Dy9loALSAy3v5fFMJxRy
u5+0dq9eoC0Axss3zhffJs5j3Uwg/grXb06pgHRSdiwqXxZfuWcVc+dxx4+nsK90xL82hruyIpzX
Mg8frg1PfVW1nn4G4Az12EnnOMWkZ1JgKCElqnTz2Ux/lsb+8ZT9QTawjJYKy1tKAmQXueKxdkyw
tRWnVCtHipfob1STrCRY836uQNF7Rx0i1F9WSbco/e3IBAuufOKyA2s1ESR/zt6eGqCURANnXIXe
+3NLyHvQjpOJCC+6MaA/KnmvECHafj579jv1G0R9snTfp5cv6rcANxaQTd9cvHCfwAaLcQx3yl5s
zb+GqKsd7JEXQY7k95cRW9bLsfiQ159K7xoTpm+NyGVym3LoEqKzRhOcYxQ4uK/3ZRIswNgiLFnf
n5MQrKuLBR4GjkmdlJRL12EbJePNDNXY2yNtP6la1+gm4LXLD/dm7rTJCEcvUVF1bkp7td5fYWNm
vYJIkkli5Z+O1rl8EL5WHdd6nDofRls6NOvu15LVqf7EPMixeOIh3wUz8mMz7ZzanuhpsprX4snT
kUMewoW3K7IJTCIzIRa1QrAYhV8pvQcVVpkmkSbcD2t1doiq44WJcaiYcWg0FiPdvh2f3wi/OcIB
+TYQY3th9bWgT8q8FfhHRFeMDFKRyKWLR8Li7qHkjlDhCMdMVY/4zeejq9dEcN8YBQZIj2I3RbT1
OBdk4rd44jv9cvgh3l2JMAX+foO35f2ynd+xr2BudTBc7I3fJDAygz2xhdctJ5cQcwXz8ksUfUCl
K4tFVJW8lyMUrB91wwHqjwVZK11syVZGyNJ0jtuY83Wm/amRZqMb/AXqzGtgXSNuCCg1WOxQBL+m
dg8JzEsH++vYThutClAWTyd4/3p473rIDE3z9LrQSN/SLfEU5v5HpxzpFtssGJJCfvF3+bk5dJ4b
MoFzwc2PtzDKpx49ieka3VuGd9zTYecjoDGz4G3+O3lfsa3GpLO45Fg5W5bZ2xMxfYptlMaJ1im8
MacJonV2uYz/tj1PHK8mRviJEygt4nyJedI+aBiRCP0WrbijC78N7K0y1AMi/xS71zPGCGSdvfNC
dVdqskAyX9t/wmtTvaL3ID/Kkw8n7R511tzKyWsVNi1X9PeeB5zzBzpuM798ol4LRrh4jJ0vWoRD
EKT8omKho1OBYGqtJ+5ejCPEynVlKPXDTWdo51ASK6gJ7qsF1stXFySJCtftJhJcg62wYaXzs81R
3ol1kDAETSR0jl6uX0w2AZGu5RBVc9h8M2g1fB/HAx1DeLmIZ5BvtjFNhNMPYTFPspX0H4OeHdDC
1o57ivwKwMYJC2PazF4tSx+TWl34WkHol5NOe++n8ZrRt8iS2bRd4G5cBx8NWB2dK9QLJ6bj9J40
O1BBBiIKLtvOePQvkSS86slu6eE1eNc566zw2/SigOsZ0t8dY39l4PAt/VugXQ90r2rwHrAmjgMh
ANERitan8heUeJJDvGCD/QD/of0HtEmMeV9s4j4Aisgy8yb75Nee5sCQsH5qvC0qtiLzqucmqzD6
vDqyZhDIbd1GIqa4t+J+Pji70C1F9zWvdrXhqbEOrZf/LUC/hslbkDIasdky6OQNWPbFgfcMeDSm
w9TBecAVVnxdXzZ4OaCEsAnqskVLS5dXkZnOswpSj4dp74YaxZyv2J52Hc6us7F8ZHWm8vdVCaTN
w11uC3vF9WKxfCJlSr++cKtZOrg9a762camKIw4mbH22MfVOh+y0ksjqdUk2WiO5lVtUjq8lWT0H
ZEDpewPTHngv6eqSO6toOqIbIn0YGlqUSkEuaDIGdRSOyGBeL8Vtq2dCQ25+lNgRpvfxbXMlTUMq
mZfqRcfuyZtgH/L0OHhBimirUYPvocYC2kvsD8TR9yfha7ExiZFvI3fDFnALU04SPdDvrkcvVl6R
hEYZuQcZVyEAn/Ua7XI9uhp+MGlW3ouTy/xncrMa/gEsb25WfYuyj0ade5VkJwrw0M0WZY9C34bg
OP8i4XDdXEzaf0eHGqzVyTbmuHFI4FCPMQ1OTmpFcDI7UtBIEKNqhqD4VnUyF0aCwWTyEPV6vtS2
K3a1l2WwkbqG2cD2HbZrfsMu8dX+Qu8NQ6DbNCRBips29zOREnViucQ+tdZAxWxcsPsBGoLmowfK
OMl1geh3cnBWo+7DTIpEkPxY1I8I4rJv/ttDDUwmNdTJh9THe7+/E3M2eb9zy6+jvy+72m+eRkC1
z2p1EUin44yAw9wRIr5VNZ9avLvfw6OAq70xT6awky1j0Zsmho0LJNzLTy+dYsdilmILWubCh3EE
m4hjeCw65eGkqRcGpfwBzFQXwdGUl2beOtEZAK1TcUrKXYjUgRCIyssyJC9+qqZ7sMmNYIS9q4f/
e1KGXmy+aOIJrQ9Y9CDTCIwotCBxU+GSM9hbMGIdNtPE0Rkw4/UiHxzOBSBnh9YdS8KLY1CyHK/V
aaCZq5E8kaA4Bs/lirtIrtfapb8EWULIl5SOfeDrp8tuyVrCpthf9gZDEosD0OJATQ/Ktw0MREOF
udMbWLciGytOkQRuKdJm/5M6eGi5pEDvbrQDzzmNxCV/mvpFD6EwWn0HKQRWom2RfTLD5i7w+31a
P3a2+bd3UWHcNZ1nqrS9hO06h31GEm9CT5M3c14nR56wb9HWpb1e4tQ3rT7k4jQFMW7s6egbVgcH
RQqoIKzO9/7jurNlCvakYiuVVfJkHLtfQ8VzsZJ2aCqr/IsCyCiHxFU5FboMWDm/ShJkgWRxgV/I
y4tRWPKCdf3qBcMFkBVVDZd7e8ChyawabarGiW3NxE0Sllmf1u6D+syJQVTZe/fnfl0AdQ9VrDol
yJ6gxoy+W1ayxSuX6QinXw98GqmE1/7NXLncp4F9bi0xdB67WhGIto6dnqXjYgZsOxh+MTQfw2cG
Uq1ZzsOYRDWS2/gl3dCv8sSkcKAJUs9/FbJIFgJ4JMUUSHgxCnncSgkEtG7ZpMzF/e1QoNsDjdE7
+ToNpHphlcqaIKjuSbzq+LcPw38mocO/2mDur7x3Dq7jbB5q3TXzmd5/sCakT8SdQbnrJpTkMvHj
xvgaajho2GpjKlBjb4T3ChF1jjC5BwlkKl369B+m9uffCIubjVcajOYS7VkcKsq4CF3r6fRG1FuT
Fojanz7YbcHUe1XL9tdao4pSJ6F4mRPuP/be4opcQP5iMF1gqD2s/Th3M798qw2lMapscBAAUv1e
8K8MRSDL/kZC0xGAaC6fN2bTJPYnafmYnGanmcW43SKwW5h3o2+qD2C9hNufCIfK1MDQUPZ4eB3Q
sT8ArIOIoyWP1FCaXhPFOlNALP8I35Xpk1ax7tA4iYyAyTd6KbG7XFiSX5RUUssAqXW+WAm0AJNE
ocVJyldxC4pD2iZdwxUccrOVqHH9QSMu983U+tPW/wPEGKU56nNAhDI/lo823yZNXRexa3oCnHuI
Ybh5URP5+p1J/6HbA4F77G+S8lpjKAXvZBiedGPJDO581fUeipROn/8FgVFuPmwJX1b0mp2MVVJT
GYPEjsqoDclqsQgH0wy0VGUNOv6Fs2YPb8V45s4kCrFATwl+dK5efSlUsf82C7EVvD9AqYpivKxc
XJ/3foVtKzpeKmo2WOW8/pTA48YjUk5rDt/F3IIoEVNd7Xt1dZ/jD1wM6EcC/Stm6yJYqR7xAldV
e75AsZZIelFaM6MBlMWzArswz/Nb5w+oqrOqtjFB7brm7cRuZG/5/KuHdfh4YCgaFP/kbrTF8ALK
H9MtvS62dPvpmGQOjig5QpvdTvJI2YhZHxEUmBuHirHtcjehUGeCk/OsVXc5vMLlC9XBhOttqnYX
7cHu4Iiwuu9MZ2mRV614o6kE5jcAf1pgEdxDUk8qvnD8ZzVvwlVXBVN9AmRHvnQqUXGZvYgvvIqe
wocv1tJpdg4mU5vE4sMB8a3D4/OFSwXuBRWVepBwpqLZgeU4wQhaPyOlEjY/V8DVaAZHP8kW2qAU
5pSV2cgtODeb3vXI6JB7v2YXZplWO2Qh0SooMreVELPXUI4c5rUUDMYt6OC/OfTkYcErNSSJhdSC
Iu810EOoY/67ZHAoOO8CeHqaj5O0ZLOjIHnAsIuB8GW8iuFav3UVF6iji1XNABJKPMPD+YHWdS/V
f7jQ5HD5DwNOFNkmBlUS96Z3T4IVkFDkOd9PQq4HG9rAVNuUwDnN63Q0GMYvxekxdhTATdGQ4LfP
lsJWbdUvc4S1QBJV/VuR419MKw3Hlqd/RpAzmJmksWrLQQfnUVrixUGq0LqF71hnCsfTNNS3wZII
wuAqvHnOQNV+DjG1knmueCHOirONJzv3OCK46vM4eLBI9aXkOlm4g+8yuuklxoKglxgr1ib2JHfT
2a33tze3CAYQkGTfgdkWemknR1CCRpjuT/OQkG6kCOL+FOB82S9Br9Ghek5KSaZIT+XA8kz4fnb4
ipN4Uj0D6Jkp6luPkbOP6nExSmB8CtUIOLLEo3pBR7jIgTNtD8zyCXaDFCcSy/pl/y/vJSjr1qGx
EF3PrmyXK43LYnCoWNc6H3kxTq6e76S1imtUVUqe5R1lcydr530JoyyUdgU52za2YRG2uZI01ARK
YAQUfxU2nB7bVb2irhlK6TsDksOp5OgdPB4PqD2aF8aQtmnnBOsoV7GkPKwsovHbxKAcuHAaXXU2
tE+WgGt1VLw4JqbWnLR0pILEYptVFejVPOtg4dKCV5MoL2EjnNfLINx+sx4/W11uHsQZhM3JXsm3
bO+DAHqW6wxzqBMxh8P2JuhsWOguo+CiMfEj0D3ZLWZWrziu0U3yOfciuhma/9Qc+NzJGzPfIXxo
igLDzZQ6on6cGCqParUP13w7q5Kkuf7I1b96dk+/ZAPKKwknvQgNJdS5NZxJFqd4bAXDmbNl5Kz7
IT80/EiSAGb2oWpw7PbOJblEoA5IEh6Buu9J2tLTVTFA6F2yCXvEgF3waOsTYwFX60imWL8BQ4J9
KuJXHzPFLDx2vsSfAvewIosCTo2jNo7oEpyvTCWlVFwlocHbhxt7pvg0JNjzBCjz8b9+rOzuNv5W
xj/YVj/s7p+Ah+hkxwvwkhKvVm10vZDCG7Lu8FLPIX3q5k4B99NcvqC5VCDXXQbzrO6YJlZMevv5
/bpe9l9zl84V3vKHPbOxzwaOffw7wfIkGxJobfneZYcrB+zegtKmWQS06lQUgeCJ5cpJ6DZpzWiA
whRd97D8s57NERjy9OjmDMce+3NhmuLRV4Gmv0+KapqfxyQN+hktls4C6lgu6lLJuNkOVPqn+D3O
DkpYJ13P3e7IIvltVs3P7A4R2C07+/vu6wi9tWp9zVsxc7jBJzA9J6h1PTXGCduDg4P5UZ+Zxyp4
8KvYo8PUve8MXF0s4nIdiNZyyK9Bxn1UKyacgLqJhLHJbAdinNrC6Db7Jhr/tun3yxIKGCE5g+fT
EwjO0LpxDxqbnpoT40gk1vGONWvv8hWm4WAdoBQUavulRtWQ9mBgMz/kV1ygi9kAvRXlS2pPA95k
TE1JLwBmnRF+W9Zg7Dk00O1WNbJYQY0Vdc6qdS2+KfON0HIWZYcSrG9bKxeUC5e8yTud7Igt5/qW
vdDnS/ahuwH4nqq+v3UcRcvA1CvUr3mfGmwTi+7sWDUREbsfbVOgzUrveQR0dUJhZd4O8kwZlQVD
kViwoWWN6CLDxYvaX8mUL5V2grG7A8KBNFutm3I2d7X8UI8R7GYsspKGajXd4BvOMIX3MPtU0qhs
Y4Im2kfXy6IaWQbBww5L5XyMnDAVdkZb7X498zYz5FCTrC25XKs1vlz3LfcMa8TLnJ/YhDGUe9oM
iS2bsLl64fwts2D++b2sd1Iu9CEqNTPNoPwEbKmYNOVyWRPwoZVZHW2sX9Ahg1jubFY5S1wt/wBH
7SyX+E1QLTtmm8+ZjP13tH+rKF7SrMLKoYsL70k11hiVflppGgdfNFDNtXLf/za/RIeBpCtGmiu3
dP5MnfFllLdFpBbs1rzK04cQtJLBQI+Hr5UMMlMx1s3RpoxC0mbmLBeTDdNj6zopcDMcCJUvAE1W
UNrJyVxYzlnTnYITxf9/RZ5FBWgcQKYfRjwzIiwdN8NGAUzoberBvxzzRm2JbOvnJcT7h/UFomh7
/zG3cpq5/tMyHwhny3F9i8cCeRTtEVnkSTLz+QGXltkUy+yzl40U5Ru5eqqQj2+WTVPBxMIGP3Xs
jJNkdRt9TZIFLdWBIa9edowzT/NIIfmnFXd4dJw9gyh+7uqi8MqCGbFlQpA4DudD4fpH6onKcZhb
/qrHi8jkvYierZpRMjx0ku2tJSWPI22sHFpQFJ+Za4MvDjeC+erGkbURPrmn47iHVnxklAkWUuRk
4SwZn76eFTqnVsdHbwm+BupBJUDhAjLWgPTLhV5naCYq8u8Iudlq1moFl4NGsh3SvcDdPPh+9Gik
HLxXkpXeXm6p74xk6MLxfYhxv7JzquiTCHa7S87xSiY4sVww+B3gasdOw/PANbibODEcIPGPr26+
MEgm/VAyO16OOw98mOT2jqLKT/wsGfXtfLs//+/J1m4zoxWUP0kAi5PjatAWCk7GA9tcFJ7q7TnT
FxHC43Z05ZHZDmKYKxZTYwul2ob5sAnsxTGM18f/krBDgDa9RluEKyTRdzndq6/N/unz1FSqpYRF
RMCkErGs4vFHZqK/atjqX50rXx46RRb/nSezuy6WPjEZiMd1ChBAq+6u5g6DYCqiuoumNEdX+o5n
efxLlN9TUMnxqN6Ha1h9QOPM1/6pBPMYQnt3MCcMpyo5VCd2UyBRJUQxGqjNwxg0tjQwAA/s3E93
DAr5bpw+VxkPm8zCSgKWTMIRaTrx0/9YDKDgj/M2qACVw1fsmAzAyPyc9MXSmdcR+5jzUz9kFEr/
KLk4vp8yZwQ9KajiXO8ueFsR9/ZnAMbev5sa12k9KI6BNDAUx/HC+UBbh/hKXNZoNWiK7/EwZm9b
qy2AgT8li+DZAxfjHEmxZr0Aayk2P2VtIP+T1dMxydoIcLeicamPNtCJpbOBhmJreXl76CrUYaEt
+1RI2yLjYz58ZlmMr6BRwDs/lb3P/N5RJg3nIfOTLhQp/97DFuv33s2YMM0UuiwHW2KJfrNgNAfI
SJL/EIePH7l/iqozokidQU88JIzV1X3wTyW9iAmX9BbrmqMIhztBThecwwQ+d2f4qJx/vQvT3wlT
I6zqQ5zs7HF8DnG999eod3UizNu1TbeualM1VP5yZH+blzva7ODwJNh2Tytu1jqLXwaARo9Ev7In
Ddwl5Ylo1yiuv8frGZDepA38D+H63ODGQDM9yqft+MJCA5k0/8X1f4DBTQ08Kf5HgqT+mrXFawIe
JG6JQmReBxiayxOntg6gSOJXUIav9U3+ZtpkoflhP+VOPgstKol6w2oSdbhpAJ4uXpXpKbY74Cl9
P3JITNPm1oRfJ9rCgf63TPB941DgqoymG13RUecNBsgf4CEMV+ltZmK+/TrntwpTI9Znj3gdnfHi
jQEJzUjvfVl3kc8MOgs69uvikds3CgUq/7yYV84V3Ke3Y7YQHrOfpMh4ndcjzGCMq6XqIkJgEdcV
oIoMK3V0tzybAn+yt+yjPsz5ht5T7QRaZ770QOcrLLE8xmK6bJmG356MW/ZtZ4ggC7HRfskBoc7I
x0pafuvYZQT/f67PtoCpnfurwcxOKJEqwmHjy99A0Qw9MNhWeJ2sMEqRNz3fJFQ6LfI/7DUmOEpc
D6h6sHcXQI2mAx/TEqjv3nSaeRzN+JS/U4MFwtLNa+eqE51EDNjwMrUAvLF+n3GgI0hQavkOttBy
TygMfew2d+dILXLq/9EAkAdrYdh/lZrTssWHhLtlJ+u1olt2HDpnkKq2OFdD+jDXqGjpbosYTyvZ
vUwsmq+lrnrE1TWgQmpHMVlOcIAQTFA8F4rEGp/YqqK4hbH/RtJNTSofXOinNPpOtuV9UUJ7PcFZ
pQi8WvgQNw5FYQOvLQuALlpxxUYnbxwUEQeCRiVt41JfvKp9AZbMQ+WqUU81jSSmmkypfgVdg+Uq
6Gnj4vqrP5kjp0C2y2qQEv6gYdUcz69atcsKVfYpT8sunkPVtptSqadvFnpTWboTQO0pOpu7Jdmo
/V+VXKn1TQWRQWgAnM2fDc6S6/0hc2DJCfvpBdl2YooIb9Xq9b4nUD/TNBFNmiSZkq6Qb9OvEKVQ
ETNcp40cJhtyvO0iGamAsfHCAx+PWlCHLBsbiWkgiXfTk4M7v8fMQq0VdZcQHdxLpDVR/R9WZx7J
qcZ+1Mpv5LhPy4jmHhcytFiCTU5gya/4cj5JcwQrC1Be9ghgKDzf5ofnHbPleQN6CL8Sf7F5vkbH
XLZwPczhnel0JrzICF0LSjC5o7I8DtoYy0fw+IafDukccxuujrmletsZUM41xxsvzAKfunngyE0S
dhcpifFBu+oCe3XULzGr80ELvG5vHjNPpHY2GX8mj6bLJE9ceIN1/tjaYdcLEScIZQFTkKaeFDWD
x6tHWY6VITSTuLkxIepjUYAEn/UyxenkMVey2vLK9lDfkzkUTxlSlUlg7Qc6nnlz/86Hj49Tj7Z1
xVHoBdmu2rLYvEy8DTHWPaCInwN0RjcgFeptjctYAJNFh7HThCJ2tX8ERxK7uBK7LaEbQqsYu6lv
IzlmutYK1aROt9oCQlaxksHAsH/8/rcjB6rYR2crcAITyI9Hw5RfAqx7nyfF2KfOiH5YrNObtDD4
LYhWZ1NIlw9NcWr1EesTo8EKbrYgZ1gOcBasSxXbSTe9f9L0WQ4eqwhOOB7ZpVzdPfNb03kYDQRP
7HQXPQ8N46vAkRih7UWwjYTih2plYn+SIEQwNbUBPrEbkEma66b7YyEdw2WJ5WTLD4IOTWcH7JpD
YUKW+HWHst+QGn8xu1G1PRovoTrtRXvFpOXPQw9MyOF/v+SCNLwsx4IGHfO+Ms8NjuJw3Wkago4V
FGKxjvp0geQv17yEEa3sOITow5zoFy/nM+npU1ssTzMtKIiD+2PyvtOuSeTHwNMvXi/Q3Ao1v3tP
8GbDddX1OGAAkKN8k8+J3MI6hplQqZkW5BuxkAK1sDlYMlOVAygtbfP4pHXaB4RufLDwHZt0gqji
yZxraKwikIEicq6TYTe2UoM8XCJjeLLDEG3nv4JZ8X/tO7/wGSMs7UVb9yBiQXBds4w+TVTOAPc5
/wLUO4tSoKiAbmZzDmzPwNoV//u7KPwbxUjjhx7jryMRLFMYWm+67g9Nyhg9WNanH5j063Yav3Qd
LpmnUziF9ktg2OmA7vX24DASUkxboVbQ2ZfjwwBR0UEKYMptPf80b3cEXUeBAsGmkHS/syDvZ6r6
+4HiP6D0hdrvD9KjvHng4kM7cXyu00++bmB32I6QZqmt8ykcygBITOey8kdA+K1YN2/Fpb2Nc93e
UsLNic7uAlz+euKFDFHuEMFeK4e0RLhhygrlZZ6lXKkvboldQNzRDkye7fc2IImJNJ0HRyC8/zRX
79cMqaD9VGaPbpDhmTQF7T+bUjj+tzT3HXK1QxLybUeRE7O/G4AluHnFTPuyedfrK0Ocdd76vZd8
2W0k4+wwQ65e2RMXFr7pp4ivOpswVuRq03EyIGoyJ7KHf8KE30+JmwDaQlm/yU/GtYz99ynXBLYn
UY7VpaIpARuipJIf74/WcVo2dHnMVHgx98eUxiBD+fXIeqvjjS7UzyfYfGcnY3K0tMgefrkoSVuq
QaGHbw5f3QbKQPUfAiD7UYemB6xJ0mbIaAuqWARS4cqsUK7KE2DHy28J641KR2N5fINgT7ZWfdk0
a+aJxHVeNKR+xFtaIlzcjJVs3R10x2DvpLggZbI9zNcT47MMVm/a0VRSULSjVdyL/2RvjjFOpClJ
dlZqusW+YTh5Pwm/FxOQo011Wf61lsXBLdVNv+h9pAHlgbAIU36leF/XHsbYGXW/dIkTPtTjado3
ZO+hGg2fZxj6rat2aIuOzNLtRVwd/Lkl/fTyMT9HLF0LzkEEEkrwWN2QJCpqg/gLqk9VVT4s9EVs
Ke1N01aHXUC5cvb1ovlPLu7YUmyWkK5jHFGsmYIwGmlZrYnY4tYj9NHSpgHkrXv5+ieFtn/Zk7Z2
S+2EET1xHFZdPUUg2CypmhGGsfjuj6kXBE+OMT/A2obMzXHFaPo3Tou6tHfwGMdlyKhrg61KXI22
gDcOg5vPpiWGK6Dd9Prwb2j+xDkAchyJoeS6JTAvB1vkfrt38A3dZL/0xOVZCQ2YYJhcsQjuEdS4
NzmTgxQ2wMNLHAiPC7HCNzT+o1bKDqmXyd0KQnvjorAEdZmnw+bvKu0tBBB+Vneq+Y6ZSJ1zjXu+
LPfTF/tCAqVTkWJVARxwpJt1aAA28gpkHogEIDr7nWoCsLItl7kFNEwXUAw63of6TnkEOPgzJNv6
XCgATiX6gqRY78VsTp4wG56Hql5qQeMbOmqzYkrm0lFHhfLNZx09FWcj2TREmx9ExV8jc8Yz2COS
I3cfQKy8TIxmNlPg4WdEOdbOAa+aYmDt7OAbHxSd651hNxLBe0TT7/w9AvqlM5xrK+Hrr9R/nQ4H
cYapwC72E/ZhjEFbnfRbUIwe5lx84+/qZON+cEKxI6NqhFaZSeX2S2fY6GGRhLYScGVG/e0M3jKa
5lY/UzDXqxYqVe1Do53xoqu3ZsOeeubw5s1OSKWmnYNNOnvxvDUUzVtGlDEwH6fLIibN51pGS6qe
kZQ5aU7YdKhg0lTiVV2T3IAYACAFeH8zIBmfzzQMgBy+JWsZB5Kje6dGVEb89XQsJu5o1x3YPb/X
UNl+OIU8Y3x23raKJK9sTWRohEXhTywa3XHk/IjET5tRSiGw4ZT1cB36rw0/JY2T7/vNSdRwDPSt
hGd28D7YhJ/wRK4wQTEUSqMbdaJbLyVun4A7GproVzl9hK0Bet1GNn6OuNKtpsLxpwgi6chDK7Ou
P5jnj75vUipUGSMCxRz30aLCk2Xwm+1NtmT6o9n+9xFb7vugtr/ghw0RDWaKFuBoj2ahx0RjuF97
zkmqzDU4pGQBaaNGSeVLCGk8j42Dm2qocbjjmxeoWcy32ZPrLwaXCRbYW3SJlfqB2Weu+hvt6br9
ysDjl4HLGlQsBDlS8YMdPomZAqw91WRTDMH9JDN25wp6GEc+RB1D9dEYNnSQo3O3dSCwqtd+NKEj
gZOHBlM3VDYbSHHu8EGfqnMinHQKaInFm4ETSZzjjxWt6m2D/JTw63PsfywEHPBEPt7qJel94CKZ
dB4e12/lcs9WMajDqAhH5iS+RH+ipT9Dd9x9rJ72FnA7enQPtkSgBzXJhaoI8Suv1sXjZducw9QA
cKLy3ymNQMx4ULeP8PhewKP/MLbHEKpdq+CVlcHMpG1sxjlAaoKXVEPD6qXOW1nBe9ET9JAeEhvL
GBxPo91/x5kOz8glT5qPh0YB4Y8cN6Jnr0CrUKYyGLGz+Q0cgrWIncEln1VXQMkG0zf4uUXoVlIp
9cpYQQq81LVSeq/bNp0xPsJUAuPN2V1eU5fpFPeO7aEHH8PipNNCTA1qZjT2tSc3xS0xAHb8RnVS
zbI91PY6BxRbQriouHM09TYgWyPVptZztnQk0u4Tpq6XSQC1x/C85oF1eOg9ozU09UNXPFHHkVTD
coRqrkKrePwfLisBi8UNljGBfS0jFvUFAvApOVe8rJGsE+jNXPlckRq7GgRpqK72gdocMu297xKp
BXaEuAG0NDO/fH+P+mQ6uvjQanuBpj/3oZWFFWEscn8e9bc4NDftfNWM8gz//T6Cjfad+5vH04MZ
rpc9z1Zq7SeV+VYhG28iqAXrxmuyhXHxuisCwXs1hdkeHZi09yyI+9WYGmnYZihPDh0qOWOP2j4t
1XHX9zgOpCsYinNxMa+irttC6bcyywF0ji56PHXz+ADTsyYo7DatGg7KEV1tcr+i4sjkg+3g0+Y8
vkrG4mc1yeE6ox84lX3nfUduVjYIlLNfZnM0DfNwAiJYnIzl0jUYlVxUCbX41TEyIc/IVyeLSiRD
2ci2S116aZegW8SOp3TQOk62oCh4y/6ZogoOVnrzbqc4Ubdc72YFWPdx5MkDDYachWQrPRexjrbK
oZQ3wvuz1PK1RS/etn3uSIqZt3zFK27P6oZ61cyG5aupw9S1adBqNriy/bKauyigGVZOB/c8ayjK
0yhOBcT6kBCfdT+4wYGmY0bMVwVz3HDQyPgIe0ZWpmGk+wzOGOBt54J68VCt2vChko7Uu7LrJ4UX
PWUooaTydY42XELxbyBROp7eaJUVSorzaU8FD+5ih9oUsEWFqkSsfnkrnECX3GWrsKoPXMsz4QG1
2sBND6ui9ai/GIVNB7Ah+m1B9j6OD2qqP94VjRQ1gb0Fv0zRy+n4WaHVuXHAk2f7PC8kQGap3ZnE
icBbQ9iZ+ZnbaXyfL5gItB2M8W+zTeTv3Dm+M7VTWwbJSxU6DAkqQi8y1b9ZKgYVtMJsGEEt4Cvy
YKAPIW3bAVSZRSN2Kko70nzAx2YEWQrL+/k7XvK3EFONGMlnBVnzW/5NvYIggzKktOODdhDTiv2a
tMGbQPcNkNUPchd+NKuVqmFE6lNJyPdMsGQZUNTCz+7c5v7miJOPxbdAWmAZyDclqNrQjzHBQBCF
ZgU1zxSgV5pta7HwtaVc4DRl/B0mFiDEruQJG2ANOptgvIOcj57VzLWRDT9/rMK+Y9BvZBjb6d3+
lqcebmCKYFyA0NTiwN2LJ1hgQn1qhjVoEkZ6vMjQX+aX16chZnniuSPtlpdFJQVVwiparHF8GLak
A20LGE/wREztTQ4xwSRcUwKGaf/FaU2nzboVJOMHBHOgCQP/8LaIrRv8Z4YaxDm3TgqR7WqJET7G
wkbVTaz8oCQYvgEQz6az1qAA4U+9E3SDhqvAekw7l+euOpRI34ZPaZoYRmuBTE4Vi5bhANKTRJ3l
BGqqwumHaG61NveKlq5pmLSKaqxQH5lyAiuRvcujnd9F6KPJbXMdcYOlPFeGDaWMbjNhiWed+tYA
PF40KalpHnrxNtqcpKnnXBJqBDev9RVKcCieCAQb8EvR/ogwWDumV3B798X+PxldOLG3gLek4n1Y
p3rOUODRl6TGBztx/5BtoJLXOFvpLbkidDBgVydH/0LS+fo86dZ6dcQy96MDeyRF7jdaJwYSLIKo
l3q8pJ6j0HPmCdwzCovHoQ5SZ2LxcbBxZxexdxkSfePtQY04aUgUcNOgop+GMwhdV0wPF0kTCVoH
jM8e5UFMUQkY8YwhbOYC3AHA5Aa5r8Ye0xCOd8IuY5qAnjpTsQu/UlY87wKEz4/nj+mwCUa7rU4O
nxnyRDtprFgHUCOUrnXOflZ+BdajSkfPhk1cCWP+yOouyDfqF6uOGfzD5Um9F891TMyuwKoK5icd
R6sKaPtpHlVFZlSf/hTKUpCjnHSETwUu79cPADIaXUGAtGORv8cZqFK+daO5MA5kG/ztBfjPliAj
DDfY6ENliMyGZZRuAYisvidfzEBzlJXd1ODZ8Tci0rduHK5EsimGGEDGs9Xu1ZNnCG/Uing7cvjR
I7qFL07V+a+OsMyIsmx6iekYjdRZXh75bgtMI3hnebStVML54bPuw0J3nGfe7fSOELtI40LVJb73
p+dDGLLN8yN/IxhFhiQPbtM0gv81f7O+RMxRffrhdUHHnB/j0cJ5tQi0y8laf3FuvHBVjMwii7K2
Ol4fbRF77JW/u7fqZchtSGJgjbnWT2ot+717dhyRNY4TEZlZ8Xg1OHZDIZ6NP65slAF4D6cZTd30
c4Fgpw+upVUCJHWYJ1wiO9XJqMatd1eovjHVzOQE9RJdHgSnhiyNteIm+KbfSZ5FErsytTAeLSh1
a73ulb/N4cp/UN/9wVqRcKRS48v+FjJXuqw/kp+s35hNUr3hNp3ghYB7MkxfveMpJCimtbhxzcSS
UOjsKGyBxv+dcDvHpASdmP4ybn3I8mNY4yQkPBehDIo0jv73tVVkdyLqpDy2CpBImHWPC3KeybUg
4w2yDREbMjI83mcJMQS2rSxSGo0wMKyObeGz+hN1bImqSl7+t47FhjuZEaaTrtqp+4+Z9vqyaEx1
/LGsyjrCwS4aKCwVnrOqlES+gc66IBLVOt/PvT6Mtk8qFlTp9dBPJyQRJHUX3PBOjnYr2wqnLNln
DDEIx2YrQ3A8fJa3qdRZW3iFq45Q6B8NcED6677iPwaqKEAs2VD9JCJDeRad0XPPcfiCkFzgP1KM
3UYT0Bi2C7ER3fil6EXkuSu3cPvDu9yPiczzLW4j+pY2pT8bN7uptWkOVjQk1QDdJ0hZlQkBZobQ
uU1IXW+KiWXkeiw8qk53wvz2DlYr/49Mquum0FNA31HAy+8O8RuPfxNm+8vm/MVncBlEdJU3NPZs
muzWQa1jt9yPfEgT9XnO6NNRJBlFOvIqkHkoIh+yL+JY6toG7oktf9tJojJGdt1spMTF4dRQlYDN
aGMbzWrkDRFJWJxLn3knZnOoiMBG4gD50wP8RK5dev0InT89m8rXiWAlE2oIWbyqmu2lbhZU1wux
NCOrXeVRQszuiwkET+O6xVe54JrxNpXs0XI7dU4qy6B+cfL4jky/vFS20FXXq3tAV5fwOxZFV0b5
VgcnCyKwuSN8S/cW8BI1lXfI4wrfKwkPcGvpa2tCG/c3ysPvo36depnpFQufZx36+iZ2a6YsEhv4
g9lLjgQfG1RbHn5jHnAfJtesWZPCwC1zRd4hXKTDK2HQ7R9JXOvhIBTOnH3VmcH8I1NsNJlXLBnD
3aXWDImMg+EOSCF3+4NeePmPxQ6dQQVw+qTZ6t1/r/feJRVU4VYXeIBl5tFqp2SeOd/CsHwmpTnF
ase3JgDfAyeJMJ2M0qq8Gb+dNQmue+EuluQb36UyvrXUU1xczlnTTNqJtnMRpZu9sOpFkK2M2lv3
eKc4PDIxqfOEnEXAfPyPhVCnyjw7Fhe5I4ucxHlsYGBntG7H5jj1aMAjVK6Mb7g4xRbLZ3TZN/On
e7Z+f5IJ+6CSwWFnqEf9Xch0c74sEWaWZ//O0pXV0o5OxMjvHB1EkcBexL5jgOuY1AqKBbTTxOAJ
4jbnOsuG4wUFKVzCRijveFIZtdwP74OsH9FoZfWIzHc24uroam755Mqn64A/Ho0528vWcwoX3a6b
lCFZncVIcksm5g7EmDqYK6ppO25qe1aPc3DZkmDHc3RGr/5g51Klmpq34BXoa37eW/2cZh9MSB2e
9qyZZAuNP7L9qd0FC5caKrmCPHk9OHRfGyPnWnRLkmCv5pfZ1p6K9WXm0HIkfT3PzYn7D3vMRdBc
Pz+SQMm30iBt3IMc3O0IeruRALyLnruLFyfQrV6UzZz4ZhPsFYaHT8zxDay5+mARKtZDlB93WoDu
5QqCvj/KrV9c74OhCc4TVHtD2JfIz0VZGRIFdeQ1XIQu9Aabs1kSqBXg4GHYHxGainZnOCW8p9Q/
6tVSWs+PJRQaaK4ZmKFIsngnfg1KMxh7HL1HbDlf1UuWXvYZWU3mDSlwCliLY6JYDj0wj2Lv+6go
aUNzY6LpmysKSWToTZD7QVkmpC2bBMFN/SKWJIjbRFCph67NEU+hV/+JrDNuY/a2thpJkRzeSv1v
85xkgpl82+BxvvJztOyr/7XoiOIIaL0Sab0e8tS0W8nba54ZA1wkZxatHIovD15N6DThtQxngsEz
feA0TvmTBx058BlvMPqYcVouX8PLAk5a5NoR4cPv5yM21WZhfazKODUHSALYqHpGA1TldvfVt4dh
0vfsO8SY2pI2sDHaGrzU6eFa7fEWc1iniybfbTdbaxbtbo7FIpnezCS/UYiuTSlZBRcWuRquHEd6
YGuxUspEOOAh1hi6K5SgdVgEv+Y7KaXBkY1qSIhTmh9G5RpnCDZi2PNh0ybTIQlO9ptkLIRpFdzx
t+Po96rlLPb9sIDCYtpJpUFs8ASHIfAAAi98RcimPQWl6Jy++uFnZOnr2OKqsInPFK7hvLHPf9Vx
q6vqKW90APwUi7eE8N+Xbfvmqz+8lV4sy75RdYPcx4XerWsm2Y8aLWv8Od/M1wi7l/Is2JLffv4+
7KQGJSVsMx8nLo8eO5jXkQmd1NGrOnQqhrIwz3rvUVtu3yMoXkK2WYUM0cO1w8o2ykrF9NvWq8u8
cV+arE5Q+jiX8kBd9tiKxNjKSWCqZjP8prIg2Wic2sR6eaBH65DPvRb7nKz1iOyEYcL5JrK7vcfz
lnQJNfOGYcJasvQokkwoUQ3dS6hXfnzaurjIZya33EUhLr1vd1FUH672ZTw9jd+kxhIj8XT1gBDy
C0MgWuD1FPj8tzGb4WQWoIKrxmFgk/IWU/oRjJP4pTDl/ALEHIIjCeOZAPTHU7J0bDlpd7ecsGtT
hAYIz6bOqfRdaZsJpYFjU2FGPbGeseIw2aJ5H/RlxvgqNnCA/tMfNECzrRsWbtPQiYbnGPCE8xPS
Z1xAczNyQmY0xntKX1E1+/wWOrjYKV6snXQ3Es1sGJNRGoupsQamWhVpE32HJog4fyVNrQAo+0wZ
gD1u9nA6f3lESY56tFywdbhnfIOr8aatAArIkhqbawEwoE3/PoW4u3ho30gdU9GHzMVm4fsNWPNn
G4FA0wawZ06dVtZTN0nNpaeYE6m/MVwib+bZKNy2147+74vVxpaMpEZQ04Hch/vdv/AiSSuRZdZH
U2cQqPhnBFGyJ5aN5Bu3V2qlECB/es/bj2en7Pbbyf26KPZ7De5d9gPOfQlbXVzG5w8LLMaFxy9U
2eADmuqIWQJsRoCZ9wErCb3wTw8mLvJdbtb11yj7gnHR6l3RhdGD8dWKdXo52/KyhxAsgdH/sMZ6
683rlqdNScwv/Scua/GEdQAtxPerDP08sMvc7Q+7mUan+jSCumXkOkQCPcZnhkfr1Dh6tn65nKFw
ouZ79CwjBWk2O1NompmHmcQptKZgy/rptfpgv8clktppXJ+iuqRZurT8vOeb3mgcxZZt8xeRNuoz
Nv2S90EpSkAegKE659FAZqWVpc6kKf+uxL/WiMbeMkLZj6oR54yxzmKCyb5RQZpWFgPPWjo7jYzu
hn+R0JRHVS+fSAX/7H4lTQqfKnuUNURmBAtKfLCogutzx2CSAMZFl2Nf8sIZHtPKPn6CRzAYGYUd
0oYDYwmVEfpts7J4zpuGHl782EmGaxmdQ3c657VtPf3jiVS2A6a9XC0ebsAe4bGqbWqkELKwvtHC
BIbOtj7CWWdaSbILX1EN24oZQtlThfgdgKyRD+e+d4bTHKxY1QhVXmQxhabfzoov/IoLN8lyvuRZ
UZU36gwcFgAdhnafLPsMigqHnu1B5b1e/YRSNfqKLW11ovuY66leITi2vc6zUYjcTwHWs+uivBDA
6gnNtFAQWhNZkOvjgWf37Uzd6nHN/MGmI+bp6O0RIUxc75Xgt2lIf5E6wt03QU48Ms7G8SFI23k+
AXmze2HfALMVLZu8+GkUtr2ENV+jHnh91i8XM1V76okXD65yEL5XjA4/Dx/Tcdw9+PtHC+wgXm5G
adqlCvTa2kn2gjb0AEjvxl55/PiNj+2gD143rx+nk2q0BgtjwqeQ6Ayok+r5mQGWBQ7tnDHSVH0d
H6S88NjXaRjLn9/V0Q9+M34t0Tb+pHiR7ljgOFUlM3acw8EvriWf8wPQLKFQhvPaxA5QeCqznJEe
TyxaaaaSA32bSVZKBvvdJOeaQtDDAHc4C0wdMgdGr4PT9DlCMn9dvOSO80sTAvGZFox6hzhEC9B1
9qoRYb7KtMZVm2SHu7rkryQYUtysQ8bMytxYSGIx0QqRdU1snv2YC6+Yu4XMRUoi0iKvU1k1jn1v
tfvH+PMFyor6ejqceLRBnbRhHiO5Ah9lq62Qg7di07EoJJEEWTg6tEUKwTpnYGTTZcEpbwkZ9WGh
EzM0aUWElFoqR6b2VdTL8G6+AM+5BKvNFUFrQXjLFkPA7oiXqC3AS9E9Nic6FMbMKDXkYLxN4tuw
4AJMRPoNs4Bh1tgziElsymo491l6be4K7pgh4RK9jlasSdZDl9ydjRzXbkzhqyTrpRUemrnVVJtJ
2gekng7RXJkDo5TzyLtEdloadsj6CuoQdL1smHC2Yd8w1wcx8FxW2RdI/OxJO/r2mHafwPsZhRf6
nWDjUGhgW9GlupwudgosZAW33rwiI65aw0KutxR2AA6BZPWuYOYn9/QLSWlVcITQ94XDnAHnZrK9
dSyX8JkLEkrjEcQWQ4MN7lRdGukDSfAyHn0MkA0FSBO3lVxWASBSgtgt/SXpWck1Ann/e8rOXwuT
fMYPP/1xNzYdU1/U1NaWVNOaqOsSjieRed7cQd/ND9dc6OLumZaTAvK+MUNbSATeMHXyuAxXhxgp
4sNcaBjFPRh9Qfg3UgOiTE+8HKsYlKxru6PSORs7UVnjFVICp7ZTIPbr3kK2VWC2OrVGWiVFz7PV
b/FlOHaJZ7DPHfpH0XyKOzYeUujtM54lfAj2Qs28L7DoXq3Wmy31gvRScNAoXQlovXgY4dtqYHyi
/CZYBDN96HDL23TBTuSK6R/j4TW+r13P9SVVTjKh0bpGsKvO0jbVLD/SDOSeK1k8s/kOYAWG9lAd
SqA91jnecqojlNL33julLQQLFxM08dndjnZ0KVx1732daGvU87gdi7BhNwEGEMYOWMxOfovU5Apf
ZgGr+5GusZD2OmgWhelW61e58/GhDq4JBVhXb2bV9UaNgkKdlUfIrRGO+/IME/vd8jTlDikcNxOO
lpefDKsajVQOAFueQjXTKrhH9dU4FA0T89/FhvqTrzfKqG1tq56hQXWeqMO+VPfvClaW1OFaSVYA
uDIsPO1WJ0fRTrGy9OVJxOqP/qG4wLXvdYQ6XWi/y/Guf76fomR2Z8xU17c+C5jnJZrjnrtZflK3
Hfo3pik8LVw3putsuH3Aq5Rig7KgyjZjEKqheZRnF3eVK+YdfwmFSnRHQMeuU2ypOOSQhoj3TKGq
zNs5ijMb4I10c8xu0nhXar1ZoR2mWpNLmTF3YT94KxwzqfRNO5P4mdZHKOwAb0lbXW8XPYin3WiY
mdk1a3cbo0A20SuF78+JVUXBjdZDiEcqDQFYiGJ5GRTkG7Yxg34Mhp2VoJOEEHRkKhWtN7YFzv+a
/fgnctk0ztEiQ2CUZNmab62UPCnZGbPvnd0/XxzsYSBKpnxvGiIDDzMXdIGsHvqxKfN2W9+2ZA1J
MW5TFHD1g6j98IUhbD/Bazy6TUpebdokFMYNXC6Y8mXn8vO8ZbYlk3dK576aLs4+IhNlK4Ohv9dQ
rOV+umsVIPM3J1MFbROiaLpFQWJZRCwqyY4Zu9QT1EBE1yLii325o1eDmh//nbtwWlqlrCuZ0XbH
1QM5vEPzhTBKfJ8ia2YrfmN2gvU9wdGpS1kORi5LgdjWfepeSSJ/fkDSVJ+dRjfYsJAJyuYuV7I0
7grxW15jEyF7/sYAtvlGgIFM4pl9k+2SdBJF1W6xjozLfXs5cO6ojSkWsIu+I9eJSO6kvMrbeGUp
lhGfrvsWqWjct0urGZcML5cbExnEes1kMSKnUfTMfMIYUy9OQl+eO76H9+lLsjs3KblaSC1lpkQK
cY9SxyJ+mkn4jBR1AN1sPjrHAJkk0/2jcS3KkJtaASzKNoAZSc2kxiH06CpDvDwYanjZrHATTne7
vKo9pW49CsiTJ+pATOBrVgbiwnh2NECBQPjixNqBZS962vOWFT33nDFzM1GB/Kx3SEBK68mfU6dW
VZsXlsEwqvpoodDyh3oAIyMKKLRGF2PD+jblJMDi1t/rxaukWX7gdF5AMmTT3m0zAqhKQ97IMh8y
fLr81TuwLVjHeRjNg4VWakpd2IEaGo43VLYVy+UANa//C/Xek75asBRJ0TH9on2WgybvIhI1/U/R
YNArXulzYWhAiyxT7SHtn20zPt79SxqOqm2i7Mq21ApZKI/ftj3yXfQU/cUFVeZjmWMT4s4pvFgZ
xL2STbSG6dlTzxp8wqh99DKXWea/mID+uDRn0t0I/7jMuK4BvDwP52TnE6bzlhD4/ZVjdvCIC0rO
YQlQROCHXSK/hu+MQsp3kZnPP432O+cWnGhyfzffqr0IYXx14kMlhxEFHgl3VeVGiJIgF2OtYyYQ
44WUFMPtRL0B//O6I/a2fv2o0xxItiGNzb9lAjkBAMoJXwi4UICJdUHZbSFGdNHd4yJOJymlK6Rb
zJK3mUYsRMiP4jfi5HNxvfUni2AjO1dMOGXx4KdM/gJsBtq0wgLuD5UAmLciTpW/fRMNeYFOjzmV
h37MGfinbhQY6MCKKEWbK6UmRVfxdaC5WWJrJ/+ejf4FniT7pPYWcWPBPHRpI81OupLfRB5ar/UI
uOpUEBYAXXiprXEHNHQuTznFPRl3sCDhfprmE1leV+2i/u5t7LoniV8FB7QJNKivM18j+dU08aXu
R+iMdKAOUpZz9egjimOj9xVDGmQq4kCsenMMez07OqWWGFmGsg23ZmQo3MsbfhIZYg2t/KEohlOM
LHZ5Cvz3NkQNp/So3B97j2q4stjGYhqhLaYkAQlKrI33mc9vnx4oD26JbbnnLuDgK1wGxJgHKYeN
4dCMkhMPfwaaOQfHmMJBwtqXEhSEARmYqJvR3IFlo0II8StgqjfImUo1Sz6/73sgJ/qjj0X9pNcl
wxQBQ57Hr31rKJXLSkEAkNVxwnhwQi8VJAB2JxDcOd5itmYlLT5RhhYuGAnh5X00sG+BJmHB/W2o
Yo3OyYjWXZwfnXH7LHMYfq4yxks25SVSqzhx0Tiwu7r1RnjokJS5hSApMRZZAw+mZ9i9j7IkEOy5
YPemI0+0z70Vyt7Xx3S3S2x/EFqxH4KWe8F4sMWtFYqRkgzypS2ophREVA8jhD0ozi+Siv/WXsyF
6SC/no+jejGqnwzXIlADwygZYmRvfs6IJ4KSX8u/6Ehfh7QUgKwUQMQQVuTOgees3DdGmEyjKq07
fwJ8/K7z+A0FSjc53vmptpCb4SkU9/CbVir92lO7EfU+X//22qTSWkBdMR+sPYx2THmHZvTTX7Ky
0O4hdBaYhCnAeRS9zynA3/rdykQbKIR28H7o/yJJRt1931Pebyn/9ojGwFQmAUBSMRcrLME676fi
c40Ba9d5LYBtPRgg2r4O+a7dimvQ/iRKjndujzE9HfxHgnsKiQtVWMR78FUJZrzsutFh3/AJU6Gg
y/DqGWPO2vHg/sqGXFz0IIiv6um5CilJdyR/g3bZSDAR6sGpHXW2LABWEiQBuz+DJupY2g5iu+f7
0Wvfjm0t4Nm8FFWKrFVGBXtiMlxSWW2Ep7YbIUPa42mCc+kZa2HMpRz0P9YrySE+oj8xuWPtW0pf
iEBq3UYP2j7crWLYk3fewh7Qs/UPdqz6ot9RAW9q43BIirTVluMbCPehfUVaknkgauqhCWkLeaFc
hDfMQq+oWSvMlRiMw/Vi5gTRaPKREkxeb9fBGIK184b8NTspHpAwnmzxXu9qAiV3vj0XPz7SyeTn
O1lqvJ7OUgXezynisWCdtkNr2eFMPHxOQW2uijjdEuyOVh/P63xpMi95fITFE761KXSGH//cKhY8
TqTpV7tdZ6E34jeY1+G2ej+R6Wyk/Vu124ggHJrLRDO5QBhJ/BYIqqaQZCgtWTSjS0CtV7BIbCiS
ue//oNCN9G30x4ZQ5ivUb+KcFByg6lixhp5RfgEuPiyWtTKIqFz0N6o2GlBfnJR7Uel/uFmZImUL
NcZWOQSmQyMWqBAAkOto6Ypv7JJkwVKkatTVNiO9PHP6e9q/qqi/nUXsrGmgJjRzHGBQUznzQYp2
GniLr4k6AZnYlDdRuSyFlHyDd83Op81KK63AjMA2F+6L5ylJcr7m28A8QCCFysoBoMghhwBJe1Lp
0gwyQfJ4h9vSCMnAxYyIf0okk01Dtl3tQvlHLj2OjPULHQ+wjHNabC/w/8Poxo3DW0cUITCTOm5x
QA0x8310qnxOgO0BU+nYYqnZ616Czhvr6NIDwTirdl6mh60GCn676oOKwDi+gr/fs0yn+qT6mpVT
An6V5aTRuNhwQMQ38yWoXDblH+Vy09t0zeaX/51zLruub3yw6ej+VnQpJzaq9XhjUZ+oGPUv5I21
bJnitlRkkUNGuDmIc59GTt+myU2HbYYAHhwtCqQ3TEVugAFlyqMS1MAQd7iCBokpCNQVPY+MZx8i
WHawXfmkaGFbCiFBjf65iqo6WepMYkLFOt8Ux2degiSUIOCJdSVGyxM7NrKqq0yDxP3SNSlERWir
VmafhgmyMtvZx1SVudc6CsgY9tzyODKjPHmI+U9INcCDDgCrUsGRYf77zRLZAwFWEvdPo8L2BRpe
IV52NPjPugpYP5VfLcbyvWqVdJL2JzUSdiZh9UseXNOT/PdvpCglN6sjcVvgo5Zb62Cce5p88q1V
ZiVgSGfQCfQ8RhU2idYzgTaDzaweAQ2grVxkoGqkw0EA8myKzI9X9PSGMrVm4IFCNQ0+Z8euo9ds
QH+NqENeKMUTOpkvLGYc4Xwp68S6EK6+E6o2q1sgtkURtts93k08Zz+kdfXvtaqdlscQ0u7tnPhq
rvPJfGn6udvI0+okYUrC7V6w/sKvQWdntTTJyRXkn4af8f0KPma9f0tW0UCy4pe7FEFpeTg4XQYa
MNatfxs6fUHTJVu39G/DFyxTUXY1mrmYMJHpSN5LuBxQT6VElDRRJEmVOLeWIC62tASIZQ/QbP+J
zrMlSTkfU7Fd2OPBRaIfiBGHUqA3m+R7R7Tol3EI9I738+hYGBpBedJv5+CDkhtfAUs7vBhpYtBR
IhJvTBmzJAyrYq8sQJiPfRoXcZffzJ81tcNPOPMQnR2Ddm5gt6WTS65YiikZCxj1551Bij/RHCiN
l/4acbdEV+0xWtg4db84P17O5roJqgwNU+1E1DTeZTyuSFGgdj5YWW8M578wILp6lcjzzWUBxn2C
8u13V2JASox8VsJ/lynOTJxLCKd8wZ45ycYhQA/cTBXwTmCOF6s9bHIf+c8apkVWEa4RmuRgZ7Bd
RBEG6uf/5xyxVhU/nsu81Wcye7ThTsD5yNld+xni9/Cq8gCLZk8l3+7n+50XJLC4iK7Qt/FKzTfb
Sv6h1cO/vOFKkWY64fA0tCgUaAe4te4CT0iBP8YOd/xKwARG/MARASgdP8wbTcVmlvyXuhiBr7D7
jKySQe+KNt/Yq/BQypg6xE/ZDMktXtSK7umV6lO98JbBTvtCYlypckD1W3NCiznl09G/YyYqf9GM
pbECXI8sPAkslKBCJI7S8KLLn8UFDuxcJHF7dK0h5RpX2dCOhKodkoy1Xp1XvBg8l0wARVIy5EC2
ANhS/s10NgrNVa8MkKG3YitJ4ggtU4JgyYwp+w15bOqPMgz2/0jgjHgCnuK+d6Yr7rpEJtk3Dnvm
nvKCpTgO7ymPTzbEiuU+UxT7dCGtFCdKIVcfON0IFt2H7iMZmTSZ5Vhumth1kXShqATc2huhXHo7
0Nt+QoF1+dnYwjTWNm8E8cvlW4skQtnKoJrUlyQsd3nd3+r9afBIwJ2ZAirc8ALT4rH9MrHM0/Rh
qk/ROYSkIdOPV5DfMJuP+RDICvZUvDYO2oi4WmS2rYhy+7A0GmD8fs3nidX6DDWa3P4MvgFKZOKX
qCkMPfGlpkz+s3sP+k9k+p2bEWKk/nsnB/Kqa8DZvUAkAXMcjBopTU4QiIwlNTis2oQRXgzJqgOD
LvFWF6I/443JeyrRUV50ahoIn9PD7pnp8xcWyDNaKOHDqc7U/ul4eO6CdS58XK0loaaryXqFAVDK
/iTps+LpxvTZI83iFMAllxMDeL8UtpZ2h/1TG4MOz5uV2Jn30k0e+SKkespCxSHqdvH34EV1xatv
tnhGsSIHstuVrHLT/4aHpWDYBJJxdSyr19ILtM9x2A0jSSCzT6gmwIl67f2wWBS+SP3WVE2rTvjw
sqJNW69UdkC175Rv8zyGize/Blrz85FZWXKJU6WUJbIyWb2QRiIYnBG1LEuaPsnV13YXJHf1uGWu
H7Wx75jUx+iSbbCic8nmS/ByDg8AWFZIkCc5LZn8+2cLApfpBdpwiOIDALJseL/tukWDS3fZ/Voz
rt4lq+0Q5Dzo6vZg3amx5NCuU1f7z2Mi7PDSzWA01mInARFwgT3wkNWJlQFzb6ZKn7cJIiNZHQMi
z2DKl09fsCPNhIx7AQ4WcotH8SEyzwiRDgGXpYY1DgHB9eNF//tSWGJDIsB0IlwDOS8RbjjgyB1i
b3owWdmPtHoKAHbIhPTW3FsC6mNFW5fTLBy/DvMIRKWEc5gzTR5bA03EBWKy637CHrW8bJAgRTNx
HP2dpnp2UXJgMw1g4zClHxT1KkrkXQfCuTdDGjRucUqWueBNUTTctZi00HOcB315eySU+r2PPPr3
VejumfXcHXKwGFvpk4sTskUZquSO+OucKDzpHzdK1d+rwLwZYbCu+x2+GCwamR+x+M6lWnmS9Lt9
HKXQwueSQl4cVR015hx4WmfereK842iEFk5S4iuKsiWhLUhw32X4tOliohLCk6nLgtPl6IiFIAus
MNKHKMBnqj9VyKst+QhwSKe0VqTExpAxDjv2TstozPdZ3y600qnQR/BiIpTlzSb7HZYn5hG0DitX
tl/0y6zOwD7XrJGqSf7tlcY3Au/Yw0e8zi4xmZJXbYE3cJXBxc61F9KECbxAcAJZtNW4OCegAXnm
czPgbK6sJ/l42hy1HumDIh5IJouq+/2wsExUIYbCjkJxGBOQfrCEWYo3A7jEs6+jyQIu0Wklrs01
o5YiZHp0F42J0yyDEnu4GfatjAISlcZ54xc9fLJt7/SuFJT2g1aaSFcasGRlow4r+snL8JJ5az0W
b6n7Ap6QHbmrbLbdPO7yNQS6aTTshX0QI9pJ1Ycl9C6ILT4m4AOVdF060b+KvaJSKTuqBSux6Zxu
ZGp3JZ04nieI2mOnuv2cFoRoPThzChCklYaeJRonAhnqjcyUIvVoE67ZNHgHqI1YWTNU3ZWMotoJ
YJ1Hc+9NgT9lw16+F5J2bx8g0e+HghsK/6E2onm8NA55prDi8B334YbF4yNXX7syN/L10Iivhjcy
ADHgP1VjaKYaY2R9ClnFgXxToFYix8vhdQpVGn5sJi7AQgplZLi2m/ItpKIdLbjm1E7YI7Amt/hf
ghhfcPPcnf3MNkYbY2ERaHJFv2qScPDupQqk2/8jSZBgrxRwpYT0OZJ9A6xDuoualmoC85C5dssw
28rNgagphVKMnZqEV18OA2nXwGA6C1Gn5vcarfAbawpre67oYtyM5Ydadj+4POoJe1g3SbD3b1K3
LlFGUtLu5vMWsEuqZB6simL9cLYdOAt+bwR8qjTQdTPit4Ii/TXzaYspTUYgUs7KaITlfzkxzPvJ
WBR9Un8n7/ZAx9kFnvtGZuZo4galTODk4502ZkcFIF+Bz2hEGw/xhhPAxyXTH5iQ1AIbrGN2/Y/f
pjCknnHoSkedG/2j3YBucoD7aiVXT6xkAFALTiFLnjg5b5ABFCvqqs4gJaqkBSwNNPcex2sJ6ggv
fhpeJLdt2vS6pjnEwQD6pCeSYXuYnHw1uIKqipeVCDCR6u5X4fkv8t58vbruh7nvwHwZCIsZp+tV
ngavhQwh0g3+CHR0aDwBdaGpIkIsVQSUSGipqjrw6S0aS5OozxHkBWUfyQ6GH4QHAlPo6/p8D0gC
/tLxCQWhwuLr8KEFlTdRHpe5dfX4PUH1ZNSAJIZ5+wUfc3/KohBCP7/L2TYROL2DdTKMQGC0m4kb
V8c6wqSQPDRigwEYwy5k+GTVBuYZxHECzXk6jMH3FLQ+54bbdiB/7vJMXvRdDSKEj7QMbkOOI0Oz
6WyDMqLagylJpuhjrbtzPzECLP8GELLQHvTBSHCACy1B9zInY5HKlgTY4A0tvJ860UJY9/R00dAZ
AuwCahlo9BjJwNW9WrNMR6eXoJics3C7IV/xEqpv26RreLas4aQaSrI5EyZLA8Tp4hX2JFNmg+fT
YtkVUSrE2f5T9SntH6G0NRWa6c5G3gb9VLzEYTjUNi5a5iSLvMgNSXAEPn6VlrCjfxTLaBFGvPxn
LZPSaHX2FJ+UhAblOOsPBp+C0bTdhWlsbBtNaIPSJATRWp6FP5/Qx/vGUzthE3W6bCjWbLOwjTiy
N2kQhqlOa2WFsjyia7OIEurpXiSuFNwF/iAEqZ7RXTiQwJSVYjTT0dkLPEHfDe5IsUZ3sUVcsNyA
cO4fkfjHKtAGcD/KRz2wOEiWlJ4RYMGTbLzDrIGrO7blBWEDCq2EjLi92DOk/CLIgIRQ9gqjFtu4
6eqVuokFLS+DJnsBZ+ZbVt41ySGUCu1jOPi1YWKJKZi/Ib7ua6V8AylJqxdSK3RohNYmURgtBIlZ
c/AWj9lKVUzwFubuozwooWXgSgcpddW2Laicf2JXRkPSDsqIQPCCAnHHhIohoEPNQJncpgHqPYLf
JN4rUXha32mlEhqAH/WiIqikVTfSbU5hdS4E2JPSf+ZZUYtK11BborXRctnOmuXHU9p58CnrT1bl
o5pKcsELymiHw+FDDVYSctBdBrdu6fEJ2KxB3sMMUYYI5NEJqB728x0NQ3tu/GlNbKIPH22l8a5P
t7JdaEXKrBNjwh59Ee/mRKOV63Gj9hjcMY1cBM/I0zya+vkmPBqC6aiXUgL5KZAPGQnCdg/4dtRk
SFCKhNY/iQTmU3tytr4Kc8H/tNIM60W544Upj0Kna4nO835H67baT2u1ImRsMx5DzcogFrxZuGmc
iypvYEH7c/OKOXmxXi55AENsVM3xCCPxWVJ4MvSQ3/MLoX0jS4Y8OWYiGKTOweBnppX1LS/pi4SK
+FqerSE8ZZrZGvYODqepy9fyQhIZ5pcpkgNCajuTQaLeSmlQjKLj6AU4wPqsXQi7FhD1QLF+wRTH
NdUT9vZMsI1V3mopgsqtG8dCduisIIL3W0VTgdd+tUcVaxSs3bLpKfcuWm72SdgH7YeBqnNqyqgB
SFCznJvYjgkvslycJF+71OpQ81sC6GdQMdJs/TAWmnXiIddRSazlK77b5ohJ1BPt4Sb16y8a52vR
g+KPU5a9ZP+N7dbYvxh/KLB/r3YIAPa748G9KWTMKiHmhfxYngIXUTLL7vIvC5fK/GgN/z4CHh9j
cWp2TcGF3Njmmabf1xqlGPc2UZ9LKefhpxJrGzqMzAdi0TuU9prEtBgE0/ofaBkWcuRYTm6d7PIb
oL2Fipo085Bh4g50BncqQ7RZoGZlUbTN6yxp01RoeCiWNMyC68YR+v+TBqkKKGO6mxAhgLVKdgiX
ghkNZt978E2diutTsMk1Ck95df7w0T8uamvKyuy5E4p5Wdu/OSC9piRaEih9v/Qu7WDqR/ktZyZB
p6VuK2xJ5d2y9Z8/UzjKKmKo1bNQVgFwrdMKRQaoLbIrs5Pbog+CPPl/Pev5eh4cYKJwZMNNAbzn
CrGmkogDdP/bf9EnnDaaeuPOgalb0uGZPplwnXHXSKHi1j7wN1jfp8unCyNGgH2Hoirl6RLRHb4N
NepZAE4on/W/TlUBfdyXYPDEfnHRKreXrmLrhM6tqjsZVHzcZlp8816xoYp9+7X27T1Gsq1pVJTv
tafUWBlFXhXrVUhXt3rThTshhMgKELY8f2wkNNWyVVXOajYhpKHoZsdOBF4BKeceuZoDvzxDxNsY
evrz7dFA4ZfTIjHtC45uiwyHNC45Nx6zDq/RkAMCqIhQLMYboGJwmcVeNB8KwRHQztZ5AeOt5sZ3
i9XLlRyEB8z4XQoOPCh3UPg9Ah0BP6YSjpR745qycqurk3AtJEhep4Co7cNkNamrFTw+wbEvHLED
X9SbCSSj5GGFP1dLY8/oUagAV2uL5W4HSyF3FfTYa+HX3NkpMOJLhpzgoDz4ubBru9I3JCUcVvct
pBKSg3kIduaQ+JkZw9Gu6NTR5MoO2/OCKiYOEW8jryKqJL950/ogKoCvlaHg78tLKCanP8FnEiGl
S/SeJn4ZUSmOFDJnI8a0EVsit6smMD4GklKzBFiffISpUAU1Jqvo0CU4/VsUTtMMx8oFO3RslLgb
VWI1w2QKWV0PDFiwjOCTvSSpODDxBauqUcEF05HqsyiZmoPUsUM5/udD2sDMbHo0bYNFCWYqdAYb
xeLuzqnOYhlSL5GrbwMyN8BX63a7UbDpqCPVXBkurlNXCc0pDA3PhczSEAzKb0wwccHmQkpJrvPK
r7/mUD2Egj0CvZ6QEFozGcBQt7AWjdYwEpUol8BBqsTRaFjzNCiull3milTxlE6zHwfBEL7WAjhM
elvtPS2lnaHPWHB3GLav6j1d/YDw8H45wUIdIpH7L75z8BG3kKoShkQOc4EYX4ch4ZAGcAKlHQRh
pXkzUC00M/rY5yrq1Tt4UkETArqP3ylqcoRxqqHIeCG5QYxkkk3jBVVHUTvHfN1piwifg9DapqzC
wIuveSlTGwGHLI1uUdKMJwSyfuMJctK9oc75g8XPX+XOtbNlo5ujtWkF717DhYNCppaWyhzCY9m5
e3WaCrseXcH9D2ZZ3MzO8temCy1M7kT2K0CIwnYtsXngRxxUAzpkDQoPj7FNZ6Lp4FAyHERhrq+6
cvsvHUHTjgAbu/g3aQYTw4UARepDKjb7eQZXwfdmEiFMSKq/JLGosjLIofmKWGAIINkhgg68unjW
FY6UI3K1U8EoU93vVO2ttr0m4BM5hGgmDaOvbmUQ/K8O8VTcnxD2XNSkvAcEga5maPMIN8F97KfA
AMJGQP4dAwc1PD5feTlp3bjwiwtktR8ijN46A5Q64BaYmwB6KyoL563SA2yLq5QootEvCU54hX0L
Z0H8TdUk3eK+T8yX6rGx8ax0UXcU/6DY/wrtsoqtebEugDTNdjlNjyTXKD/FU3S15Rv0Cv9dc3Ri
Zh1sV/lY7xBR2fM1Di2xHCji0AxH/6uoTp0vVkhDaOJE4y2xQ9vl/1Mc5lTkYXV6+I+VaOlyGCBg
HWDHMlP9l61gu1OYmGabMUScUYkrpDW8QTQCRTY1KERnvMqUpTHJTpRjbdWPrtttJIK0NSBApUMY
+gx7RVKdvn7JgrzY76WIZH/F5zoNH9o5cGWhBuHu/RKCd5KQ0cUBhew8MpwjN9MF+Hb6wCpnhfzh
KsE5V8gxEKgxRsKXV/WAcS13wZ08b3i0kxo0kuLADHAaQRUhyCfiAg1zYC2ARoYkw1z0/9R0l9bZ
5At3cvdUWga4dQqz7WrQbFxGYucdYrgbLUnjyrlrFqklHylqOj2uXDZL8kq9UaudabvvB8WoKLBG
N7EsD5bn4aSOtKpBItRGTdZ/NJlEDV7/8ZFrbZ9JF78AIuNB8ZskqECEfUfuJ508WqhLwbHMTO1C
GulzpQ1G2RF78gEP8eY6hFGYaj30ob1ResEgdWQMuw124WklcpvxNMZ8jPK6SS/8sf8fKiTvbQHa
sQUV4wNqKVykyDEGN08rQ4o6GyHEJ9P74lwDgAmqkfqIdYIEYXytkzWo0oWFd2CDMIRP1DcQTI4f
saIU85RlH2RJrn3Ze4+SeYmJOQdH9me4qv3Em70rn7mSQsR7/JxTIg3TCNfhMUZCepTvGj+HwH+g
tv8ZpzqR7lOsSfRoUxWHcKPSG1jd9agy2OXN8aQeWX6YQT011bYEK02/Ke+adceH60V9xoqbm2n1
zhskUVyglpGGXoFA2i5ERjFNuH44cUF1ufwNMPqUmYGrJCNj0ZuCEmaU24I/gRBtnc0tWan8dMSA
SLLXztMHaoOzYtBXb2SzUgG36Mpx79y++g8Rsa6QVsO23b0i4S3IwEdm7INsK9YYIE72w9VoNVyT
+476k0gbh2VpON/4GEXbQTfiJsFMOcTogyBu/jkz8HceRkb7fJ8ph9ME0oW1J3g51YIuTx2rhkvO
CcM4ym0tnIqm44LSeV2BRa99xaocz65nY4VlQMUYWuw1Buv0A72Spo0kPFIDUqdUldOdwBdITt5t
moObXe0TbfzTZGojRX7TAMKdZ6dDnjhfO7W7sT2dWtXkrrvOGqJ75XU1sG3u1x8gjzYAkgbeSBgX
VtOHsjwNNRB/UiEc8ojVbguwzUrWgINiXrKQtgSZouN+hipkCAxHSabFsK/TZvs4azYjhxk1jtn8
F253s3GNnT/M7jbWxGNNxR0sCoLpNQ23CgJuEPe64E3pu08wuftzADhpW2SFWF7tzZ/JczC31Smc
5OFjfs6PAvRm4C//K6TWUH8i3fa2uK1cQpOB2mmscHCwtKJg3wfw81lB3OqrsZ4sVe0W2SkB4wS4
AO6B1FUTZUXAiHTZSsOVg9W60h9vO/Ish/YfNev9xV+KWUmPMIqWiPVRZkJrqbDxIY4f+hy6sGyC
zwuugcso/GM0fxIzOrVvSTLnGFO7935TcPdgJN5f4xDe9pgubwiq16VccTmOyWLdBOj1bO72ga0X
XhPYzAuf1sl3Ir0fQqYc/4AW0mbJSYWz3rKjCeRmiCsah5qlDoWDoKLfIlaUNrJmbArHx7VFz2GS
OehgzjqbFtcVXYAgivwPQRSytIooL4/h+K4i/O2fYT4MFSJrtJ0+CQFmk6WyF7P4CUCgkObTrK/P
vjXkoOP0RwfQJSL51MZb35hv8v+uIZusvijpAbJGFYvHu5iK0BJrRMg5o7bOAixNSFC6c7PiHfRa
uIAhSToKRZyUQL2N4mjLxGdJoKRA2ohWVWUURwg7XSrHRhQnK48SDv51FgkDpnwjhwWupH+tHukr
6kdEcrVGr4mk2IvNxSZ66i3MUdSbO4rHxyrFV8gA7RxYx9MJAc8xqp0mrvoZKiq4zlFW8jQCDg0k
jY7W6OevGhT7a/HrQY2nuoC+x3gvoguo6aW61OalYTSkZJRhs3E+bUhLLZZDvnttnJmFr8dU4SuX
PTmoRba2OzX9fu6le4WUatewA8BKvwXtB7m+PwtNpA6Ya2rBhkKe/7lz2glc5IUrmZ3s6lUh7K3z
+aLDiDeUPpy1n9ZAfqJUH1B6m3D5H+2EpBPR0h4b6Vadptse3XEGuo0RgA8IN2IrrlSsprUN+nQg
GhzcsKRw5FlEtf/lrO16gBw1+7XekRzQp+xxfhW2NLTBX4194VAkij9a6PvzeYcH/f/BPgOoojr9
HoeMcT1sxPpJabd8GcVOYTejx2MAqRetDXYi4R0cbUn6dIkcMm/nDGBOa0jl5N9GmXcyT7MbITnA
4exPhuNgFcNrcFvsoIpsXuHG13DXIFSF2PcT9fYMkp0OlRAXYMKEzMkMa4nvENotHISW+yOHmtc/
sWJQFeoVvbHckMObpDN0IJ81F5jym/g+Ubj526lSePM8LKxCFODAawTaN2IZvd83RSJ1wb6zmKcN
WcvGujUou6khlYrRHNxkz+4TVi+Z1+MAZKEVpib7b3/ouq+Pf2TDLneV4QpWadYWEL1mHF5UxxL8
MRyENejRl+Fa7N6mSivNqXzJj6tJAYpwFKZuh7Iw97pZzfQORqH3WJMs8Qkmk9YQUVyp2OvQLSve
jNMNCPLaHPgGMViAZLsM5J6VDKeyJb/CVC8qT8pZdLgezYygDouUHS9kmaFzAn9BEzxcmhYALgrN
o5iO1PfdXoU+HtcwPccV/y7Vw450v1BET7ZZ7CnH8B6XpL6L1Mut/DzLDXcfEdDZfvoUkcXkiS/K
C/Vibuhs24dhlQARj1x5EI60uoUTNDGMcUcR5g4NNr4TkcDPa6A2epEFZPYB9YnctnXAsfxupPdx
ngoFEKMoZuQLy7KgkLp+0QeykUBJSOLzTWM+q17liMmJG21Y1e4uStK1Ydly9vUuajthuFM08iH+
YzAdK/l2qs/opoR40OF/DwUq/dnGn0z2/ilux8/M4dcj4krG4u7/lnn7lEOq0IrbBc4O/5hHSy1T
Wpepsn0qAx/zn+RUP5lspq4Yu66+BkgIzTdmaz6Z/3AnDgZGb7BD5a59dT56mCx5q7tpV6e1g0kB
qlp/t145199yDIL3SIWy2IsbAg6vE+FMUMiDkQe7E51wVnDFzGIVDt5uFQu0W91BccX6pXWWzJu2
IOwX/R6Ipi7Rf4OlkRKgZdwzX+0As1jBxqhZN4aaNx9ypn7OBKU7yWvu0xIQJ79ti6gfT5KkGRj1
j5oUhHhSJZ5NjzYmeeZxOPo1AgObdhAhDA4xAHEjfrUSlV3qy2xri8d9yZp5LNflYLI5HlQenVuj
xT7kkN8pKIKgfGjpHDhVTPX5m4/WUdFByqfT0o0VDIPBrEXEXa7/3QJFPw4ppA+xDGkZThxQp/q+
cRaNvKN4EEue2V2TCgvriV/02coCbkV7a8qTbV1bnefaYAQ0mmrsY5cAjjSg4yrMhEIl8kQGasTN
bfMiLHz89aTJhReosaCYTLxeoFnOxP8OwahvPBu3utvYLxVAuKxMpfxODbLYt57VgaNpXiBeLfsk
HADhsHxaYXvt/uTz9Ul8ZT9SFpDhzHYVOTPeysKPPjFmdSG8WhLQuGd+j7gx2cQXC9PXGi9+NtFU
U3oysQFpDEgghfCdD+2mu0whT0NROdR/haPgxQO10IWTbVK3k0LBehcinwRK10daNzRLexQkA0rl
VngOiz+KpEE7pHMGd3W4SAkXJFK6irLZguXCQw3YjttnkY2VlBKUZ6lZ+OBs/Gphqxdh2Cp+TwaT
tCyvvLFDLD3thnHp6M7MfMMaC0KiFa6BY7t37UVji5TDBUYPcPVgyXFVBwKmqGy96k7tMYIpjnJ5
tdVgv24rvvmKEiKSHk3wNPpNOmO6hTSJUc+RYpSUHZ4rK6apVqR0xbPU5HKq1Ploz2MIgNSLQIwZ
dda5647wIjew/OpKC06z+A2U5CqaxXV8dPiD3lBFY5chktXjgGSKJOiNhCIttw+VPQqK+3JZODbC
KgHa/yduv8z2vNnvTbhpXa1BX1hY3+Dic02ucwEmLUFI77YTCiKUAX7GcVfQWKi0fm5kfJU5zAL+
HzNf7IfiSeJtN/wfeDXrOi2mo/DRP0hyhQfIUo8OVJTFkDmfPxW7jvJ7Ev2LTHWZLkQcxUP3jp21
gioXCzlzGonB4LOHOyTgqZ8HqriuNqI+MyfwX/gwfvG41wqic+Cq8jKF+RRl0BDXTtHBUWazv/sY
4tot7zUOAGLpvJWAhnXu9jH4hACwmqZ4V1VzgXfx8O/d1wBvmjOwWUS98xYllzcpIjK8Jaiazay/
lsb/dpMQb4bYYXJhJ6wsmXjZZtT8NxZuhMc+gRKSwoXS0KghxsXSN3ekOTtZ0tnuCoh9oReO0aDM
3l3bM5bEwWKBvrfLOIDHieXr+POeaXTJ9pUqpVci4XjrIKqmWt4aZH2IIRupuqNiYwqSE4PiFjbb
X/MNe6QT8ch/uZTiq4Z2SfqAVO2Y7qyOrPNZNdRgmIIeAQpsTapSuUQLam5whtDNGVRy2ZLvI7Rm
cZB6DUyE6899onMfqUTBXfKhThWKIsymffrhadHWlj+NnUQPYzeBxu79hIrRymQIyuHGImfbwZ+8
6KOm6gyKPNwHUdaQrS8zzx1Jv1+yJBhsAvQBLy3+ebAOHjd3MXU4yon73S9DwMsBboPxdccsConq
4kDo9fNXSXbFJij3KI81gRNUTY0IjDXWolF3BuhLNS5+Fr6+OCG9trWLrHE/aABN6ecjMJufuG0y
MzbGQLuAstFKsI/j5caSSZkbz4ARWMplhuujcTlwg4Ab6t69+ynOxo7B13N0KDua2BGLWF5hI2BI
b+vN6+UdJxO+v9ExavE7VYZQt334RvZktHZO9uFiWt4MQVDhGiT8w23BpWMcfqwcruiVW+caaRqH
R99UYgd7wydbXVZXIN7OmLsBi8mCB8fMMYw55sDRT2gXdZTbFGYguJVtX5Xrq5yvuUZ/SwSrYSws
quK1B6SyNOsZ8rbu6yXqNf6xmHadIgXtLbtXjatzJz3wlVGuxM+4qOiiNebTKX0A5x99WaR4EDsd
d9f2AnFmlhN7pJGsuYrjgzB0UaFbglLtpul3rArt0gu8mTDOsC8tHnNFCQ9JLH9mj2MnRqHH8idJ
phQeb2dyq0lFm6bZkBioAneS2LG5bUbVa+aBzHBmWNA/SGgVHBAZjvb1R3VvLUULIeqeacYMNpvW
qvrIvmc/FfNotWHrfxqqICDsfhp5mCb8S+RvMgqkesaRFT3g0QVV/v/pwgdjxS8KXREJ3Qi27Jek
YZhBTIU4tgyTEy8Jr73s/AJj16+45yf2hk9YnE4+SCtIf0hSDMjrxvmEfBr+AlBD6aCyVwHvyBVI
RPjFJnJMCtf9rtxkpOvP2rklMftRP8ycvpK1z+mAVfGqM7GV+7HSpHwz+SAVUiFHiQZF3uMqzx6R
eSxT2uF8cV85t8vTTBtWRSOIjxxmxaU8F7wCq9yB8K9/4AmISuSz5LlawJQhdOUFRSE0VIowFOYX
yv9dU9vC1WzeTe32IX3+pb2W88oiCdrbJB3yzZZhBfx89YKW0t0wRta2RSqamPBnK9xEUXW+XKDR
WnYTkFweMoE+6BYL3KPTIfr4sMjiNvpszknx6gFTgduzjIMDgH5XGqrDXrll+AsZmQO+U0PAMdNJ
xRdp1XjVGP5lmtg2Uau4FuwJ53pMh6t6wbFdx6te4SxzL+NRrgPRrTAKSazFeSbppb7nHq0vz8A+
vlNLcSEfy4tCtnD/7sh/ziPhE4fn2DgK2Hotb3BbYer9T/54Qo4pAjQJJ5xxfS2vaEvNk6DvvGA0
OYimshKFGf5ZDGDhq7pMBRIxh93Q3fqPjgimHknVsI9JbC4c+jLIhGBpCIypxzcsXn8xL3kFgfSn
OUvpZ9553NOA3oxa9dABSmZy/S+vFCittTlpjS4xkKhg9KJK6iaX8+HbE6DC1qFmpv3wQWymzuv3
83WI5+8Jw5M6Wum2uZpRkyowq0OxwQqpu3x9cOreR6fFiAve/+Hz72v98bc0jmuFj+bLiQtp4LmX
NVf9rbb8Dk7W5IZ9FkfAQWbeoYK7N6XgWCDqcLzWOym3jknoYwucsV9JRRbmxmpKQhpWzQMPVIO8
K62uknJuYg0tf0QgRViaHhl0jlv4pCYb6Fe7UlcThLwdPIqDGYCCdIMBcnvHwCXqsmoqat8R6ud+
oNUiLKe9zkA6rIAfvhN6Frz4kdKcT+Vb4QZcRDLiPoPETZveD/Uyl+0PTWbUezLIkGP5qdngerc1
Z7mRaYmgXtyo2ySlWjGH1u/kkrStOeWlGOGJnfDai24siVp7YnFGhE/rdi3bqPQRxsjqGPWeSzA8
whyohUZCvlKqsip83cM6Qq8Uz2s2nZZllwON/GjTOJ+D2hsJIA44XT1j9HmV3BWsRPRxpqgmTPsm
mVOtSeKauBlWjfzXHM7xyATQGXz/jColsY76ZazLbODDt+3FQbsrDxLHTNEdzHXDpzJE8Zq1XtB1
h2zgGdmGOsavHizY59rZmLdRcYOVCg/DfLOZVxYpgcceluq0uSeL2QCFKOtRKBlAySpkES1wq42E
vMuWN/cBhEzYDuae7o1crGP2FPd05UxuibSKbbY/i4TQJu4kBZW5l8cEeLTEqCeevryJetYetRj7
J73aDBzkAESWwKaRUm9tcSqywK29b3HoOm1HsmXhZvOE6LRd98xvXU9VsqYDytcPy11ni1dkWEjD
zK1ZcHlpkwwGmnB11+YAXaRzctNiasBy8VxSuG1CPaMkEWhPRewQWRVUKRKwpz/DAkvkstgeSEHz
9Yeak7ghXneYQHEqbnaCQVwJZWolbCNfKN2i5CGbdZpV/yvbTybWads6Vtusnr+w65+3d3/Sf34k
+aMNiBzEDiiNSNblR+OdRu611R8AHz8p+dzuadi7/A+1LMTHnF9NRKnYTwI/QFXDlglg2bS2ukCl
ejaLEIz4svGaKQDlVEfjkW8dZfLcpXy8TmwH/S0GweQme7UGWLxBxqgB8G0SjyDKkSvSNKelUDTg
BWjXiGZVeNfZ+wNc8fYD5USfvpWHBlVtSQi0cbrRp7Uk1V/THfhlicvPB7kjDwd+PonhRxSBNzoM
KVPH3XfJ/rsTakdvP0ANsXYZAN/8SJcm5S7G9LQFrPV+tEEp2KYkW2nN3hmY/0mWasFHJShNpYrj
0wGD2HTCTAXQyt8P/ncyAOCC9Qnc/TE4/lGuiq61CV9DIwR8E15hepqRkgW/cNJbqzV8POwS4I2+
zzFjzjorcjxCGe+QaxH2v3uVGtB/2VCtXie+XdlV/AucvM+1cZkNuBCMiG5ZTpXEQGNDl/MHrSmI
dXjCYL3wZAR9/yqRtk6ci71LMXfPXneIwtIi29J8Td92CzWqjx0qRJXRgS3B9muSKMRVr/09Girz
V7ilVlFN4kdOYseMyGX+2vAGGkiQGHtI49Q9TXRwUElryIjeKbwkywY3Bl++kXHS/OnAjCKZtB/3
G8Rtq0rrxqVCwH6xdIs861NDVaO2gvUBliV0af0sHn6Kq3b7neDfbT8nnKQlsNwguFFwB6F22MNR
0khEdzWiVyvO8H6ydPyiEm/C0djUn+XDbrMZdQKEclfJMxtS5dZfTiK5ydh5taFUl3lERaiu7x9X
dEQApROdRK28BI0Jpeqf37ZImvwfY0YbGxnzV0F9K++7lxXq9ZcwwyATvdmHe7894jg+8insBH3G
M9K1vhTeZWJgYRrK6qA3DS+B29LL8frv0noj+qgtbOUj8KXpTeArN6i/jhp6NRR0+egtdf6m0glS
mutF7UD1ztJ9MMh0Tui62l1c++pAU9ZaoOeHUsnq4ogUtPGXRChY0YMwezKxsSUFsD9qkCZF3vWi
2K6MJMSifpc2Gby9vYxITmqZ7OCVa+BeZCaIBVkhPiy4tJiLyKvlZ2KggXdSrpwQFRrmqLiCBJw8
KoGuoTAmquqya/9GcvGo01BonZaMGGbDVgfGdTz/w1Yf8JFuP/ag3071vhmkMkZvjjDsHJ6eWm+M
2CWfkvqIbzAIGOxyM9WhHPq2uhxUPLkAiA6+0hs2Z2cCW0b8LERdIFhnng3nKNqOCIkpvVC78hnI
mnzJ124ocIWhOjRr7ba4C+Px1GFlaFF7H6KdY4H7+e/rhnlLkk874tJ/4FNR+Xe63Aa7B+rEEcuw
YKyerNMg4NJDPiEev6z1HTsPi4lpzmhBjvMJULOR3cdK+pXv3mGW4PG/G53Ny2K0f12fqyV6m90Y
K3EIwM7atJVNPj32L28BNqGyCHf9pPhuyz9UiQMVUzDm1Eq59VI5BaHy4VJPCvpvnivrX/d6hyAs
lKfGWoPUG/33Z4gp9VsVOZjaG0Jn9XMPjLZCP5mDd4PYU+WazMH2yyVNZYqC1NbbHqE1mwIyBioo
DvBDV6VI7toovYdFHjOzATuthYIlA34172p2+iI3scSYfrqkvjKHKLmJgCbQkwYOUken4XkMnNQO
ytCNbJpRU3CqctRn/4woVyvEMPOi+QQJ92UUWBPBxWz6GtleSxvR/vrrM9LgPuJVLuJgj8n7c/6+
35eJIxwsT0ttCbsXi+DHblGyC0fUOzXmN9KFJJNpCq1i/fLlJ3hzAnqCpfns6Q+Hilitq7U4NLfQ
ZMrY24kI/H7ibvps80Lo8GqaMX8Q2P+pBJkx5gUeye3mNFVudiYvP671l+JPdARWtGsUsArokMcG
AboG5V4l3A0UhOk6bSg91g8y+GBulvySRzqBTYiIsMYAUwLKFUMFGpH3ROCaEZa211w8wjFINWsW
YcTRsxISkFyH7WwyBigi2fA3Fk3TnHywJSw69Bt7aYYAmvvmiKh9rNfWsXzraHBCrwHccWwtGJBj
+ZN8NMMbTc0Kd4FOJNTf/7DWmsZOgekuI5SFTbZXyq4IeJADIxHC3JD0LGnqgpnXjU9RGeqwFKqE
LsutlmhmAXPVn+9yfZDavJBz7UTVTF6o07//BX37ZxrBsLmUu0MCxNc1Gt9tbz8UqYZHXkRJqYFE
pfKPO7Y/mu260DmVTQYutQbpoc3Zv09PrOif/ihCXIGWT76hszPuFN3b0Bi9IIKHh6RGxLeViOo5
DRkmCONV9B9lNs9V0p1ChG5CaHVc5bLiHXlTYF/7VLdDefRXaa5anNw5D3yoU+9hFuCwGm8D3Q7g
2UvO/AaxyIt/tbkgil59TUiIaCkiJvNd2eTaeyj7nAoGZD5I6Yit66TfQMd3WMHU9AymYh1CcaVo
YoxoyR9mpaz4jVF7JxADtT42RgdOieUgYJfsKXVaeLbcfG/J84mtA4ISd/CQ5riKMM6p/b71L0C+
w0TDEgwSqER6JDJVCzrrKdmG9UTcsOBo9qYtpKVoE1SU3tSEEqYBqxOWIuPvHIkzRbytvTWcQI19
7+6Ib41rndWFaf4b1aV90nXlegLJrIzj+iYQCWhO/3BE6AssqsaSG6mTHMfIOyf6GvJstbA7prBg
sG78kkI/DoQKSAftaWkSOxYDgof6ky4838VAbGSjoQg4aWjHECuuOgogUacaITGBjRDI8QM8lxVM
cKKIZhrru9udvZ/2Vk+f1q/Trwi162YRr5D/HbJr/OajvOKvUg5Tf0uM6TE+PHHWpCdib1Yb5501
3CcvDlAqc6NGhXs/rvcC9JGvG1erzwjojGeVfduvQ8vgDRKamzAhsZ1Z+Ac8DVmFNGtiqJiU1pxf
x+f0Disf+MCkXS/pkSZnh1Fk3TP5uawOxVy8CjO+/giggeweHJT4YKDY7njxlQBBivyBXeMx56PF
+jLc/mcpPYaHtkNSnrAQEoFNyV+HRNrPyoxCF6SHopjWad9vUzKj1frcyLR2EXeur0hXvFm9wD9o
Ce1gY9/eqDaFMRugRXanBSSx9niQKtrxuUPrtcAxQFpOYvfxlKTDKxF1eAByCPRvb3WFggfpcXsT
c5EKhL2bDQljyDeYwtaWiWGUGm8s1MNP6gELFsImorGL79uD8rCSLJyM/HSR9bwNyruNAOIlLKuz
N4eaM9Ga4oXvLrq0QxI28Dy4pYV9nmrk4suUj7EVm3nXx77MroQdAj5vGFoAGHOF0pa9Bdk3xBV3
mWHu/b0oZcAYfVjB5akyEmF4qLRcNaW/b+wrkXMk5gG4FpLJWyhuqHoUqbi1yGM717Y1XN/geOXp
tsSr4ZEDf5+jHlqXItO4XyB5bQ8bJ0tPeL+Z/3K+F5jArblQLDGIUdcj+5no4Uxq025S4gVY8dba
vWWyVQlC1j/Xe1aWHiqvFW4ztq6r0uXj/TKdSqGyzgR/mEjPzI1QljK6+bT/efE62D+lOygNPAgj
YDKnA5P8DedXUCvoI5FlF4/QuCAZsXBYOvSw4j8/rkVH3ptNjzn8sZzI1dpmL1sRi/t7t83jedau
E+z48khyYWcOvxicarLI87hkY9d4PMYOiLVaJmnmFcjAbrnbGNSaRB9Tgk4QMBUP78ms3ERTBCM7
tMxPdEzann1daTo9W58hW0e8uPJY10na/QEcE0pyyq0MrUB6MOixhWq1RCqOUXW0ucUCKd7T8/Kj
zd5EoB/1ToPFvYhkySsL6/GzrhMiR6tLjrJpMch3JisD42GWuWIImqhLLrWqDKtCxaiBvvOIJ+m+
vRexp4QuI6AjlvMOykiHGim7flFM4MXxbZbzUW4aeDPQLpLswhwJLx9kkPx36V5uOj1d7PU/0UxK
kAFiy6enRz8ncbOtGtvRBXtIjmSh+pkdlAs/ZS2EfEJx+zgYOR0CJZ9JiIkAEzIi04zu9chHjxzJ
MgAMk8j3Hc8iabIec106O+o+dfw+F68lMZ8VhK19PnTbNNQTBs9kGCKQYstjB86gkUvSk3YafMls
Om+u/iHJOUKLT+Z+o52DWo4h46jVGzLb4nlQZWjNJnPWUlNGMvIi2CCYvSSmpotew1rgNQf5fyvP
U5N+qauiq4+U04chjXL1E8j09agrml9lHx8UTF0QS0WrUjwZHnaPRzhrNCMuwuzQ+jLPDOqR70mv
QBoyjHf/pRBbWYiybsG6zw0A7Bf+tux/AC8d/aR+bzXJeRxYYqCPopu4tFmETccZjVAajV1Ia+57
sSXsrZjX8AiU+J5INT4DPZUpDQt287bOFKiZLuY4amn17VsSy43OyLppgYqqD9PFCdNITPVTfDzt
RDjP50ir03X+2IiBP0EZYba06/ZLvH9/l7Aw+sjyLuNMhcTtSGNx/hEY/KkpEA+P8nrNmcisXK0J
UOzywx187MQPTQUmFu6vMdpG+QWCJiGy8RUD+2LT8smNxX73izZCTNUzwNI2PmvrJ/aZwJpKT6QB
/Il+xr6LZJ9fygRTxYkydl9ZIHYpNdZymoNXmC2z8rigRgA/NIwu05qhSTH6+xEXyMalKj5FSUMs
6M1uI1Xivl2uyROIxgtpyXKurJXc92gu26vqfOZ5b4Qmm9HN+QWjgFcskOb1eFWzgcgIP5fZaMam
RgZX03DOFRvlSiDFbLijAOCYa6xIsmQKLWmTe7kLQ4qJNUlSY4N31YTUdaw6LDp8U5wg5Hy06ev8
3zXQqwX3ksOSZfjr7lfsBbJYJ01qMu/Tbg1bzFmqJUABAUqhBgWABv+ZomoW81ZTDX/Z9o3CFhxz
VRBhH3Eur8Cn2mHbeXIFOI8Bf+BuRmBUF0gz38zMtg8P6WaDKTQeTPr6QRetul4YugxtlxrZGXE2
C9NQXdyNnJH7mO9wHVy/aHC7T1p7fpwmnr3C/1OhuuxaTTmdhR+ztjim7GT90PbElhqWp0AdQ7ys
ZeR5vEQpXOklkpRbWdKV+p9wV9TxEYmhSFM2FKMiIFDi4GU+TTFgPLctythT0Iy1QQpn+fXJSHUo
V6N8Vn/y3KKUoBmayI7wqH7a9TIlZ93iLRWxf+hxDwVPNAB1FwXI3m1Hm18xZoEckLKNqJ0roaMt
sOtle8bAf51ZVnZQFQzDNiHE2zkF2+4RyT4LW3bWbPVRx1zk4cj51AKNW3dgoW+U0s+83EPGpoC8
ikZ/fMpG7wnAS9oxPu5gjsFpVYvPfn+sYsndOxYU/2FD/hUOsTxJ/syB81UupazumOADmWsxbnzH
dGpelaU4G5y69ShZOwNYGYsNvp4FmW7wn8zKpBwgtcPRjATMS3Dv4NX/cjgMYXZds2IMP9tfICaB
ztNWYjBoveomw8f6y9HnJKUt6AETHsVvbVL3wPQx3ooDGLJ4Q7vLROyHcR1pU1N4QmPnuX3Q/j6c
jitxvA8arWiRtaOX5O8cy2ipfsh/Tx6ea7tsF0sP9Kbh9vPRN5RZrtgDQ5JZi+eqvL/hSDahaLuW
Kt7oCQeu7B4hzeLOw4uA8MILwxfdHJzE0/RY5Rpd/uE2BltgOcbGX9FbA39JTdiIIysWNTcISWwR
RPwfr4yAtwDnxw7oQMmsR3DyE5dhFH/sWcUGIDBBTRUgtbeHKiWO0HCfPIECdR8ViotTcyFG69YE
Xoi1buXYIQrEkgHOikhTWELmj0vdRPN5wFa92UKZVH/rZ6E46aRvxVmVW462cHee20tg8F2VVnhs
yFcsi8Xal7JdkoCxFh7tGcHzFvITs5w12OtLjZOGjL2Xnq6N68JSlP3oBsi7+iJfWRugUqWyvSqD
PunT4CBqoiGmRNX3ftj8AUwppfyR6TpxRCRfLbGmZ5fDCO5O9YdkI4VFbyHo6jwir6a3tX0EWz7S
0zDWXpOQ/GqWZwJesA2NDfDkLGnHOdApi3lxKUY9yKr5bxMKkLsmo7UrJfJ62/4v9ZBDz7yIq4xM
+9fXEeAm9Q22W8BXei7zKMR0V0NVqnnjO1BdZIdSSrahp/KWQr2Q2AkQZR60TchsXvZ/vrp849/y
2iESI4y5kssUH9qQdMKMXF/M1QdN2pB1T371gypwL9FKgj/5CHP1WnOCqWh5yPXsIVOeBiukIW60
I0CHThGptksRbzkDWBgQ/vt1R1k3GxR+amVN1/7A3y4Y2+lMKkidHrV8wyCHG37d18EW4VRQOrXh
Whz/FecztM+DuxRrRDyeO0BGo9jXNigIe0vsosvucnoaKL64Y97RGH++M7tHUs/udptakfwONIMv
hAx1MxdUWt6qquDIboisxZZA0DjvkPfZxR2rf1lihK81fICT5+UHNYeO4fA7fzMRhnguXB3ZKSfb
ijNelqGR5hHtBREsbZYHRglIIeUGdDjS6NzW5+ydbhp2yg/zB/pIj4qARoHjS3hfvedfqVWxjxGm
rpoWxem+biNvTjlDnTp2piZztoytknkSJMveKT6RdrD/zwhEltUFpK/Tf4alo9drw/O3PTyWWD5M
PHgWPLYYiqxaKyTToRrIGf144hS3n8TNZD0EQCsk8iYuEunfqQtT706vztpSGMYSmGP5Wb9ujt6z
sbxGzju2yUHn1EXy4DZKohWU5IHNhIBa+i3HwYqz9FPuuslUpObm58fdgo3t9uWysk0AXjASafol
ESQUs3qrNYQSD0KRSomlyuRfQqckpHYHQsSG4rri1XQimRG3uTCZGS9MY2lZJm6p1orBUSS/zDkY
+aLdjoDd3i/67LwTh5aIPOoHpU1NYiXUWUnhqVG9EIuPe53DGW0eveTy52WHmziGEgfcfT6KOFhA
kJwQGA8T+ppeBJMPpSifaAImuOmLeSJvjNm3FuivyVUNsdt3wPGzq2j6GHlRH4PLHm3VNYwJZ/g3
FcqlS7GYmsYKoHEx5yQPV1YxRzcyqZ/JT/WRK7s232BBKvQAMCMn6kRkvqrh8vwus+Ld6e8CAT5u
Pce/oujbZ9GpRTDZjCeLHXM5TfQrB+JP8O+1TMpwnC2N4F3rKxhp8yqxRdGsNHjbcbIiTlnocRGF
X3jg0dpwA21KngD/qtanREYwyEazAxMDG1PvkomPtqHQ9UFEZf2+OMkYCaSzBngBzhFsN3A1pxyL
lje8ukIJHnh+G+9FyOgJjT9yJeW7oQv7BhIGV03SBRC9QLjF9Zmq1p8cxA6TUeCfbXHnikbE9ChV
wFkujgCB+FqXN6HrMM8tUVckzfEDCaxRYyYMEg+9oD6+srdCk865m8tcGSu08v8Akj3EwPnzSng4
Cx2s8Qs1ErqOZoKEP3lbY8rRWTM5fMCvXpD5DNO84KbcZutAa/aUxPdR9u6YiYHw35Xz0h7Twb9Q
CcFH8tipdRsUVnbCsWSBgMFdIXfsDp1OEi+l8DKUCgzxj0tLJPOfqzcE70I6aRaRFQPJYz9XPykn
G+pB1mjaf4dLnwW6f8kMHjSS1IldjJ+yqt8fM5UQ4lrQGl0GQTe4swbZkzWBiFdeLBtEx0ESnepu
WKI4INPAm8LRwKxWz0HqRdCqtvFocvjeUoEtH7caW83Xsud7EoNjGBOTsMAtOATpBPTz2MHgnAuF
ZsptmDZy7LXt8FdeEX21AoL2KRLf4uicSUdfX7fIYor0uNa6oWLicSyvzvKZbTLfP7fDcgDz2oFv
dxR/QngxAq/MgA4XQO4w8b52P+oeylZZYPUU8ruIWveHnwzP33zcBkhIzjZJV9VbDzF5Wk05khAt
g8K0Bn5FzoCm1mZWRcrjY8hobdNUdnYFSccMsd5Uyj0WLvWftHh9kQybbidUW4bTsa8LsjkJBuWW
czsGAvHG3Z3KYwiH18xJplCFKVVA+/0pVEbkFHmpzOO61twnp4tYNv2HQLc4Q9a08ynVxPuH946l
5bSrrg8y+sFjlQAhBur0e49eWosKSI8joiFMiCPQhsQ8kuouvFjvseZK7KjGIlVEiY9/X2p01Q9w
2FlUt7SVFfpPhqzjB7YKg8A+yXpjpue/V4Zohjxin6qPdXzPnzhCrXjtf83KcJCEABxrackUi2/2
1CeyxxQKEoPX15ONmzo51xrYNnQF7XPINRUuV3V5HHZSrWDmSZcuhKUGFpuYI/i62Gayx0Fxko8N
u+GahadOYCo87fKevzdcTdwFOgrcPZh3Y9s2wPK3zxOilYSI9tmUD+ny0P0p8QjWp+qtR0n9p1Qb
Ejb+pIV/CkPfpg0DxSHo8jAFbCrqZibg2a6qTV2F73W5SpWHPC814le5naF3GvefSRKW9YCIVTn0
zik8cMIpDU/FPhFlFlEuyS63alVXkKEFjCZnPvE+AYtYuD+pGnUjzSzGbqRt3racjzAPTf988n9D
gfWWZnCiYWoFRti33gysl+5Q/DgKlP6YIIFKt2SGPiByzLQNerIxDqJFWuDJN5gMbBmvX6PwJyza
nO97MKrzJDPMvjuJFZ/Gzv2PE/7Flxtxd2ifZzBKSsYcpS0xh9t37N6IYhT/jajbqPlEWJzlQ3ze
ovPXXkfAmwMnb++++DrvB0jn+u8POmPP8fOyWPtQ8LrWUc9aP6pC4gU+0UVehFm7I/XsvQaiHrRx
Q2vNf6mEvvi1obzUj7BpCUhJGuEgUdH+/rOk2JtwXYlyKXk/5MQY74Hw34HzVo8duPI4Q+2Nj0e0
8zfrPgmU/tTpQ6lmi0LpBPOU8cF1YMFGEjhMjWSVmNqT3Fri/2UPTkkt2TRUDpYsrfJ4KU7sipQz
8IY3jfkgooKqxiKEFjQnJws1FIqEaTF0cF+VWqB+qBc+k1inqP3nTPGjwdlJ7EnUMot3uJMTZR9S
z2vx/m0lXkChmWlDgmz8h9kIx1QWgAQoDxcjoPUIagc0FrfrA8s5HfAIvKukgselQKZ22rSxoaAB
VMKOYGBRSMsRV0jioZAOux4FSq9RgKAfD9uY3OVX6Bc298O3GC/bd4yv2gqL97i+sd9+q4Cxi007
uiGSs26jJq9lv9LDRGBGWpPdtcAriOc1ia8LUIcpgTOHhCbqe6KFnH4usQLNdhtbxZ2R51CHG5Bx
y2Kp3k2Qi1KnbctC/MCOgMb4gsno1qRW0ZdAFs73vI/pWBnnlf4TbPUgW7kA2fG+rBKREDxDekFB
uV/cA2bWbUtJ82DoLA6lYFZiHtsZRDQnGlxm0KiMILecYQlFtgRye2ipyEkii8/gGNsrQRx3SlAG
efbalwFzIWKObH7EKjBuiFZY7THVX+D/fWaf9Tn4QvbTw/MxW3thoBi4/WXEHVbY7OfiSDvuh67i
xlq8DykuFClPvvXzOb8JUfEsFOkswpczNiYSk2MMJP5KKd7KfBdurUUBgg0mgpgyOpWdLnQuKcYZ
0215ERjqLOvkCIHK0HixGDRGbXzLFFXOiJW/Vva53Jgj/vI7+Uly2bdoynPbJ7DfKLApnnWddkl5
6dnojKUKvCRRFkyDTs13UEaN+UD/pnpOYG9Ht/+W3/4mq8ilEnMDwr+dMQ1CAneztJ37jJGJEEJm
VXlGTkoxKad5XyTvTZJ6Qk878qYSkVEZPR3GOYeJ/30NjpmyQYkgueRXapNeeVLgi6RXxgBVUMlD
0wXtnpzu1L1/3KC6m7JFXD1xPkM9MCWCQUHitgSz6UAbSHWn+bLjx002cR25IUanMMryp7t8mQ19
5j2dmtNljJfxExK5RdsG1gAOThgmxSF6mxv70RiOQ4cSBAfwwORiuFBFGT8jojgUnfvV50YOUwIv
wvxdEsVoDfEEugHzPf+OeExy3w7zUh9Y4MuObuMUa5Y0zHZ5fDSJfssLslquUPdLxWDNKZioBitj
pqFgwHpTm7Fu7JAoRa+nbpbyJ1Pq9izQ22wMVKTILObWmBz5i9m/Mqo9ybP0VHgWl++IPVVrefZ1
oyiQy3D2s16jbyiRvndQ9tHf45G+vv0NIeJ+DCxs+bZcMgRJOHjj9A6yol218JwdPg7xmsT4RkRz
xg8bQdLkrP5iC3CwiiI4oB1OPR2TjU6+/1BxDVi4sUmMr0YmUncxLC39wgUDDyAOOANBXbu5Mcya
M9MLEk2cP8bdx5pBDt59ZSUFiFFe2eb1VVmUpE0kCeycul6coC1WG+bWPeZvTokhPT00kQakYRhP
afZhiRXgoPsyeITUrtK0mS+9EQhZb0ks74ju90gsIQSKUJWx7+V98+/qPdlWyEgAaypH08bj2YxM
X1JG2gOJa9R42/pwYub8Awt7Vmb7o1vEf0uIZEHDioCUyjgasQ2+tr9UPIofF5K5hxOEmc99GfA+
1Jp3YmRISGi1mPlX+UQiH26qcD5UEg1XgqLofJYlHriNI2kiIyvyu3vI69TuxXxGMRDGGR8kOMzg
yFwvZFR36oy+XdE3Npjw4odYYLcOuaxGZcWhQTtxV4kd1fMTEYDd7Suw22hgiRRgUwL4SgwkQ/q+
zmKKeQUY7qy5sFOHsciISCf2zCsttfyy/l0rPWbXxdt/31/3JlwF885Lij+vaxRMLzLBfURwRLnU
+5bdytIEQBiMkaHbAn9g0xSy1ywmqKImiDi/DLgPxVfPcJUhUUx1jq7FcqDalqdrMLLwONQtCH2D
HtNOtzoEH6q/aUQYrWTdCnxNL1nizGoZmWuwc3elYyjQpUVrNl1LMQtrEIGY1IF4ZcI7rY8/wJVH
nz8xZum6tTC2AT//3n7hLaEgo5J4P+85USmukSdhu0iq2yyHbdg96wqiT1XusAwoKwvA3LRaLtiK
mWYbeBVYEatcqHkcFONtCcCQZtYvalfdUDLChjEqzylDo5gId7X4YkM2PG9DlilBWQhgxfOsHcRR
GFw0kdM8dKSMPRqOI8iS/j93Yz0iPqbrLPqynVbSBxQTTWJdstwznVQnbd6eJjLUh8E1ogBOV5KX
illHY4O5CqrQVd/G4M1NbExkZsnh/+XGleYqGYWR3iKH6tVAFh0XUhA3741SnH41OaXCBAvw5omA
zh/to+SvaHWHp+CjPG+QDtWkuHHu8wYS+hraoiAvwuouRjS1YH18gzb5tyN4upEAJTWhTKRwe7t0
Tfs8LKqgZX0qp2gK/O5BMZAN4WZqT9EGnA9FWJdGATY+eBhUWtiFmyNnSwCxB+Immvw39r8jq/yR
8+phiLbBSOsOmd+zaO6yEsRZmlmPB/awX9N/WxGvDc10vvEvMlua8LITVf77RKaAMM/1K+p1BeEt
BYx1xo8CDH6hzWDKYep4bKawSMnOSHVY9ArsSdIVglPkFzQ27K7Qlegg24g1mTp9vRgl2EqyjidP
2l32HHKfUV5X7v7sIWwnYZNgrKruMcTgCMF8dMalgFH9P+gYCwtIXkrrj+wWxajqkRGVZu7awuJ3
BafTccBms87gySl2F3E6ljvvZM22kZV664pmJRgZ4+5R49T51e3lI3Fep8sps2IxHxFo4CpbnMBy
56v75MJ26OjfnEqdomnfbsyEW1yTp/p20uzZTRjAbL7zLC+VWLnFvROlAKZ1hqEFsz3sMGWec2Jl
9j/10qvAK7HHbF65eu6bTrx4XfYUd17/jRpJeISeWGald1DwrZiEpJyb34/OxbwkIOdPfXgEDhN5
+QEhZ+65DRvsL2c3IhNlNQ3/R2zN0lsZImNs032DJL/L34bbkr9NlQSIyzlOIwMD75GwISKj+i5P
J+Sn4XOBBQ7IPaOoNUiVjYi/xMOjSFw2C2SHsaksvnITHj2HWFxT6YS37/5ZTDZkc2+t5Ck0ObI6
3Oel5njMcq3g5xc7sXZjd23C6PWrnV7irjgPwRFpayrAlAexrZE9rek8JAbAEyEu2gDFN0nBYSXY
y9XgUdUrzf4Hi2PmvzKW1n9rhuYvOuA6nNHE0GaFhaQMtMvUByeMCnb6sTwqG7cLJOU5glp+6J+q
vOFD7Lki3ybcRYO5lH6aHFC6mK8JgFf7L7rAjv1NzBV8udbK+10SbL64hsxOrAg4djc2SVY7d+gD
5WMsN/Slp5N+/12GD5hk9DCYB632Fj0JNGieeDkbwhQ5trI7CAcjxvbPH3rjwihYyMDQT6K35dJr
L8GqeLVVzyn5N2xyY8bsYZeHarcTp9FNevKUO7oCjBAfSSWrX8//7FCEWp/BmgTkCQ0ScMOlG4EJ
52BJnO62yIKRkHykqcID8UZoWEqelsx69Jesjk0BFomqXiLpw6CbxhOcleUweHahhikxL4SqK5Fl
XGVob88jwcrUkJ05lCoM04oCxVOm4a2xie9Sp+WYPgyOWfWO3mkW5IOILMaq5jPUnCrNbXulRG1N
O6NnQnR6YtLq636JaqoVkVTDzYAPRkrZAMoimYox4VNlsiL9WjY3VBRPa/6rSjVruSd6lnEoCaQt
eCmHjEcihcVaicLAdjT39RZd0ppgs17hKRuogQg+Bmz1sA9eOLn+R+CNE9LMzb+86IItB5nVsDOB
mNWlymb/NUvCiP073YNnuXi0c+LRJdIJwv11oaXyYaEy7BzNaOMp9u7dOv2LMwNn5WreBOhIng/a
oYBKzvnORnb7QWT3+uDiku0Hbje914zltCBnh7J+y6aqpYTjwM+snoylgQx3T5pAQzsTU4KPF8Mb
Fgawf52MoaKq3ymL02I+/+qcZCJSH/6p7yAFLPDMYRTF4M9FmnPyWv2rx5ezF/O/3zMwjBagzjFQ
+IGCEN7YuKl0fygN32LDq7Gd+0vRptWao5ztPplboU/hrs3LdDj3frhJNU/yXzMJOmAYwx+Bsr08
/NMLuhcW/tw66DRcD0Ee15LGrW3i7euL2Ij3fvLtiR8naz2H8LStizgXACjaSOx1OQtIdmo+lUgs
Os/obMh7Ff+Xq7BzoUBsu7XGGJMBHgKd8mhzhEaIvRCnew+pyjSZhRRWr7q8HjFCxyttdGwJoaiq
FH/GDn18DGQQcycESwEy9dUM8tbTZ0R8PXgU10OTF8s6t9y9akiYaQKS3XYqZW0uWKv39IHLb7ls
RaRBcuBBSVj66G8P0laC7V2XtKAzdGKU6wzpVUpKChyoRYtp8KcnueCtP9FrQDPtvkIP5Nz/kTNL
lIHj0acMO5zI5ak8+bCO7HFFEEttNp3oF9M9BIdzUqp99YiYaSig74Zxx1u/TTx+MMiNdSWoUuc6
4GwgX+2zo49i/vtYzgg8vP8MFqnu++H9Unq7lOHHaiD/hv898+YmBL6wYTeXpsYUcvBNzi6wjCX+
XZ44Ij1Po7q7Pmvy+0Ptg7SB7I3MuXLLC7TySUXf3KntiwE8v6+r1ok9aZ/Y95zHP4zI9HHYEhIW
lK8P/1A8Zs/dEpmpVKsfUlfemYRezCgTm9lB5n5VDjyIEVlfbEAvyXHMkZyGsJCVmQ8ysEbA52Or
54PT3ZfDET21sX+gG1p8tfFpDHmBps/jhsTAGJXH0751berZYQHxdDmZOXw8kmLhW23kfkDZprNw
CPZ46CNVw6iIFloA+nFrsLkHwXNYO3+AnyQbUQHH8o4cHuEsLFNWsG3ysXHLTWGrMihO4YKTqaX0
euLo3P9e+nQPnJlXqdNU059JjZTDzzGa+9fNsfTiRqMRMC7fdq96iulHE1xez1M1wscQ1gk44Ks0
VMrTyBS16CVireiDCgtsCrjXWz6STimOsNuquErU7mGzFmjkQh5QaOEi4mhs+TdD+aifUhCLpscS
01mqUI4hwh+V/Bqezvo6q4iu16//8fWTzqZQLkFWdsVBP1ozwkTcTdrArjS8BLWDhdKhTGzRJu2t
B87CqrmoJZoK0qDn/cyTyFloDJh+AESMlT7hySsefDM/33BvfBnebtszWIrHWJj7VA6qgwr+qlkO
RGBJzVEVArSCn8A2/Q3PfsYQOnimqN5KBAz5Y3z+KlraSKOyW7ex/LLJ+OriNpgZpykf8Q/Fn2Ze
gZ/ivoszdgpONM6kawVWfo2J+QybwBbOs/RNPx6t8jQ+LaVJFqSr2N0QIRx3Y1O4Hk1Kdm56NhWq
Tl81K7s7oXv+50+BGwujKX65M2vPPenA5c3wHTZbX+SClsTvppQFaqjkk5SevR1GeH8yBKgMkXy8
+EnfMorBo5Q4fhTAfs4oPivf07A9tphoL1JJ/DRcKpHiuWo8NPcmZhCUGo2tVTTkgZKEVINvo7JD
PLPpgYJvcvsEvf5Ro45A0z7eSLsYvQmvs2ex5VKMKRgsq1OwNH5opQzhAThcj48Oe1RHX28paMYN
x8G0M84DmPt5eW/n9AJGu8g7nCcxeHLPLKha3ESG7K4kJXYDadBwgBMchPZZFyn4NXclDCPsHG15
3JQ23fZmsey5iU0gyLSumQGgqwcsJ+JjdB3ggA5DJohdiV9oASeFetditfR3B73NB3ddow7IMxJX
330igEv18uPmyqkukH9oYueiCIxvBxzbblE6S5B95gLO6qUd1DIwHFv/M64kNirgYv/he2Yiw8Hl
Ib6+E40OCcN7vrwoVs+pbdYlQS5iNThRLUO7VT0ELBaKVXRqWMhA3n7BdhNVLd2s2uN4nlWqx729
bxr15YazumSWXocCAo882u/dx9pIvdMyDiSWror3YVvdSUR1AEG2r+FDofULyjocA5+RQauN4+vm
wYQVF1f3tPDrGmKu2qxi4/EVHntvHuPbtPN7+pRceO/IFZs+OkfwGBOZUiggDVVb/hpBTJyEQlvi
2PtA6otRXVpw2nCa2i6lVPJ//OODQ2pvvSXPTpMtGa/ptrwv9mzHryGAhcj1fv+elmbm8uRfOp0M
ZU/cvu5qZZPJwdFSZMQj5YIxsrIJJJh0Fjku4HSEKAZ/DTZhd05d3Jqo7n+o7TO8Rvad02T/DV+C
43lK47nUKjjdePxlXR8wXBHD2kkSdHH9FtKSC06uIZiP22XsJwnFMhcTGseHygQremp4YwgpmJ62
s2LjCfeiL4edf/baclatW0/j89S6BbMhVfwRB+1HjESmfHSuCuHQbFr+HLZn8v1tfH79RvGHrsH0
E9hBc63geJ8qxlrDJubfvqhv4uoTMnieP31d7lwaNuNO3qfnwJsmMZlRECbQnAYQ3F7umptqdQ4K
YqhXVffREzQuR2MdITRulCcNA5RNnRbRHAsdQqjKi/00O088hiHDibAIu1iAE0vk+4scAl/8WzE5
dpWOo7zN/bQKLxBg845oo+I2c519z+pq61wU5Juh0eFv2TkLfLfBu4PkDBhh2De4XjM2n2v022Uq
r+IT6TxlMcdkOnrj3Q6tuh2Ku21H/6IHdsBTc9m42OS8Do7iPfK3W0Apux2a5kLYAGKOGY2U49Nt
d/xxY0Gzp/d0uy3my2Mzd2QOB32uLVOyUnEin2uADL6SY8M7J8CQXCuGoejWmwbRzZ/9HESwZXRN
efur54r4TWz+Hx7eyBjIYKkRTlKdJDVdQ6tiudmPU2melZGDQt2YC51Xmll/zBHUGrdq2u5dQgLY
5UPBSfBTTp7b4Kl5I4g1MuKG1wIfQ57QC8hw5wW14epXlOqEGlLseEdmL3hG4tgYYIHP70Jdu3V+
CJUI8/2c5peOy0lvbqUU0aGCeO5e4oD4Fx3CPmGOxV1zKuq0DznkoLKGKLexUYqw4nUHPvyYVads
Bfa2LLE2pTzCwyGtdEmuMTqVnh5ZJljss+P6lEsjx8s8LJFxjQMHXmJ6AIMovYQJeqUHi8Cr0sYk
iCdWw/3y5TC3eW2wN15gTSe2GtM5CHFaChaDa/oJtjZJNXml952cUaepl/w8aAMKpBjccuzgRwub
o0BkFcqyiIDT9Hm8e+SGkMWnTbrKRHbZLcgEHLAuNEq726Fsz6TQdtiT89XIXQUN0iORTXtAotMb
GXgQ4RCoRhzrzVU0Ou42Clrw+AhRTGm/y95S8eu9YXhYwG8oKY7+sexf4xbdVfFEPdEeiJt4VOfc
bjjL2YoU5y6FpsZJymcSKziFFJQzDKramPYt46nxuTHuIaPDLFlSL7o95iNDvu6Oot+cYIyOqoVQ
pGPZki36jxTizJV//Dzjegfp2ZtqfA/nP7GlMgnToNj+ONvmBbYV4r/5AsQIX3hXJl5zMtZHlJ7a
h31h0hHWX57cq4C8PuR6Uk7v1FxwSKLg/jxLpgsoKSP4qzEbQNMaPjjP8h1XEw0UnFZsEsvjOT7F
Y07Vszc8YE3jtNGmuh+xqDae5AtXc+2rATAVHvGb5drpMXxf95QwR5GGqRqfGXsW9dqpgqCtki2Z
y3JzwZgSfiBmN2KjJ+mRzf8kP7or+W27o6lYQRhNnEoJB0nDuscaNqbtY6O2W7POA3E3thdYBoN9
wtU9kNoqzL0u+5o1WBQib/O2blEuzmPiwtmoCPvOJ1ljt8hIKqVrQ3itvcoSHlfLN9Rf/jkQSzsp
paHuKxveOJaacC3ABcP3XDgMbyszFVjtfzczRWFYUfSBZ1fzzOY80cRNcQLL2lzQi28Z9+inROwn
zox/OckbY+oxVAvKz6x4RPxik2riXEULbgPqoGZR26/bLKAas2QBEGyRnxDA3Sc4MshzTRW4rCS+
kZC6EvnpZ3c7U0vy4FqwPHhbcSNo0p84qKQZoHMIpVBE8V1BJrGiVCZ2uxP1pWZhXFIYEctfthy0
kt7l79GhHdROAw5Kx2fHpkHNdO/e0e6r+wPwq/Me6RPjogjuEBPFcTAhY07lg4y76Vqrg1WEqCEY
Ord56YQ+RCrEuByPDB2h6dNu0ddHsA/xZyfKOc05woVWAS7GF5YQvqg2srcA7GwqE1GKL0uIObsv
vkEc1tbBm/AR3rOioxYcThoQNLU1Qh1CuRPvCi/nytMpfJYowdy7DCqetcjw2Na/BJ7VuCEPGJVh
euNB7pEiMNsBccYpTeCEODM5/sPhtq52wgzRXN3ZBPUoUtdnp/X4GHQlDlw3mDVyem14RB1HId91
VHUyYWdbWgUuNxHUVJe+0gFO299wAdeQRfnhMMEcDTIxAOmxwy3NLGN/9CKKoTXzZXJdInqOIWlJ
nrB6L4JBZIeIvD2S/EbnRahwlH774pzh5U9FMwtQa2V37bB09QW7qQmuiFv2rBAKDaOchh4WqYXv
HHdanU0ECw51RdKJIvO73vnLIpnhGTZDPHIC/OItpIaiszadm4aPya+Irz8KX21yg+5NWDKqKBb2
+bf+yabCbO9u5F83ycgNO5MGj9lKVLv3UQrYmv22wuAe7aPUerSVVDzW+g3d3lAHqxd4BJG5K9XX
RbcwBhCHVtgJvczp7lZj6uhBYsFLrUfubFB6eYF8q5MNi0CMHY+o1JOmKuZdkQEebRJ6XmMWAduP
xUHGHPHwZhWzEne9B08QRQmiX0CLO/ipLg3qGb/EuKxgzembHj49BXPuH0xngw2/uyISPiB/72CF
GiQpyqf/zB7Xr+RkHZb6JLq6Zyf5uw0wL7Zls+rumL/OMMPcYrUQFr2kH7ajpRagWOMaxYr19BYI
N9gRdJiahG7Qv5aLVuh4+yomhCArWUr67FGgaFcCiWSzlUpu1JtvnZquSfaSdMxzJtETLikZIjjG
+YyL6vMKK0/XS8kPrXGwlx8C6OG7qR7j8UBfTXaLwzYCB/yVO7pIGmL7iPIIFGNU6vghopA3BQfx
az0JKiENNZzgew0WSVKx+TQurbQzcbBdVakcwq5ZDS/EP2ysKlERw/3GX9pRsbxye+UzI611qWwl
bzZtMa+bQxMX7v+knX5Mx57KnA2JBJ7K0uZYUg0Vh0myGbmFcpUueJhFIKSmNBD5jCSenYi9e0z+
I6ENfZkY/ZLd0O3rfKujMOZOpzstVdekrC5zkbcKnh6ZuhA6D4Qpu9BhnaDP6pOgEOEW2DZGiN0V
p8f938hJM22ZPdpwoqj9ykRhqlceGGmwG4CEUFAXfW5jQ+R36XwS9aLKh/M2acNs9A8daqLCUcam
FXFoSRgUh3IKOs71gCIQCuFsBcdA1iqKzU1+7VSEHFChBRhUM42+zLhrlGSdiKo/tzVgNvE2OHXJ
uY8vYFS2wp7FxmvEQxAzK5HmL01jtaZFfQ/lINzrFGolmuWFsOc8a92dcr5Nq0sTiyIfHwzbRGR9
39bbAURy7gu8wVva4nmdbiVbQPZLXOELYiPDGhfKcgWRlOpDG0fjPN9roMUJGW9JARpALiyG3UDu
+X5XT8tjZGbHj+yZ9uoFYEtdy+ENAoMlukuNhcUeLkaoMy3cEKAsv8zNYW/7s8O7leosjKmAkTW9
Hb6P21aivCqMlzhh88jKz9Lspbg7pIfmNBF6BXufKh9PLI/moL0Sn0yqE9i4gvgAWTz5VKmMilET
L7Fbcd4r+EQEcCkHhi30JXtVu59sfzoRZMj+St/kfq9uEcKyQ81+O7lguJdYnaKquatObgNBeXai
jqSNHowEU2DZTqbXRy58nQWACAUpMBCMwmjnwPDSYlOvcB5E3xeBjiifSPfXrO9sNVvnVPiPZ7U/
cGrxuRnXxtMD/LZeEwJy13dB+Zs7m53ZEkkPWhyUgfXMS4TZDdEuRDxIfmEV+Z1+KxmioJcQ6gMW
rAsne7coNF55Pw+k3YOyIUb5oPrY49irbEakEXhY5tD8uv15nfuMQ4f2RwCpGeCfFdzNcajDO2p3
JENCcSYhljJ6bmT3bOTo/KRmMcdiSYI9n+U3D+ogDjA/XkrlhEmJiWqOKcdEuhE/RlKG9rjdGKa9
eCeFZFzFClGgNXLwwn90vZwCzVJjlRo9xNLkJjAP+1pOvmW/T736GeDtTahWuoHlJU6Av3uh5NPn
ajgrHSMeO8cFiJGiTOKBHd+BRzxed2MIfuFLGXGqJRThH8oSVcdsPHb+l5oN8wX1sM+Z70e6EqGj
9gVYhK2lKTmXItBZ/jtmsR8tl8osQVflLQOBUgIp0hRZWy1DTrILKQdVeImm7rM4cOUzosMZZT1s
7GbtUXgAkYdDblfgLvPtmQ1n5zuqrf24n8WbDOYmL8YAnWDPD5w1hNy4YWOt1sP8R4S0CnA+Ybf3
/KxARKsJ8hFzZHWQkUGYrMbTrTlFxRhrRG6ukoX9MAQZBjqaOvgF7JZh9rMKOVIDrheTcrsOokvh
5wA2WZCoOnLYh/d1nnFry0F7IW16fgOkvAetxgFIFaoI4cnLBfdWFhWNhfnTIBDXlPX7x9opPQ4m
OkCnEmxbWr4ivUjtK9IIvpSLDC8GP/Rp+SQEOOI8NjEC19MTG3KtuB7PN1Qo9TIDtk9EyVQ3uAhq
hTz1+hJKNsiNVPJX57Bdy2n0DFJQ2sXsY8WJfNWZ1ZYenrvNoKj3ZFakGV96obEDTY0Q5ifQ4c/D
ptEwakGVh8vWqf6tl6TbUrYai2tDiNqnIks6WFRUdX9yTRG61ooUMbLBhezXHohdHPp4AvjTtvCR
pGav9zkoKGHg/VIodeO+kW2iUduo/dHEQBxylqmWMJM7D7GdugLhELUlcEh9vvBl3Uqw7gkr6UUk
ddf0THXb53gxq6HIqx0tctbx9qlA9r/QGVBfgQYlPQFmb83ki/SDlCpxMlZ3h6T+FxutHha11ULW
0VeflAq99TUAz2zcNHIj2gp2fLtRvH9XE55unjyaRrDRZQhHirgfTG9W5oe947g3S9k0AJGiS0IO
cck/jsftsPRH0vcjLan7O03Rk5N7SXp0oPHACywdBxUaKQLhPiSSmGk4OSfcZu3lwoVbFs547Kw6
DPNzoKnLTyEHqqi8rq++vhFUk+1Fdza19qC+uwtGrBqngo8ujrqnbCzvDjvVOKLKMnTlpaBQfAyH
whKLnuQRtwR9VDNogf1DJmaknXosC56tvl+7LnPej8SHhj9ICjPtzuAzL4mopvwT6sYryYqT6DrX
OEzPkSvnkbXlsHYcJMMPTWnPJRzPPUv7hbIJuy2woVO2NvcQnl53b7+GZpSPe+C31GefbvDkaN/f
8ELG9pDlNsZku5ZpgNaU6O3OHW34Ea4RA8iCyhUXKYJtJ0UjDBWd7CBJUbi9sQxwhzzdAPIfqv2e
i4SOGBwH02lrVZtc/DIBE3JaNxCTlq/K5GZtnC/GcpPsOrtD4OEvrD/qJJWrE4OzKntULTZbyooD
iPBDN1o2G+7p/C3yzk344zVWajB4v5mPHjro3QBZFpVZOdjrWZciQ0hOmGruvlVCpBa9EH7Pn2Sv
vbBHaQz0u07oSetkVAod+64Jc2TBLhDyoF13mxJuft4zLG6W1ik8Ig2syl3HrbDOylxXegRd35Ao
t5ha38iRqO0OXh1b/hEJ6RHMgP39DcwWU5kjTg0T0cFc60w9pv8NEGLxx8r5peTIvbMqHIkbjy8B
U0qp8xEm+rgEADFnxc/hVySc9IR+F1Fxq+knvHzIDBqWyPPCmTSWXMJlRJcICLfkwjLzjoZex5kW
UTRsLIyelz4m8HQYYsSkJt0clmatIgj2BOuYOrG4WO1V9mJg5p3og8zAnx0cyGWlVaMFmapF5eop
wFuXuPkWv4mNazpaAhrJmFcaNBaP736z4p0YmHFZsq2ILELuSJxKLwqHHSGt03W6XIEpVGrc+Wrn
bdZfklDnHx+r9e4g5vbaAINDFPLBaDncu73ZaMBXsknTyhD+Ah2Nn3n1Bb5ffa00DP91BXvo+/t6
ZlIANNewDEgDmBEtA7AF43aC6f2W3Vhj1kEDbh3+zIGG/3wQ+rd768vmvbd1xcKMav3cDQhHi1gq
eyrr0sLfKKm4+jpEhcr0zKaLMgjWxMHTp1nrI+g2VImMNo7lrjUXM8Jrcdrd7Y3LMKDoSx5FeCpR
iGjuF61OOtHUInh4Q7hu6xhxWnt0KGJgnTPJ2LSSBarbgK5Y+Z4u5t1buOreZM6mQrYqCZ+Gy6No
oQ0CZrTR8QuGmWzth5m2319gPIGcG+uZcoEYFhWKxda9vTxHmMZ7v42ncP36Wif6XDVPiY/ndQRA
eOtEalY7E0BxEYTTWnyfHZvgm3Z9YFSXkjCs/u3TZQh8WJQSAw/Ot4ZdYR6iay98yOR6e2ezQHxU
kqENpAA7WE8Oqt4jOPHLNz8+tt9b6h21+jjW/NF2RONEGOKwwThujo0bng4E3tGa6IaWouGf4jbh
ddVSmZuIc5XOiG9ilUfkTnCLaMd+wwfW0ODiYkgimiuYvB5FLzSz9dZq5McKEKChfoohG+FFa8sr
SkCp0kygNfUmPUClA6BUg6k/vdLl6Q1eDcgpEnuJbMM8Tpyi4npAZX3b02z1+RePWMAxCpf0TPEK
z1i/wNh25Ag2NGIyUdYt72qBlcv4rUlJX4xkxJMj+gF7Qnp5260cW4f7XKGBSc6VOw17O43NRKHh
kJhTH6petEeZ9LKFS7CnfyHEajMi27RFvL4kjDol9SHYlTkSwd65YX7dBMORMqvC25+R1AJXVMwS
L7vkjrVJcpywwMwoGZA2PU1yMHpzkONluhTdBLQcDm+KHc6alz2ODEU7Ht17oI/oo+MZg+b/Tuos
8VgMdVD9Hqw7sdwnlaErS8P7iWADQ6kKvTenzkai8zBg/kYWviw0gvFP5ObBebJ6rnvHyzl5vrqI
zC1Bs5anJi/1DK0lI0SAChX+gwqJKJ9mzIEMJyq6srtxfMhTXsCeV4h1O6liCxYlwVYxc77mTo0K
afUONX4aDYB5WUIqW3iRq1O3ULmqnrtfWyoXOwVChZE/oUKmC4B6H0SJO+duo7HaMtFJ/98I70V/
agciHhXHbv4hRxMat9OsIKOf420rNXzO8mWYDAyphMgtbOMNRSvau1f5qt2Rc1OCUtXfCIEivZJN
oXl99JWDyrhSnH1AbzzVfuzf2TNpZ9zEonh2xhhgQwTm2X1BpBfs04eC5rmuzxt8vpC5hVSWxxbk
btulD/Kef9KOYPx6cLMVX279NSQ0TpmvoiAqwAtNDg4G8Ue2pIB7OvTihFt5rd8XAmIrIe+TZxuj
jXhbkPkdzFilfdVr01bLdKUs4kVgAYlV3SZlqZuuE3DW2eM4oHepEk3TisQTD4ZTjQGTgeRvCU+b
Ar0+WhYZvfTtcYo0it/dU2EkdlAhKiHS0Gg5Cs+3EvVUy5eqIGoP95wHqE5ocq9TvtEALaQyf2m3
NtDDGjCKENLoQwwZF4mr2b98BSKIuHLRkTVYEPYAsGR7RQW91zuF5A78juOqkji3YWY9ZOFc0dML
iSY2Kx1+P6sRuyJvF0Cva6vlUzXLWjA+p2JU6e63X78m4KG40aAf3l/1JrdylDRu1e0x4hu/mSeF
e4SdEm3+Z4AoGVo9yH4i2h9egD6VxtjNszikji77DFG8HOVv+iDTgDtg7I6zjJVG46qhNOkf7iyr
qSkYMEFcftQyq5yd4k6o3eW8lrAGJ0HkPZOgRfTPLtuVcQa84JoJQwKHybp1RRpCR/IN5PhLyOMN
B8/Ix/2UmhEdI8I5kSMdiTTK8ECzIN86U1PghQsjJvqg60aERRpRs+zC5OqYGhZzXOIb+otsx4Gv
9c/o0zYiEp8RCIrTrxuDSPryQZG9VTJxtSXFvKHvRlVq5scmtKEUt9o/3beuQ8u/2V5W2j157hYq
Soda9UM2dvW3flC6GgM+kv+D4/cn2YIxmQMnFwZWZKkDoTgS84nW+rVY21ZTZ1Hp+F3dAUsoNj0+
G7cOEo0q4zo8/rxcURcoesCRhkTpgUM2T1gDOs0i2VPofsShMe6JjfeQpqjoqxbQCsGuxrWjKiFe
zHslQUNaIe2Msw+2Y4zeFwYCjtMvClzOeJRbZVJXFEX7UYuZHsVCSO6O6hyFheQmi7wgs7p8dCJd
WlNxBjOxCsGZTGMPw/SQG2Rz4Rcj/YFHRf6ATvyeYp3FTyd64g86iCfVavMN/4qjbtNA8pxC8Ys7
YUy39hVhiiuHYCP1OwcBhNAYfASqdAhGPnZKuZyjzuPDt0vIMIGV1g3TfHPrEnM90m8pBvfafPqh
8G3p26+po+Yje6Pc9x66ioEertvKwuxP5xPOH+/EggQCQeR89WOxoeSbYTyVJy5eoddZ+ZyiMpFq
iYu9JtFRwDo0fGdDFsqek3INjpP6Xt6nKSHzClYqSXwAdQTKjIxFNgGqerEI8vwPEd2nFx9lhp55
Td8aY4awI2zA0sEcoUqrEfdC8OnvZWTGOcY823q/pN2PW54bJtUU9OAKe8PAxd4BBF6UlZc2QQRa
OeiXiGzMoWT5AogsuJ59muWAIRI+xlLOp5WIlbaDP7zDZv8M1qdEyFHG0L40QvmJEI3MjqdqnpFF
KXXk+yUcI8QXUPxJqA6h48sN0oBoZKRTyNf9KnJBVy197gz9fU1N18PJzWC9Uw/yDgUGrA4q/aIv
aQ83MyCu56xqpK+r2/aWKbkUgr1to9Ltqu6+JXheU5/EyUnyi+k0oyoTLqZPgZFVqYG6adV0Cw2L
oy+jyW6TWLmCGjxZk8sJKklFilUa9cD9e2/MyZc6fM/zWW8rGg1mDx95wDHXXEecz9r56JsVPsQ+
ttURX5xxzJw64Zw0ajIAxzKw/Gh2kyF6da+rkmCQKc7CP3UgeHWs+24C1+wJ/jn+bFXlmOltmIYa
tnF3ibpE80YWpUGyERjpaolOucilqQ5mSQSwdDLzdh5cDymalxm1pTWU2isg+maK2ZrUIZdS2Rv7
FXRY4D7p+cu82AZURXJc9De7YEUXvoxqJhH7CbvXMp9+T9JG7D0nmF0q2zfGqZnKVrNKUjil9K7R
P2S6eWXOnF9+mT3QmkSfm3AMRU1EhOGjU+X/oSNRcOMG5ppYqEGtswDME1r1rI/MHZqYZPv5xuP6
Os20XvE5YEuwpNitqkgW+nuiPl/3BPbSJZ9E5TnnHHOxwvWTZD4K3IEVI/Vdkoin9zWEF6z6HPWf
WS4K+0T/+FTTRLDhRj3ky/ebgtxK8ZuGmwX+n5WQ7dwHTo6Xf9p7TW42FO9/KTd3Rv+4qYA45geB
ZtvQf2Q5spj6DzFn6yoSRiQNIbobi2T/aLMJWAMP5Ll7+Ho5UKbqNqmGyCL1FVsVkyTwceQbHNvV
zoqc5XjA7/D74EoiisJaNqYCt/410OKw9Yc90leBB8vdZ/eg6uXtruf5eVn3oYS8yu8G4tPbvNpt
vTVVfEi9K0AxLcd6arIHCJ9kxBC9mytB3yBBKBZcHyLvmKfDvCfMEK8KkbnZqOfClibWCWtgILxD
la2CCBZhg2bGZJ1wJ566F/sOIonFXD5cvTPWx5v1ipWyZ8gtKWyOwqN2rt4gR/UKZBeDIhfeKaq1
DcHMruKhvTiO+z/DBmBSGz0TmYY4ipLSDTjX9tAVhpCYMyvvOe98tBtIKt5f/+k/4e1J6C9oNhYH
2MXk7Ri/ti1vX4Osf9wYnJdLiaviF3IXmGp3UDn9f9dxkxUmck/2KH/wBu9zgPlCW505lAlEAytM
H4G7+0Ei6D5Zas72gTl214cZP3B9pDeYdj8GNlUX0Z08gWkKS9uXFSj0y5KT69Y/RXWTNxxgiWJV
qZ5nyBQMcfUjO3cXK9fpPKkb7v5fII1UQ2BCdSqoR4tw++zw8tlYWfRIgx6jWRCBY4+rl1SbQmLw
7o0lQp1LVnOAt7vcDjla4lADrpGsMoj66qWCRMffI2wWzpD7aEfDAJ8RpTWVVG/OgWrArcaS55f+
6MdnQzVFxEpcNHdcKf8VY6bl7yOq934lxYKQ50NSst62mENJhSi1dteRFdOILP/Z09Sn6Fh6GNck
j601VsTQ/CksqDtrnHsDdPuytWVwsM1nbwretOeaBu7D6gSfE7H92Lcr43EVyVOi5o9wq79QpRt/
AI7BTkDydJPdZ19q8+Gfegfkp2cK8+vKSeorgnuCwLoN0W3v0VpWGocbW4XeknMoKGgVFE50qLjb
iB+rnYghX9mJPa7B94VFLUUfZ8Mx+bYwymUh+NuocTSMlKZZ7tNiBOyKpp8QVUYBq0B8SZzSKvHF
Yq8vcKuR7bWHWVg0ViQpnupyNCIx0YrAZDgfaFO4fwzWwH1mrWJWxOQic6ksEGVdzXiJm/+SjuPJ
blH0yx9ximXBoc2koxau2ativ8lWmSLkxjlnX6/x1urDQ6TKC8TqWc8FlyT3aBQahy/a9GJdpUcv
zR5/5qTQZqVaeIBDK8Cc6grgpOvf5oPYi4EkK/y/M39MrV03HaY9MkQS5mTn09i5h0YzZ/8wFSCN
5xXIoUGzPVuySoJxlszEGKeaO/nS9v/Y6/xjZfGuJB9ICxEnWRORTeGp9i349Eb70Sy6wC74+J45
uKeY3ydQrnw9ezBcjA/DzbQMCE+UdG+fuU/Trt/lX5jwZuehH4vX9+AtEe8GDQmTjz3LRrF/mlcT
zlo0aWY0knqBMn7MjSQK9PXWvLWqEUC/3TcT8I2n9a/KJVQumByH6lZYQHwdYlxxB/lxk8BbkvpP
jHgF6vunRzlEP3j947ptAVuwGRWOR0LtBY6ptJTc7yb4QMUcuSGkfu3plJL0YsGQS/F8ANH1LSRD
jZaUpThpK0WaHOcYtyzBS10cWqY8S3AAwBdagZSSxVZolZTKf7nnG2OCI65I/ZHZFBnpWmXK4R2L
5MjCPlQK194vCzydnnNPY5o1l80I4DlrdqkaYYzxkgcKllT26mNfyGMr+8chpY+bzCfmD6PYBeVn
E9khcSssSULOXK/uk6tZfhXvNwFLdB46y8GEIS5q3xDS3UovZfzYwwa0Dzw3vIiOcpNrxXBYpqZl
ScO+Vr9he0KLpJcVpER0ihn0ZovTCAwNrj2r1e4Q0+RJTopOtg4WGDskNhcesxssPDE64LdATRu1
O2RTczfcU0mji71GLu8HPvCo8SRoT4OF9LC7ZiGB95rJB6gK0l6kWDbSjD8Te9AxwwZoai//0MMi
ljpnz1yId0/75Y7kS/hzs1Vb4AWqKnDrSUoU+Rni0AbTa5Xzp36v8q25Un+g3ztkS9DnclSyLq1W
U3LtkjW96aYqTbo+nCGOqD8gqdbPWwHOiq4QsEqld/xVSxSftzc5pfwiNYLhWOkZSKjyCf556YMt
mwwqjCp1umJEYZgJ1cPGGhP0p7hAgpsmeLgepid1kFIlYqzp+3IKvSmzNuEejEHJmIeM5lEKc+qS
bu6kaHxD6uM2+B3g+nJf1/jTzu4Ymc5NPG5In7TlvYZ+UNNHZpzQbFf2X80RwITqegxOYaL+omxm
SzO26RawiW8k5W9Z8OclueQ8tt7bJrEcfZIWTxwL+J/xDp8s9nP60AB912mLGiahIz4VPTt7kfMh
KifCsKE7L68E3/jgA4/UutwZqqtrMBDyFo0PWaJvWUm64AVNDHcXTEBqNX4K9db6qBDu+7NvEiVg
sekWZTZXamqDR2CNNZhx6fRtHbSqqhINHhWvB1WZxhyUPy+X8LdqiYmvOYiMihxpM7sk7s20wVBP
bnaHhENhT4+pcXzbveNiX8pgynIuF6NcyBi70A57qPEUOkrxvhfIA/62rZPmyMbvt8iIbHWu0Fhh
gQUnBws/wAvuEFci/LwOF6i6NxgH3ciNQUt1/G2+5mNWwDhj5GJTSsFaAaxoG1tIJLDQUsJlv3cW
Iy4XhIO8Znvytr4X65k+FAhjgiKYfQAHfB/ezSXlpfyf+DD2PJ6s0j344yrDIlq9wIRquBK5uDpL
6OBVMBJ3ZsX8QXWozjSCXacDGr/G1vPhRwOpmD7QoHG3wcsfaMhvHKK/JSQwvo2Xw+G+kVHEs0lE
ldhmjOe0eFYCI4Uv+LDGhcu1YnWFhWNZz9PgO5Twhc+wtZXBzZ2kmB0cef4D5f25b+JBNPukM4Uk
4ThnUGPU26nlrP6hGDmC/RO4Ot0NBF8EluAcO8PckhdUMZoForM/QNAg5IAo/UzWN78T6AegBnR1
E2Kq9RuFQIh6ACMsLMOTuJfK297jiJ8heBb32Yfd2TRX7InQJSQFf/iE898r2FgjFerREEicJekF
q48nITa/MaHwIzh1UynMiteNkrR1v86Mp4MkGIqMOQ5yJJr21YQB95BrF5zcnAHgX32+xoPrmUTF
ol1LUN+f66OrzFB36s4lgyjZaCBL4Rk1VU5dUZ/Ls8UxDaHOLPGqKwNoWP0EGWLXc8z0E6G6bj8o
+90dQq+lcGUC1GIAV4zQEysrLGBZiWOPOK7Nvp8xEWdqdnOALNLOddGklGBPWLWSuqdduQ3C2JM2
wVaBkIwJ+p4leDy8IzIEUkCg2LKsT0QnkHnwbbu4UPD0bcmk9o2M2zDhH8H00i1f0M8kN0YMBGrq
wOwKFdTa8PDTG9fTKkfNA77gf5sGakMM9s2sAdsPf6N2orYsIlSIUEWFsImfThg06LXtHc25tCTN
cO3pug8H8olLRkqkChe1o5LjiQi6QnGCdGrZ3ZBT3ZB4UWCy2LazyzK52xyJK0NkrBNZXTqRSscv
7KuB5dznGHhhhAdn5AjZNjsJHdMXAt24e9kR5b5NPB9K6SL/K3e92gFJdWBW3RBunBJOGIynWljW
B+zpyGrY9OAFfNFa7mm5cSi8FRFQOg9b/80viPC18A4/CF40+1iYMcjO0Kxd9nnQMwYsQ+oPK24W
K2J5Qbk4ULYU6stVgJxwa5+qFSTdTArXo+QiYqBe+cnldbIG24LvWTxP2+hqwl26l/vZ+NiaP2b8
xx2rHus+i0/1Xt5WNj0Pro24PgiofKNQ2BTyIt63yeGp0Zq+dkA/ReGD9C+igULg253OtSgvkJ+V
5siG/21uXHklhZq1fvFCje9KcGoqS+2Yol10tUDwnGVgPIwLHVERyPcxg8+OWo6dOcqzmlfTxPci
GHrifsr8B/qa8oPNEIIBc5VClOc7iNPc9OSulLBWgHo8KBiRenASbRI87efSFZTGHS2Jsv4YzquL
JTPebfomPARNpEfComypvnD8xcXK13vxws0kVDYZVIG3rRreddK5Lrm/oviy+9o8+A9TgxoFS471
DtkxfZ3rbCeTeS7/eUfArnBzROlluyo9RSCaLyMLUf8Ld7UuwRtDBTVh7pYLIlHEFETwbfHgDq/m
6m7cIpuVNtl4lQ9ClWFzGSsC6tQtH56YS0rwGPtujdjN7wCTE7oAYs/SzQxaAd9szHmC28vzQh10
VNeg6Z7vhqL05L7T9wrdXxSrb2OM6INgPkmJ12R+pW03ZWH9mk9JMulbLtGRKQWUhrWnbFxvTt6Y
GG9fLtlBPbXRlpVN/Cv/ka/WbhRSq6eaGL5CWNVJwrUuZtskZnkA+Z6EROjcilh261va0RLeA0El
jID1TU9sHdx6nvHk7U+HMQ1MTxTQcUredjTppYqei9azVJ4UYyvSUv4Z9N21pKO3PFw9iiNzeW2R
a4wjHIrcjpVGBTjBrJWjq5K7Th+o3Kc1MjcTEWxIp684uWbt3hVZ8GoZXqhQb+utZdqPpxjQ3WI4
l9HtJRXkMdoS5yMpAnC5I67pR9BYRS4zIpcJH/Cqg8voO8v5Qaat6gkdAU7aPeKiMee9wgkBKcmK
VQWOmvy8yuNicOivHNZWJoWB4iamNBp/h93soRHIVq8JoGMxhbp2mbFtBZC1zyszhUKdWGyXBjik
IiAHfQ6bc4q8hXs2A9h0lORC/JAszNZUdTyqPCcUvogzc0d0vYQIAZYLyeKdZJlKmNTSr9dfcQWS
KpYpVgMcWULNO3YyZN98czNAufDwaHiZmbU5ldmbV3ZqfoYhmohd3gr5xnG04xQiVe2iJGuy3SMh
VOUtUEAlC0bBoH+ksYsOYoGFg4/WR4YlV/IF12q26sGbjxr+BYfKZMx0SU+HGYbTsT7b3qpUxr3u
bVf3H0XfK4Tz4o+MDgmV1PQO8Zwh7NL6XQXRPyQzSymawde9aVWQk69ecou7Gj1LOx7KDmvibpA2
KJY3+8D3Lb/NBaa4hB2xtYf4I8rm5phnZGuZ5ewEhrqnVHAUNrqjA2+5JG19QUTNcXwOmJTP04q2
678MLTpBua8EQnrshZHbYJlHOdl8ug3mTwIMDOri/lYFQEFu5zlhamGcbFM5x0bdiOXqZqyzT6bp
ndWGceUu/M+gyPgLw+YIy+3LUsVcUapcbroI2rThw6FCG0WsC1tg3pVGsPs52NX/TRVC0utzQPu3
9jZyfuU1lifQ6JicS3alty/ww6O+GzO2NJ1kRyJ+qp4eVOL4iBSefZJ+rxjfLedbhzfLKhAYqVWz
1QJjXKLaSydfmd0V22kBMSKKvniWjUCaT4Y092+X+6LF3ZFGSVysuAXa/A9APE1aGo7eTP8xT/0C
o5RHmgcsQbbUgouiO0+mJ87de7VmI1G5oWusnu0Ei+frh4BitanFbxsNj2JCgFMDYyWu1AopO5u+
xutuSpK8n58npi1fNdvY4YKHedbSRn7RbbE4p/xoQXZ+2RroeIaW/Q1ZSozike3FPW6RCcY3z6A8
/qIPRkVuye5D03IAIH0nVjAo9CiNS1qn5KvYYqukzpVuZZHRuakkpWeDnn/rVkB95Z9QE1CWHDnv
QX6D7W1e0+nEx4+0lg59fzV+bDHkYlmADDAEoeRecXOUqhc/YRX9spScf/GuGOlrPpc26sNcIQFR
XlKoaEyRSRmSBt5LHvscJb6JfK3tk1UspSYib6dqoVnoqeUGt4C34SO+8pMn3ql+ZXL38hjaXbjc
fMycq9iOwnddT4ptr+WDW2i4Gq9Vxv1v8Uky5cnjhZYCQ91Jigs0fr+shgXhtyeu6B4gfLQYQjfZ
3Y3IQlURLa+nIkzlj++oJdeA3wtquvravKh/pTovPUtinGBfCCG1M0nhlYEuexFdU1yVeHTcN0g0
zwUA6at0zGbcUyjy996ERxjcbXRZJpVUxZ7vVvaK6v2v/VQ3PjwVILjgvWNVNd3VQC8//bqiH/6P
rAms7+KjMdtEvnG9RLNXH1TzeOFl6rWVZwi61EkM89qhHj18nx95ub6j+PNUkjeoV2z2rpeeI0gc
a2oWRh6PWI3lTOsZc2xShw3ujmH+jLrgznCYuU1DwomAeIy0OX9zGPQliFUcQWpbGweq0nuFwNVk
xj7I2UPgqWCrN+7s+9K/7SLjyXZ6JNXwX+01fgaW14RJ5FUxPaFwKSmlbH2znco7lxCkTsiRoOno
k9xEJOw0mZfEO5APw4CZEl9NxZXOVs8mt6yCWKNxtunjlBg3744Shl4a6hu0Y5sfMKV/asitvwQx
Em/YY3hgHtgo+Zw962R7J/RaQnsZs6ni1LlE5uOOKKPyblfjEqxRggHqPeOrJUbN8GL/MpoehRDM
ro54zookQmkTnxoAs7E3cijvf2zI/7q+F3NGJSlL35x2x7uMOskAycK9a1g7DeF2FlUnqe5fakmA
Pjg1UbLoaB4YkcY0pD4Kecd4NT90LsX3CkLcZscbmJcYte7LKptOMGJ4/49UWfYSW84pw233TbKb
Vqmwbt7W3RzMm4h0FhWErb6zlqQuVstSw6/QJlwWnr1PQ9MUjKMSQweKZMinSO9GTdw7XJhyE4M+
sxQG/GtPJLp0GZgyigHDzErrxW047R1OWnlE30SqrisJS6b9iBAnYj+hdIFaVq70pULOzotodjm/
5R0Ear3xFIyEWXDMScmIBVaM9Y1zfjai4TenoxTRSrL83esWCnTqvJ04mz2LCAjE8ufyMU/xoj/k
m1+Rrm8Cu6D5bcC+rih2pZF9gWf/b1puRcRgZI7CWOJAzSWFTw9elTmDWNxMA+bgyw7147Pth7Er
j7Eqenj1t5OfSCkNFuE7a3v5WYKDqGrr3Mk6CNWP1UwK144xmlCPIzTEdLVzvKF5ENdOZ5rPb19R
/w5xLsV6zmDuSUJkXR/C7SNqmnHgN2DJkM3wEJ70lkYOe4O3QP/JKmt6HWmB8gtaadsC4zmb1GHA
QOd5UqJsvxYtSZYrh1EXPmTooaB9DxsEpnsu4Gw9uCM27vAuKZxTvhnlbPDpP3NLfaS+oEwJSJHq
DWG9YzVMdAfdXQ0C1fi+Q3h8ee3VI2c/ZFSqkYahNplAqw1HjGY2s8YJOAZHSN48ZZnknDGNIwyX
NubC8t8w0vtxzYUI3LeIM5xiaEAApLeWLnaWabY+J8BaLnX+YrP4SaUcsymJ2p1IfZLWmH2gAUpH
ZJdTSBBs+nUljG0GhUHeR6pD0Lf+ohqAKq0joYLMe4vFHZKnuQ+7P+/GUpmTYrDJtIQAspILewV7
ShHaDvWGZPnj3+39XNrV6+ebERx9NU2+7UOfvMl7wlO1MlylOhuQI3b/JgbKnZYM0wONHdIwtG9b
hPCdYOC6hqcm8DU7GeILqE7rtFzlvI+ND5iAAUrxbSkYtICnqCOy5S/FsVTNl5/AhZvKLNObsyqk
ryqZcrYrpXsLUXoZFjgQQOpJ6J+FUiMFuPxNAfwBzzhzoeCEeMLZj3/ePyboYl/gwn3aR8dqbaek
j73fwYJ4ulZOODrco2Tq5Sd6bJ880hYO8kp/TZL0I7e6hYIztl8NwvT7GPmgm7ifv1oYfyCvI+Re
UwJaH0ZEJuG887iCYEj8kwr7HReiqJ0P8Z3MCdW1qNplGHx2vC9wqjO1zowk6FVHxuYTj9h/70v3
3KunjkhTA9JD5b25HI/qZOCee50/dGf1Zkt+6IVRDmhBjK1QCw7aorulaHYaw9YMonlmBF5mYasZ
/fVMKdj3oMy6V35D3gwd3CjC749sHz9UWMRHmbrBDEcJ2VLNSsNSMsOJZPyIcVGD4MGEUFCoM2y/
d87UCc7u+E/KiceinZhYRZngx2HUq4fNpP3cvv/7xLh5X8LnubD40FazJBLZGoNvEHG/WFGVXMVE
mGhq7YjMe7VGIiLcr1rcYe0nNiKuzfs2/4eZKQpFrNanqUia3dUj983v0rNTJ/tbkkvaLkqWCIse
75JhsvRBcVmO1cv8933/yK6hA9dIxtztNxxXay2j36/6BegkbNQN1s7g9+J/YMysNresWSWfvrMs
9VRmgNUy7V0LBGwt3af+S86vVpAOSfRpN1BOzCLdmMgAN701jykpnalh6pnXVN4m3J7E8VPIWHh2
kqG91DZ1pGd9fexIV+IAwdApJFjqHDM3yTg/ibUDDCGXx7WK+XYdlYPPn29yA3+1OTFa6LyySY4T
s5ssZmtGuEch6Ei/zkWHhw313v3pa7vc0ADSCGIcriiFyos7ORTyLAdoew3P/861h1ueohDsVi1I
bj6ycTkVVpDjUyb7fflqGOICjoUiwsENg03H2tiqwpec9OgBIf8B65mfn5GmAmzrlU0rZCS/gm0m
Mt/wJsUxMt7dGGB8yyJ0X9mUKQ8zj2EweyRNOJ7qSXUpR23/ttBMbU7CcmbZmWNcEEXUHB67MpAr
7jKO1HcscrCkjZ9tbRRlH1jsbtop+Z2yQgt9SERSX5QTgwNqOv25DC7iJ/Ei3Cc9c7QlX/M0bXcs
x6xcaze7GcpdUZZb3XCE/3ysm++zKBeVVXcOUZJQ5IY3PRIrnAxyqHs4bgqUcWJYwsUAh3H29EbN
VsbZqQGQrYdAWchl019B3WrLakt8ZqyKWjA86EgYilnwbcE//4+7QFYG0UIA0Czo3q/mPQ8WC7za
r+KGGbJQbAF10yOzx0Ot70sLb0M8G2EM4jv2XrJHHLbwtKqhTp5sA0qyUB3JBzdSX4UJh4UAlWDV
SZWqxQsHfSE824jtQcJ3VG+EGvLkHq+8y2OAi7mEez1NmYQZt1ba2sxvY5JBZPgiHAzWuMJ5m7Hh
/jvINQD8Km+Q8rlVdCgQo7nz2cAiJuwP2/qNMd93TBQr6D9CPzTi3ZwxZ028DrnXJ97/FyfPCdy8
G61X2OcUPFy4HetuQPQh0NdGQXZAj6tuRATvdZujmGnVYcGmZ+ux+02cCtBICz+IxcErMf4xjD2R
YkUkXLczOBJ+ATy+Zi674BTq20oCoN7KfneAAH9BbcZLhL/sjBS5Cs5qEJMc9PkLVskBMfBfuLCV
HuODjqz9pIjbnKUPD8O0cwjUXXlt8uFYmEL9K+yGlVR4YBPDQh3JMi18YD5ZvZ4d1cXBw6mjjjqq
ESQdQk7GoWanAFMenAyQhFRhvtnOlCm4OKUO0ruMvy/hS9eCM4gSIxXCj4ku8ZXTkPRhO4Nd8OIf
X0fpcw2jv2ubj1DugpHEUNHAe9rocfoK1DewG3kRXO77FhqY1kDFzK5gTQp8x9aKc6VqzVtjYX6N
xXGjV9/HviF/NBou0dUTUs8Gg4UXDBAiZa2jVvEWlZdc+A9CD1uSpdaPdNPwUk5No3agETVfWYXm
cqKj/wu7rvTrtldL/ZEWKuuFGbO0EtVw9UTWkpGk4UIi69WBS4pumLlKCXwWVXeux2k9C9CWqaAf
jzjXrFCU9oSi0sQP2Xs2VVShwbwLHTVtgYEAEe2a8bGFSUMUD43hV3XgSxIrqEKrKZXlTsert1DT
7dvhYf8J700lztlDspfvOBoObgvdI7NjmeeqMDCltuNkCL6+kS7Du2s9jA3nidubgcDbagN/2SXV
jV6ItYLKhliTYzesC+LAIbIIva2oolRwe9C/EAh2AV+7g+01PMhLNR4sTEWndpQMv3bLcI1ptyX/
Onx5Q+YqmVl0v9tR/kDLV2ikVH/z2HUuTJWigULtgBZF1/R0n+b2BCoWDpWABGeKoQsYgkUCZ7Kl
tbjdxXu4evifZe3p9jNZnLj/B+7K32r+A4gtuhhPz6AEfEOrJovmzk7A14qxPFoiRY0RM/epzWew
OJsdYA7FhpNLsDkmnRxNYHkCIO/97p4LWMpUzCRzRp7tXFHgUPuzVS1T5U17ZSaPYhdhROzDIqWC
DLtg7XCWZJFsyuhWnkQDUF0E7kMpT+qhtrwfJSfOxO/e4x0iozArEVj6dMqtXD+62nLen0w7SKd3
IZx9VIChOwR5G0UisThWVAmTxmdZPromxTxtgwiCheQLnVMVkZd3tjCHPe366ohSF3CxICgzUTxm
TEW6CwvZfLUYMYymwL+JbeiZCzC9dnWFTyGcZWzuuC2hGtZGDGYV+t+Azrm17P66gOy5OrCq2FPA
CiiGr0OU81KwE8A/xl2R/SxLFryCiMR5eglrt3YtxqQ/dPh7wmClq6/J74ikqJq/apJ1jK/Njx7q
0kXRH7/AQhFNFVCPXxU4i3JJrmpiSp3HQdiTIdd5NZurzHoKKk+pbeLfDPAUQyYTnOWh2Ky1xrUW
sgAVOqyVepmlIhB4B8MQPgj5D8xmyulmZmn4GkF49GZD8UgKiN1aQFhwoM5WU+JWtoSe6eaB5Ovb
ylImJ3yyVYE6N6VlO00K36I29lLLbWukBJQG5O90l3ICU57DCGN0xx0YcIlYyRsBfd9yeaFAEJdO
cK9+imxZkD0WdWCUpU2+s0iN0D7gLR8MXpe0R2DM1ic/3Kb04SQUSJLPF2HOBq2M69QOEMu8pyqU
N3wGumr074bqIiDt/LrGydWyyXCY2c1GOC86tLg6HxCZzAVQcQdpiGRZwEiAUfR27OssM+riQbnt
p/t/sqtJ2JUH4l9Ld2A9NqMO+0i2dX8dkj6jZAukajFCQCJyHRlaQn1cDTXI62j0x67fedJS6DCS
9XH9A3/g9ofWyLPQRQmG85ULqv5Lb7UlP+s/yhJrqADC7Y3eSLbOtZb5kRiYli0rHw+Wy5tPWrz5
uryygResEnnEcoTSh62RP45u6HH901tbuzD8CfiKdY5GJ6fhc8VXhyuih2+7dXVfPlCokgLq1qMI
+rsGovJxOB0gjxx44dpH4Ijsn6CXaIH4RYNDRFsqeSDscUCrgYweOWczgbl8LLAA1EjgQb2aADzh
jWSO9jtFzkgDsjR3ikBvsEfwUsPhadCA3W0VzOdvOWNTs7N9i4HJHcVymtaqAgExMm1T9jEGMhR+
Qgi4mttg2Hd0jOdp39WCWxs3szgmRDiU86pG0GgWz4w+SxUYr1MRwvn1NpkSla7LI4T9h0kT4Kkc
ps16I6Eij3E9daulvd/RjRU24JytAxz9robBynCpcENExy9vo5ukkKrVeHxC6Cl69Qte3QXZodrp
jRTR6P+C1Gkddvd6B/8ySrsfSnnzH8YJM4RPgA3LNtfBbesuI4vYfzwUy4dMRMHjO5U2luIr3f4P
U1DfjtPT+46te7+Goe14D86GdPe6El6Jiypt42Et3rPgURnqD0iXgZb3CTBZSMeLyujVQl9HlP9P
HkSS87nn2ayn6dIk7rV5o1rWB9UdyS572jJO5U8EZWw0W6ZPqOzB6D/tF0qNm+piPWm2ZV6DiIFH
lpcJdKtoNuozIHgNRzG2QRNTgg1EDqttUluJMQV4n+DPIqEGE7/WlLhn0396Jn7VCbQfTo32Xx6u
qa+MZv75Q5jHksX4ZCvxMDz/osA8U/G15JrDpstETD9/2slUnYHhSjb80CQqURiCD2gP0+MEQ0AL
y356/AhHSvUQF86z0ttVt8ysjitDODw3zFVMa/1ovSKTGeASW//LfNjCiXj7DTFmlP/NEnHTPBcs
9xL9nTGrbLA57ADmboFjnIF3X2VOBtpR+t+U/d+XAr00qEtA9bnW6Nvi2svKMnZ03R0+JAiz+f6Y
snYhWn4xA4RYUVogOH29vsxHkSFDb/yDvK/90vHG30+hfTO8+MNgZLDKfP7K8d84dUAm7O8NRTc1
ogWx5GDs5MonMxXF3rsEo+e7p7t4W+E87uAfhWMtVF+Zy+pNqlyHQsyoGd1ysPGUEoMLHu7VIO3r
qTUpSTcybC1reE65D78VLVqu3PPdsbHfIPmjjyZFQCWguxavqQ6iL1sVIVcvnxnMAVJvusuBJN0P
qetUTHcQ016lIo4fINuZ2n/1/9/2WKBpXk3Tzuua7Tb5t3HJXXsq1+gill2friTz3wpTUR8dWi7L
aC2Ps96XgFEXxXBwd5KuQKNy0F9ldZzwrU/BCW4fN6Bug/cdReAX/g4+AJngVnM/bO+hvnqcOCUl
9pLCoD0VCzawhNULtUFLzfSh4pKOkV1afsdhif83GT0eP3Rx0bcCsxgurFjVtJv1KeO8ABab18j2
4vqwbrNgUszEBPAOdnNZUmwgt6wdpUw3z6rplDUxU9U/riG3Nl21qCYH/d+Um2KlXebZvDoicrfR
MUVd/pKyS8MsAxQE8dwzjfZlQPpPBFW4xxN1KjeMSKtRmM6d51HSTexfBmEW6dUT7kXvnVIZWoIG
wMJ/sPHl4nbmu8cRioimD920qlFckbw1RvzbognogCZKzewVBRaCnVQg+qFdfNnxEyHZcQXPhEzt
dXhyvwzMsPoM2iP4KtEZyTSERtV4y94Mpr1oC67AOpc4Okx83JpO+OQpRlXdo2PySjEQEdwp242J
Ogv15PBkdPB5zkw8cVRv8IxquQUC1/zN7dghFOw3Uv0an9l0THMFUssOyk4rBz6dkYG+tMdzzNKC
Zh1O1urxh3JnxSztoFse2R7oEU2gWftlhSGbG55Q34IvEWmTv43EsFuY/MWPVprLRd0du9m6AB3R
1vCgwkOFtkuupOJHPpFAS459D+YfVM/2OlhCuqBuWOMZSKTJbfARX6QGOdzXIZ7MzmMdArbSkZYc
qOvbPG3QYYNAFfq7BX2Oy3jx3yKmNInb+V6xT7DfLL0aaF7Vv/g9V0QiAicEOwXCK5oBMmt5/b2T
XRq7wdIGEQTAgPjHU7lgV1eqKDHrl4ry945JTPWsrNFnsQpjAcI7xRtSsxljVQKcHbRiQJT7v1Dk
GsPq1SO9W28PI4Y4ExHCtpAwMYKY3/g6JRFG+bauJ+pO9+W2D8rTSC53EotP1UJkf92mazOXnj0A
bklx1U7GIfku6E3ZXLPDPOQOg6jAdwgcVLPcccKHGheWSxjeC5AJRlPsUy/mp04OLsSWdrQpCcsk
85jmxad9TuoFCaRldERf/IF7Wzva7zDnstXE/uP6J9Xg3WDVaeEZ1r2mQm/bpHx8ASCXucqSTxZe
IDokGg5kgGto/asLC4zUYthybX/4R+IxllANakCW7xl8hyXNZ4d1LnR9A6eHpvWgk1dvrj5I+gcJ
cj6GcfsgEaqk9BAgfmPI0Q8LKtLNLJKszO+wJtUXCTPh2lNFpjGPq/XqiYr4pzIlHULXHH3dcMCT
vZaxzezzKrYvjXL9h7iuxvDAVz+45Dt4qP5cRd5jf+RZtref1FF88fNysYBlHZeYGOvDcuD7Toct
/AsHXYxCLYn/8/UBs1tXU7bgjQZu3p37Yx+PisLY2Ny7xRCrXI+0NaJxmfV+F9n2A8ZwwNp7aF4Y
n8GBy15UcLFXlg5ukg4rPjfvPW1noY/iuUr+yTR52ikukfLnLmZYux9aUoOLMsg0CMY/eA5SHeVh
mQvazCgzQNtvdQufTS7KL3vD9nBNsps0bEIxc45udfYjZ+5rcZbAE95BRx6Qy8gDYJrtZrWh63GY
3D6RmsVupn1YABk+eIbqEmwbJ0dPLFkzGk8VRHhMVdVZRmZbUx2BkNHcEyGB/cPQeBcYbR7k5h2/
rk+gcSpXeuFTMJPddELIYmzOvcecZmr8XRKwW+tzuYcPN2Yl2NE0Yw1V8ZKLIRBoYK/+gtUlFcoX
77/oT2EMhycTCkaFVCbRn/G5gjHCZmCtPyFc17Bd6ljCNqDa6aanoz/1ZCnypjhN3bjX+d265ISJ
3ItiyIwCFeAE4a8qV83oxKIhO0/61tMnVsYkzxTMTQ/luepXz51dAjwE6PS6BeLyE7GGh8/hyeKu
b0RC9O4UQ5m6ofLX4Z/alxqz6gEIFjFQjw+Rale14hBygInqxoG8inwM7vSm+PgUFrfyt7S66sha
7QCIoF7y/rblelyO3ItU6hqxw5zoIE5ePx1+13XUDpPbXI38yn47kRASYIUiIIhzAnpwBS9uh583
ctehv+ZwGvoGy65+Kig2yUpUsdmISN3Lq4mkhjh5B+sWCmnV+oLASVVO5WVZpQOXDnHhJ1XW5urK
+5PnnmbQtwE3K93hCdOHhNIEa04yu/3aBsaWT2Cxz6yFJvrgdWmO0KqQ3cAdquuSApSHQPnYJVnS
h2qYbkBWDkQtSkdD4vpsBvl6eWJEDV9TYJrkqn8leGpr3JessLRkSObNKUEbSD8SNNt0oqLko1PS
gGbwQctsqC2FiKVV+GXLnEDXguTplUzQr2Bf0xLYpoDVnjaj1SyvuHZBmhEEb38l0Q4r9q9aFnx4
2UejKoK1/7OzwjFGmVYlnIbmnzJYuVdnlbZcAgATqetFuEeU8yOXrt4ocIi1W8Zp4dRgViEwEaBk
4u3v5XgMu8djp6aUjeUmEAO/UDoVTn1Y4IBUD2jFoy+VGOIhZYpXBoON1q+04YcBUKF/CMm7ZrEF
0M5IAdgNqKQxV8WyW/s67C4pyHsZ4d17cdTMeGJrE4wyMX0N0l3QpnTkYKq6hssFO/YvXvYWubg/
pyKgji60yK1IX7bmg46WDaYwtkg54gkT7fLmNrJ+YWIJ4lUHjDu5cWKxNc7dbd9Mk4marmktdgei
RW6/XttAH22zILxDvL+v3BofT2Syd97bZ8edYStfL3EOW0yEPKkY3GfWLnT5J6R1TA1IW/sH8iHw
uw9WPVuFbYhpY1SVO5pNZ0qWtDjAT+E31a2fqUw+7WE+U1YcvVKW7Sx0xYc6+9sozCwomcFsHxvt
74Q9fFsZml+zMvTsR5fp8T460XSyfG/8U/vttPHSkjvvKAUjFwzlrxHNh7cWW4QTs6HWpfvtsRv6
k82NQMpQC7S/LQIbqeNez8QKNWViMKYHvZ4tHb9suT3NK4GXnIP8kwtBMoOWeycfHUShhP5t1FH6
G+hHjac3V6IYU5KhrTw86+7WKI+IcFWOG3dMviH3C3tTuaEritVDcN8zwzXFV+HcE/iMWTvFGUWG
jT4a8Fi8HNn4fnk1lafQykxK2gMCIhzCGLDW93iPxZqEYnBS7I8sXkmbJzNKxGWDrzXQ/9C+cDSv
xIqd4lHwZ+MFabBhpQXyHRiI/gqvQUUBJdsowbwtK2FHZDnbcTaCO7f5PpXYB0u4YsoEvTwi9pL/
oRdpl3atcT/HWXERyw3cutzar837QokXc7unJR1YOYOdRTKTtCWBzKmLAGGhrdVPgGdEC+F5gMLX
s9ZEW+svq3yfIU9BBpYe599uW4Iu0BLnxy1O9K4n0IIsbnWaw4whFRdZMs9DStyJLYaR6VA7ZaAW
kxhP+Qmyd9Ga046XdJMh4ZlTIbauQRtVGrP1jzIIPm4Ni1gX1TIupDT5F3WODm4QVX3ZWIGobk6N
tip8ot6keoZoMy3LmeQesAGPw+OVPXpj33J1IbG4MG630tg56Zl5ZOnmfjpqP5X8vlExaxOD/s3s
87WxsCnU4KEiYA63A9iXWFmpA7os4OJVmz0X0KwCuErH2cSKXKAQdgHIwvuV9VU5kjQFHEqrePML
7IVKMswH7tRPR3uhyW5AwwF/cg6QSPVnthftFnlPtfKz3ldiNr6TqpjM74A9xewFOcKKGasb3QXF
daPUoXnlyX5hQUDK4g3nSTIeWfJUi0TaEOUVexxa/rL7QNeBxj0bJh3R3iqHpf/REfbzYSjVtO41
LpTg6tzWlvzLnvAhlatSZHyKE8MnWBpmnMUywzzaxuPxXU+jV9A5FaAyTv99rDyXhXWtdQ8eKs6g
9/1mvyMbt/XXdKuytJXzsnBFNwLPLwE0jOZ1H/Rub5Xz9mnxywWm+Eoys+OHBmH1IJ4RcUNr87S0
vbccqFwHaVXkiKU1il/npa09WAjFPGOvJ7JtmfOmq1w4MiEW+WJJOkiJ89dVvhUmofX4Vpuesulz
2dm61TJtaRflMRkGy6AfUwbhAVysW9CaFxEC4uaXesp3tlzHUUkWoWWuf6DmdCjkc8e8DioTj8qq
IEyWD0IC5RQpt29meo2/UtcFaBGeuOOr1DMcybIjHfFtiMu/CmNVyqoJZu0luLdZKHxbN1OzKOOp
WnHhH1C2G+Ga86wZTF0rUjspi4ngOc33AuxWurs6aIle4+EF7hSGsOqVRXynvpWFO0Gu8VLZO4of
Nv4yK2c5p5orFm2eYAsbKNmTW16GOiE+yUzG/f10V37q0I17VevNA2DGBE0AFsRtTOCESJyr+NiL
eTNPQONKKY1Gig3u47zx/OEU6xew47bBh0tAnG+QuOzU76n+gnMaK1qvJwjjUyWQdWK1okEWRbS9
AaR0rJXnXfOlw/foCRs/TSlyxpO8jhP7pV+d0rCTbHZ+QSJ55+s9/bOU5m1L/UpQ0+UE7+4hW5JP
wPutSRi7O7yu2SHd4T9QH3dMUwy4xz8YqfeORNXnE34uGOqZ/SaQKgFLAA36gEcDYknFTqLr/FM0
OrXSEM7aQBreKZeNxMoHkr4JMYE8f0Uzf9qJGx1mPm26eOCpQ7BDKAy9uzzrQmpZdIAU3IAJq82d
u4FhaDIkfRCEsZvmTZrLSMDKLoO9HjRhgBJcWGjMt9U/653NRHrPWuYdff+W+/5UQluVm9ZDpyoi
P/kqzQiJooTRlGiaOOPv3mCuv2qWUDGj78SsabKYD2z+zsQxxl6zq0NF6xX0sJTJzLVugbiqAdtT
o3IleB/yw8gbIf53q+ccDZ9/5U+JoZewGOjBrx+YpPLQmlPY2f5A1zHZ5Rwyxg3aDuv/w32FPSzg
g+aGifEMNKScmr+Ht3ylAaldne2N/cdwcyAyVDWc/wg8EGuluIFe30WWUa01+k2XeMFn03T/PNsJ
yiBFiIyRX1/2c6RSpcYHbVEpEH3yGVPdVwx6MYS2VH09++aLdFsuT0DjBoguSHIm3FnqCSrMx3Ct
oCuXz6l5zKnxPm2EnAnijurFj3IC/XnYk5atXdEqhe6ycOEhLgSNnzxmAwo0F2Xt2uYpkHf62bZj
FLvcHuxHgqaIiSMC82KL97SUmtzAm2nJaIAAHIKg9ruOsdk5K86LjmPC0aA+cKipymbU07WQ+L2S
In0gR5ZoVJn4lKlmlhcSuQPCZmxArqdtBDJZvmLj3Q0q+Co2HuSzoq/brHquagmEDcogLRy+yToz
QazGUDBquiobUJKboHEnr9z4+OukZQYMqeNlXRJ2t8fQARCfUObCt3HoZRNMd+e2Qg0UEfVzzk+5
mU+/9ZR5IQq7OuUqCwFceqopcrfMicWIi6kDRdbNRjmywg4N3vL8NxqcnEZ2KFxH3soXRJskTryy
A6qOxW0eG9AHMYm/5oV/XKi2TvkVLAtKT/0/rF8FwvS2gbewb/LIJpKGNBET9yGNFrjO00OjmtRH
i0uiwmWHmAIN09MqkUSTwe4lBxxZcM8lMkGg/ImUcN92q6xkfeYEEHvXWSX946CR1eMhq2MFGfVS
7Off5jCh1cnOGkOF92GL527vC+cO8mGDGU5a3JlYxJJ16Q8R29f6Z7O6SL7TmOG1BQ3j5CKj/wX+
CwP/bnaztGVCvkrQ03NjhjY+9w4jgPaZwevj6SCbSoXNjSl598v634DaTKvOHMac1rQM4poUUedc
7adwp3zl0/dvpzFhpQQdwgWvKsaj/9RJcqvYP/+m7jIeY7mTFZELN0JPiBa4M7mRMbwSd/tB44sv
7guRDoTm0RREbyXYLbgTQtyJQVNVA/7RTmYo0hmCcMshrX2Ck8q21pMSI7ss2jkJC25YfvILddCh
MruGrpXvpMfJEEfgDbJtQWwV0bKzVgA8Ra81DmlnbUq3vgNepCHOvNkYrPlzEMZAx+gj6k/EjMzA
eP7+A18oNZKzNts86FWFTZRYNDJupqQidteGqQbUNZzi8WfrqXXMRH+XEwgmVr9B/4zgbtK2XTFA
JpizypKJEVr0FfOKCSQFCe18oX9J1MeUEp6R6VV27oywCTPUUV611udHWbmSL43iZuoVvJU6DL6N
gCeirYNCLB+cqcbTPnbHutOAy3UxoEDd8z5xpWjHyVJ63a0CZQd2Slebjrtg//eqILBxmtLSCOIh
rpDfqs9rFC/GjJ5hp4ICzELhO5Oj+94FYe5GCZKcYsK7rhFvStlPHPpBpYsPJBmU8bybA8MyQaBj
B4JHqx4c1+ZZLTyroQapbmf4NH8B99HbbZP7vs466/kZ1+rfLl89oeHkxfbqzlDoJGVuS9FyDTLV
ntfTJGVZs2QHhbTBo6kvOizCs/7GIGZC//Woz0NvLBJx7vET8/cKfmUBH7aaxT/qM13Ibs7ShQGI
dpV2XMTmuZLqtNu23nv9aynGlEAiobQbMupO3IZM8Mxv0jdbT1P0toknbwSzhWCW935X+VScFSnm
Y8Mf4jMrrMAmEh/Z/EN3Vw26XYXNNOJzZZ6Tqc/T9Jn4niTVurPo0kDcoMCI8GbPFmw43okq6rp6
Mx4lSZkfkIdwU00QjssFfqIyf8gRt/XgvBvuwLEU64y/AMUnoeWakud1K03ivuuCmq7LML2mtksQ
vqnS9jBGbU6mKOk6sonVTJnvVeGIYqud0bR8DT7mk0nRVQDNGlgAa7zsoVYrPdunVCt3so7dfN8H
N0AsWOJRGja59CaSBSoJCzBUgfeVaS9y08QytgMbXWEAudjyPSgR+zW0cW4aWJGNNOrJiknwAfkW
oGkBrSELJOdAlto34UVf19IfAIhvakxteMvlno5CMRo/6YdMLZXxUH8/BQMOV5rBrncjoOxsute7
JiZ8049aNICmlFpLszY/diWBCLNqwZ8yxTS6qJ6ExO7SvwFfzZVhEbGyDFDlv4g9/GF0/zw/Xzeh
ngEDNQCu9Rplpo1ocV6nd43MRcWBXtmW9xO+vzisFWP+82hBFf2bnzrGhTtqv6i/R9IKMi01ovRI
FMLM22A9C8vDvRUVLX4ukHusaxW3rqPufkrFIyJzVAzV1EEE4Zgnb50mmD9kCKxdDDB5GPU3xMQu
tA1vokbUGiGmvAnwfYY6ErHnC4OdrhUh+vgWrTOuxWEA6Im4+wr2oT671EGS63AcJokNPGgE+19a
G5ffdPWYiW0fsWRTOOhpDH6bWRf0O8i3CqrIcrE+0kUnnw74RrEo+p9RU6ii4q7Lcn4wlbr9iTC3
t6TnxN3SKue0oV6KtGFj9X6jiK+X/OVAOQLMA/u2GeK/hMBhg49k2QJqtzFeyyyZJH5FvtrQ+Sbg
PKAODP/JtXT4Ve6e3NrOztK9tk9uh9WPxT2/EkBnA6fosR0eb1Fz7i6/1tnymOIrxpTFHqLEY7MJ
UpcvboFimaEsHNSSgmhPvrVrgWeavai8ahjwElRaR17X9Ox4i4U7bs77MeJTGZoCChN9p7F64205
DoOV8yYIB+9GwZlzxoZe84mFMw5dL+fYbSYQVoyMhJUZqKAPYhCwQMW8buhcdvAG9WUxS9g3Wh9K
T0qgsQbCDbxF+6qGhCDwCrWcEZWmFAuuFEbuXHeOGufkhU3O3cU3FLxMosEq+V77BAVzsNznGRNF
Hi//ZAcs/jgsRUUEzkp6cqbcZK55GvnvLVIJzdtNKCIyhPkiw8b2xDeoG+vJKs8BUuvFvfmZzuWK
H0UNy7BsK66iI5HGxINmyHlK5nsQcRrfx1hHoscJReDRh+qBryvSC1kaWWhgcbSbK3WCYRqXVt3U
IFymtEaasKbaSElOgwh2aB4H8TYZ0ANJ+/59BVF6xTX/+5dh7GNywLwpg3WhKVLVCiT3rJ53KBN1
PXFmBLBdZBbgAOBViLv4zJq31cZ7AL1t+NbWJ7XS/LrZ0Kwk+kxowRmTjV1+H27Y6yzYOI3wk0nH
LJ+/C+xKvP138NEynlhy+3BR9vM0+OnLJaW0fkhep28cuuXIJAnnxayBbWge8gThPGm2x6iYLVni
iY6E9I/IoqGrNyFhHoI9lZkj2to87x4rm9EkO8hCpK9dB49TsRnZSCFcQuVLedgBQhYC2x4fvfFg
nLHVDmL9lOHdvuVi6cRN5tGGqYgwlRYC/RvtcElmVhSQn8VVJd3sQ2fOUZAY3kAT0xLl73S560FD
4egR4JlOVRzXJ/VYwjXXkk071sGTnL6xT1AE3gHJb01n4/IXJSqY6pgnIFWv+SJytOYz+DtD8Qbt
ygpucRTPtgX0SxMUyxg1mykbG8MN2Hi6itpN+tuQNvWdE082pv1BSQUAEKMKRcWCkJcqsyy+T9Ol
jQ7LmoqurDg72s4igb0nlUNKDkZFmC8tk7mOPRLF2YY/WA+Vexgj47oy/b9MjBNNTvQ899dZbwRy
RBZVfwd2xEjGXCKpu9G/MAJk/SEux/HOxvPVyjDIOogIsNpe+SG/oZULOjWptRy9XlZTYPAiv+bh
IpOdhQy0fTGM9wNAn3kkvBZLN4byqk0+tGmHfWuWgJHs94uPIdP0PtHpq6yVU5jzu9imrj64QAF0
8SAKsZY8V+XYDBq8jN8NzwbVmAyAzwIc+o3NBpgJFn7MwT5mnyaW3q21E3IEctpiv2XPna74WJgo
qQdPKSqpFO5ERYL9baZLTdWTzwD5olYb3mH/vdPSJt+FLUN2IggfwsyuRvWtk8lNuGTOvv7gseD7
a0Z4Qq/ZJ7cc8Q7kFjb06ZX0SKIm9jsspav/taychJkOPAArwyMZnrykL5dqkTKMLpwpGV4vInGf
u6ZLGS9jZ4q9DCd29NT0wOxLPW8PNff8wvD8oo7gHgls0zV9n0PAF4Y1CdczwlYuGlRPbUy9EXc7
ZSjNmL5NnJS4/ZAFP4/cBmVUMXed5LRfmGAThfGXiimPAzNDpb1uLk+X7wgACCanH3y9El0Nn+M6
1vjJriMfHuE9jDGTpzHLWlJAMwKpVWpgre+9EtJcj6yZMJOovaxo0DuckV72m3ByqF2ZhQ84ljZ2
zu6ikSW8X4mC77MgAowXqpGlscnOqsxvrhwhYA4wBzpeL8FwR3dTJh9Chhvvol16zor42vf4gcON
i+gRca2KKAf9/Pq93uIMTsl36gO112qvrWGDwDKdL7ySUnJJspg+kmjQZ3j7263CX9z9jltf4gC4
ZBRJaQcPDWz/mCBrkQ4wtC9N2SmekHGeCog1vhGjFQH/zMGIe214ii7OQjm5Vj3x215MYf08Lrfh
7+KSh7wEw7n9WefCtkbjEkLsg4nHAC/RKCkMF/G9NxMNMEwX/6T2tmTR559g2x0szh7ZVeMV81gf
GaqJEejWBBasHHRvm52zUpjLvDeFGvnSz7YPbXXDov+0R/bJ5jD1Wh9l5axUlkn9YLvmCBletx9X
OdoDwifkNVOQi6glhvHCJVAA/Ps/GdFSJl6TcQtGNKWXoUe09yEnZIraupf4kehKqC5YMA/5/855
xb9s0az/EAiuJ3e+BwaysGPMZ61ZVhfvqfnBzaXthdO98UfK9rL9VtkwmExmx96J68OvHOOZDUIr
ao6dPLPv3eD9e/9sLhWSCz0CxV516lRtIdOdV4aD7yFW3oyf8oeVhmfLtxjQGEbJI8WNt2X3WYTI
5/E0BLg9Msx1AeISFM0i0J6Q/Htuum8B3wTi0gMD9GEJ8DLgo240l+Kv93OdFoBsrzY5Ah11tIg/
RhoZuhkGUlW3yyn/1KkJw1p/TPqtJlBZjjdkOreycXJLsyedFpWGDaYd98EEynWgtDd24d7EVPbG
N2yEsuGqzYFoqDXXRvbMAUL65J28fCfpkmOSoEtoHcnlZvJDqluXe0A1fwDaVjaPUHKK7HUZf2Sn
KMZw5ylIgkksgrOVK8qPnkB21oWB/VddPmv/uNfohMpxOdS/d9iQa+CxOCJHwNrs/Qp83Ociz+zc
IE2z/woefdIkHbFMf1mErYih5RQ211nASzM4j7lO4T7KV8DY9ghTg67XGvW5Zi6ffp0zxyJGpoaA
qYkt6YuX7qhmA28uY3ZBaUa5Ol5YjXdK+0hFmSW04uKVKIcVF9spHRwdZVP/Qu3uqwYof8d0KBgr
8jMuRt+SPIJpZQFZAimIX+ttfbB+/usaF4ErK9wxI/Dp22B1/xi+K2+PNvLp79UlnGO6U1+0euMA
Il/fNfLeEZ+VAwDz8JCbsD17Iuctem+Rc+3BMDVzPzqDt6ItGY70sqr1k9wLF81XyB0C+VRVf08l
hG7TymRUqzuS94IvA4Ha9dgIEStNvWaI0fvHusm7kDVVuxWLf5YFsdsStgJuAn+NL5DjyhZlu7Pg
+0J6YRrfSLwlSp4gNAjBaZOyFK9mNbwMQX0zjkVTcfTaUfjUOU4du1fmgIssHFLNxWmlACFp9YbY
yoqW7y1IzWQ+deH6dFuEnus1hft8qz+DOFZ3WA/epOllNiN8YcpqhjttdZId1NydAAnJvavZeQ7W
mOJvsxkxlT2Ai0TmzhWBnWGzmXmdPccjyAnVNvBYHOR3M6O9h115isdOiRgZETlzPxrD9u7nLbrh
+pJLlSQJjseCV4UHShrKQ9WfJJ7s9sAnAOGzqxRg6HO5Fdm+JA3dcJHWw6/t5rjEHShq8Eu90eMm
D2MCFR7M4yB8uQpkFnSD1/tePUyAZEHBXJrcfh4g3Whb6mzN/+kihn2BF0kQ3lJ4qs/10E/6S34M
7yfLY1l/3FVF6lIzoO3Bby7Fz1mRVbRJkMtgET9VBMLuogm6IushGkV52Un/7aI7Cb4XcuQ1c5nw
cVWYs5GKNv5Alt/RXWTv3o2aNwGc+u7dTxaDroRSVJQSmgTJIJY5B2PtnWiebZDZScTdfb+uCTPN
GmBY0BXn2ZXJfqLAJRGvBtdaUMtelb912PTb4oJn8cjP+Bs4VcycjIVolffxKK28VG839cwbcSLz
vzZcCBoo11ORxiCKabL6JWl6Ek7Y63TEZjDm2hWRe0kE/7p+nwCt0EfkzoJvCIKBIgm1xPahQ0tX
DjI/tCGuP1jOu+XqQEKFGgueUwPOB1YCwaVKlzj5rHlZEr/+C7FQlXTGHp5VO9cAsjkugtHRlLu3
ycPo9aYX4KFo2xdBg0oSXEjKcDi4g5ZKlKC+dYQAKxhBnCOtOZ6XQbkwf/Fid5JL4U/D1TfutRag
8oAl5Fl/0troY8fo44vdzdligtaA/N6ZMGbXlgbYX+E1wgbc/QYjYr4gJZiHf46yc1LnYNnv2ee7
2jk/qRXYG33XdiQ4RNstJtbiao7JL4Xtoq7xAIfwPW5XqEheywKd6kDQv72c24uNP1kvE9dKgQ3P
VjgwNUAx+PTc9ZPS0NBaqr7lOu0nVSX5zLi/nWMgQqikPDJWWRQmis2ync4/PKC04k7qPAB4IXv+
9tzoEGarBeh3rZduU6VwnOOX8uqjwPdTRh2QRqFLrHdGkcReQ62suVfD/OV9WEKvQiBPfqzOUKMv
UECoeJLP60v2C/teGrrI+SxXDMw9WL8FtsjXYrUsmZ6hZpM4xJI1B5Y7Getp4s2Fd1VY8OEALQ4c
f6N92xS5464go4Xsbi8atAx4Nvw7dgy6t18iO+j82AKnQ5Z+SDrsVQ/XupEcy5632pWzsE9Mh7vu
l9bqpcg1iS8sK2YmqziKsTnoMrTPXhmFsuIJko1MV5bqE9gvoidbgssCZNkbKRnlZuvOvQ1IWnKG
5QBEhvd9AZ0UZCcus0LktFrVreHNhLdDHmphECh64PjafMp5dUbRtWpSCb7+QBY4aPf/pM+FZlNi
82je7C5fWx2Bl1/7Unb5Pr3O8QKSsrh0VPwYLX6I0NmL3sCVH84IPV9sx0VmqNMto31/uHA82Q4J
ERU3D9Jc6KVDG1DB+FRQIQi5Qeo11oSH43Oj0Hc+aTRk9lfK0nX0tLGmqtopbSuBxOdAhUi8sWVs
c+qSqmPH4kceHjNc/blz5N5z82FttljFIJ/fcnRp27gnQ/8A+1+rwuuyzA/aUNDJA5Dnhrky5Irq
nu/UsJj/nGE0+fSizPU1louNQop9RVtLgCKAVKi340i5oylcQ9JD6vnGYawUE3BtwkISplelrhSH
skO5gUnyli8wCUo2zigoIW6qykLbdLICvr1unIpoFNjwYeCAmoCF5bOJdeT+wwHQKz3Fd2z2bO/L
VQu2eYghFMuHnz+rGt26XXYF+8CC2BvDVgLxqOgv1ka/VFIXoOajC6gsb6cMabMWEDJme7zyBzyo
2V+OwW4/kXFhLBgn19HXEh5CKBYX/6B7So8ZyGVxEh+m2z+K8WD4AhXqyxQACseu1uEsVRSjBdYB
+BRBJw2NZoGKFzwMAJKwGZQ2dQ8whA+2VZYJmU8wb4Ll+hcUVUmtrmb9dJ2yq7rFgGGYdkmF4aOl
DEgQAfbPvDOGho8oZkfd3zM5chKqqCrkzQVpkI53aUSlhl1zmPccnefEoVSMujPqRr0EVbx0Ioae
r4UgA3VvRzr4QqW4aWzsOJ4nm2QIjH5QTOeh5hVDM9Md3m82t7J0eWr7cxCPszogwE9hcSgv37qd
y6FtyE4vUcytpt0L9v1pCR2GaRxLxcrRU5q1v7FP6hK4WKBhfC+9PnFqJLfapYCVDtrXGPSD8NDc
IEyShZ++j5Nm1g/CTySw9SPUfI+/zyrznLzHpk6Hsblk8fANS0GbC6Vo+31Oy2qFKuLWv2cW5VpK
Ss45KG5hnbWAPqsiGXv8QC4v4Q1S2+b5chffUDwAc7Zkgfx3MAkDO4MfMHpz/Afdzkse/BEIUYJd
PxUR5jRAe/m/ZjevztnMetI636X31jvhD0eQWnHqZ4tBhGRM1UjjoFnNYIkD1W8vo55MutnHdkNi
kf3v3dgOVUgC4H0A4PzBRiqC89GtiE1INi1urM02k8DsugtOxxmQQ0zWoF6vcsQPHnQOTCWl7eTz
uVn7B3KFhWK4wuyBN5+0YpdnNWLrg++Jv3iyzfD7Frlj3UPl3G2mTm//4Evw+5FBu8wm9a3Y5I4p
imKnCTeNkmcEcz/pX2wZtliCRlZF+ogRVoi5kIbjr8XJvjlaCSvobKJ26FTheO7l2+LUnWdgdmcz
R1oU3y6CTjFbWG+AdiNorAg/vcfpzAW2AA8zoG4zrCLqZkqPvxlaXxH4k0MCuSfPdqCVpkoiiVhT
RRs1NniMabNeWB/o5iPGSFWD3qj4HypC8Gs1t4MkFXxVSvS5fW3A1ExI8mT7CtEK81JE+dV56ACH
fAXZEGDmNL68FlhvxnKTXsbFe+42IWB9NEasVhi5/c9nHR19ay9SM0FkjY+7eXNYRRaASeXByGcN
bIYH54cK+h/AWF1koLt0Dg69UeWsAVNjujlxPQG1w9I2oWTHceHgYt72oYDZb40r+6Ck325lL8UQ
0GeITHIl8H260CmKCyjMrb448EXeUGVFuyQuRWcVcD9KcQjd/Urthqtb1KBXq3KS9XLIi/v3otx5
7flIfKUAbWXAj6ZpsReUy/xehKvrn9rJ5UAXnky1b+JVz/3YgHhZC2Xs925Eu/k3U29x6WyU3Kde
QwL3r6EMN/sCBatKIMlu9opMUgzo8+SxaF64dU9ZNOBhQ4d4Ic/iyF8UJ17FuoaoFsxxpWAZWUuA
fRynliL97Dq1Y5V/R/AxbsskBVX+/edWsU6B9GBdCyYNrWFgxSUM544XAn7sUKTTidZlHVyCAANv
cQHjGFRdXBwWNT8RVAMzPrfRRlopY482aJmQ2zzg/qduD37bTidFvzEK3BMKpepfzM900wisbSav
m7i2PFjYjOH5QnFcjuWnbMtbe1QtNqjIDjGJ2GllqA7Wr69Z1aCDNUTzWPl8GERWr5Yfp+1HmUP2
9/LfbyW2Og34ZlnRhFfLwuPVIr+CKJC8fnXY1T/c1f/rS3XLo4jLnEmshIeTkHnQuTaN1QR6u62K
VDp7qRke475GZiOMB2NZogWYaMTmNrn0MdKLx9lS1TmxqQQz2DN/bigCq9omNJmjBLthlWlI5VcA
B3dDzIMeNK2M5vTWXcIvtQlge8Gl0BOM6jJvRdKZu2Gg6A5727fHEBjs5yxKh5nD1XyDItOLFjjA
6LCpOhSCceZyiIOzbsTMKfv/vB7rQJPoDvxmDJ1aiFlNhlsMAwWJyHyzgN41kDabuen3jaUjFIbL
y9hvPZKEjBbet+KrXO5M780jT6tCq1h7zHXQnhmFaNXxPGPUYaeqX09UzYv1D+KxtVvEw4KjNbzs
hzDSP28KhNYSCFQ3efF+Pr/xZP6ikzDWH/GGCg5piJIwrlQcE8V6YA6ss5IJok69euEa5xyRh9uI
7yU7OP+pFTaiidH+cKaFpznwYdKStOxMGoWs4KfAUPqOrO/6vVc1u5zsXcZ9O1AYJYxIGXdP4SLO
dBEfTXVs8wFSUxQ9703z0SU3vS665UPv76KWPiVtpkXa3ssj0qdBwE8d2ScCqll1rbS2mcWnVAQT
b/6yCCH61NquX5DHy2yLemXbqhE8y6TtCARNBppYInCVNLUwHZYIYHBLnPJrAeaZwW2taCw01kgp
n4Kz6brjmqdq4bXZWEQ5yN47nPtdgaYl3PaNg5N0WNo2NplOUNQTRYMRuu2iCuxEJh5WbvqiTd4K
TTlSqpbmneN62bz94kMXu+K4bSGYRPIy8NkrL4mUa2yAuuGUwnRS2RNsN5ETK6EV2CYtfx8hfG2G
2mpgW8srGslQ8v9ahm95IWAh7KOyJUp/fuE80/Dt+vp+eJ7rHOh7qqskAn+QXo9YItcKr5/wda/J
uYQKL7t/gIT2SX30S/bugg84+tAN9F1Rc+N3XhqOwv94pVgYviHuigNLOHR9RgvsTKrWgs4oQW7h
Y9xLQev4Lu0/0Ctucsj+HbqRcTH9nxgMu62FJQVtdPRTSNC7lcoa+GQUDPbBdpdB6bDJuc0+YnYi
9NwsGPsP7g7uZ5mqBWEINzfYED8wKn8ShGKmPrYTvMc7qEKoqEI8Ajos4yTZezMAQMw82l9gsYbi
PKRxdzjfyjPB1z8cWraUdLXfUFaETxZHmRUGP98fKYxtGTaEEpnv3WXlJg1ASTYseg+6xsAdOA8/
NNnD8zsav4Io1OKVmC8z67KdH3e9xoRmuXWj5V+4Q3RQsxopLZx12iHQb+t3RZ1GAO/zXteDwo2r
D+/wy9+KyM3xhGZs5naqil5FN+WTZRFPlw2aQZ4x99DTLhlpH9445Z11PToLreCvGM08BC0IgvuU
oPc0rXOnD1hSmSoXkhK8sEwDTqIUC8jBjmlNKNJKQ0cebamFnyBR+wvoL3nuN/h8cUIF2hIPPgKW
fmo1fwFtsbyKjI+/V8htDj2yeHZZnQa/bs9+SfwHzsvl0p5QudGx6tle2eRbLo9azrlpXj3HFLoB
gNJmLaGeDeguO87NrlK4di1V3FEN/SQWCMBwOUx+1lA6VuYZtl4e4UN66hR86kG6y1gHOpWFrbeB
EnsnptxgZQiiWxU6uTd4/vo1dqcaCstStwdsXc4gPAu34VeISvW+j/hApSd5aLpPs5GxHOHGZd2N
6Hp2LQXLSa015nOi/+b9Zxdxj6FdZpcl1E3zs22auZc2fm4Oiy7wJBC/HJa94vc5166F2wILiidR
Lw6HUf/V5w6eoMvGZgd32wQFO8+Mw69gnn2F8EtvETpSJeIfLVFDSRLegccFwWwG2x0r9XksC5+w
2UxnYx7TUM66nXfHRVpGX267yWnX/31g2k/QSMMqvenxPLGkBGMtqsugAWHZH4W27z0I0dmfIdz6
Yx81eZnLwryzS56M4Jtl2OMylEZ8EujT2WNUmigqSjiQxlVpVAoOKhOvmJHtvwHypWXE7hgOiDD0
m+ZGv0LwaElHHynlekws5LJyUKI0qE2vhNIOKabS6ggPZuI9zCoJlDHXA1ZOWbzVW/5mrqhlaINd
a+TnySf2MFcSEtrTT/iOqIU6LR5e1Zbja6KyE4al2eYSC2VDqJ8SC8hzO/ZBknumvd53P1xQ5ZV/
mT2tzK53YClubwXz4/jhdT60xwlOZ2JGqsOgloOK8itswN+BAmBjgQQHl2vqVj5Ms5QakXEI
`protect end_protected
